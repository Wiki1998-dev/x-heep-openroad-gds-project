// removed package "top_pkg"
// removed package "ibex_pkg"
// removed package "spi_device_reg_pkg"
// removed package "spi_device_pkg"
// removed package "prim_pkg"
// removed package "prim_cipher_pkg"
// removed package "prim_secded_pkg"
// removed package "prim_util_pkg"
// removed package "cv32e40p_apu_core_pkg"
// removed package "cv32e40p_fpu_pkg"
// removed package "cv32e40p_pkg"
// removed package "cb_filter_pkg"
// removed package "cf_math_pkg"
// removed package "ecc_pkg"
// removed package "cdc_reset_ctrlr_pkg"
// removed package "dm"
// removed package "addr_map_rule_pkg"
// removed package "obi_pkg"
// removed package "reg_pkg"
// removed package "core_v_mini_mcu_pkg"
// removed package "power_manager_reg_pkg"
// removed package "tlul_pkg"
// removed package "fpnew_pkg"
// removed package "gpio_reg_pkg"
// removed package "dma_reg_pkg"
// removed package "obi_spimemio_reg_pkg"
// removed package "picorv32_pkg"
// removed package "prim_alert_pkg"
// removed package "prim_esc_pkg"
// removed package "spi_host_reg_pkg"
// removed package "spi_host_cmd_pkg"
// removed package "soc_ctrl_reg_pkg"
// removed package "fast_intr_ctrl_reg_pkg"
// removed package "i2c_reg_pkg"
// removed package "rv_plic_reg_pkg"
// removed package "rv_timer_reg_pkg"
// removed package "uart_reg_pkg"
// removed package "top_pkg"
// removed package "ibex_pkg"
// removed package "spi_device_reg_pkg"
// removed package "spi_device_pkg"
// removed package "prim_pkg"
// removed package "prim_cipher_pkg"
module prim_generic_buf (
	in_i,
	out_o
);
	// Trace: design.sv:1654:13
	parameter signed [31:0] Width = 1;
	// Trace: design.sv:1656:3
	input [Width - 1:0] in_i;
	// Trace: design.sv:1657:3
	output wire [Width - 1:0] out_o;
	// Trace: design.sv:1660:3
	assign out_o = in_i;
endmodule
module prim_generic_flop (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	// Trace: design.sv:1670:13
	parameter signed [31:0] Width = 1;
	// Trace: design.sv:1671:13
	parameter [Width - 1:0] ResetValue = 0;
	// Trace: design.sv:1673:3
	input clk_i;
	// Trace: design.sv:1674:3
	input rst_ni;
	// Trace: design.sv:1675:3
	input [Width - 1:0] d_i;
	// Trace: design.sv:1676:3
	output reg [Width - 1:0] q_o;
	// Trace: design.sv:1679:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:1680:5
		if (!rst_ni)
			// Trace: design.sv:1681:7
			q_o <= ResetValue;
		else
			// Trace: design.sv:1683:7
			q_o <= d_i;
endmodule
module prim_generic_flop_2sync (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	// Trace: design.sv:1697:13
	parameter signed [31:0] Width = 16;
	// Trace: design.sv:1698:13
	parameter [Width - 1:0] ResetValue = 1'sb0;
	// Trace: design.sv:1700:3
	input clk_i;
	// Trace: design.sv:1701:3
	input rst_ni;
	// Trace: design.sv:1702:3
	input [Width - 1:0] d_i;
	// Trace: design.sv:1703:3
	output wire [Width - 1:0] q_o;
	// Trace: design.sv:1706:3
	wire [Width - 1:0] intq;
	// Trace: design.sv:1708:3
	prim_flop #(
		.Width(Width),
		.ResetValue(ResetValue)
	) u_sync_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(d_i),
		.q_o(intq)
	);
	// Trace: design.sv:1718:3
	prim_flop #(
		.Width(Width),
		.ResetValue(ResetValue)
	) u_sync_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(intq),
		.q_o(q_o)
	);
endmodule
module prim_generic_flop_en (
	clk_i,
	rst_ni,
	en_i,
	d_i,
	q_o
);
	// Trace: design.sv:1736:13
	parameter signed [31:0] Width = 1;
	// Trace: design.sv:1737:13
	parameter [Width - 1:0] ResetValue = 0;
	// Trace: design.sv:1739:3
	input clk_i;
	// Trace: design.sv:1740:3
	input rst_ni;
	// Trace: design.sv:1741:3
	input en_i;
	// Trace: design.sv:1742:3
	input [Width - 1:0] d_i;
	// Trace: design.sv:1743:3
	output reg [Width - 1:0] q_o;
	// Trace: design.sv:1746:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:1747:5
		if (!rst_ni)
			// Trace: design.sv:1748:7
			q_o <= ResetValue;
		else if (en_i)
			// Trace: design.sv:1750:7
			q_o <= d_i;
endmodule
module prim_generic_xor2 (
	in0_i,
	in1_i,
	out_o
);
	// Trace: design.sv:1762:13
	parameter signed [31:0] Width = 1;
	// Trace: design.sv:1764:3
	input [Width - 1:0] in0_i;
	// Trace: design.sv:1765:3
	input [Width - 1:0] in1_i;
	// Trace: design.sv:1766:3
	output wire [Width - 1:0] out_o;
	// Trace: design.sv:1769:3
	assign out_o = in0_i ^ in1_i;
endmodule
// removed package "prim_secded_pkg"
module prim_secded_22_16_dec (
	in,
	d_o,
	syndrome_o,
	err_o
);
	// Trace: design.sv:2493:3
	input [21:0] in;
	// Trace: design.sv:2494:3
	output wire [15:0] d_o;
	// Trace: design.sv:2495:3
	output wire [5:0] syndrome_o;
	// Trace: design.sv:2496:3
	output wire [1:0] err_o;
	// Trace: design.sv:2499:3
	wire single_error;
	// Trace: design.sv:2502:3
	assign syndrome_o[0] = ^(in & 22'h01496e);
	// Trace: design.sv:2503:3
	assign syndrome_o[1] = ^(in & 22'h02f20b);
	// Trace: design.sv:2504:3
	assign syndrome_o[2] = ^(in & 22'h048ed8);
	// Trace: design.sv:2505:3
	assign syndrome_o[3] = ^(in & 22'h087714);
	// Trace: design.sv:2506:3
	assign syndrome_o[4] = ^(in & 22'h10aca5);
	// Trace: design.sv:2507:3
	assign syndrome_o[5] = ^(in & 22'h2011f3);
	// Trace: design.sv:2510:3
	assign d_o[0] = (syndrome_o == 6'h32) ^ in[0];
	// Trace: design.sv:2511:3
	assign d_o[1] = (syndrome_o == 6'h23) ^ in[1];
	// Trace: design.sv:2512:3
	assign d_o[2] = (syndrome_o == 6'h19) ^ in[2];
	// Trace: design.sv:2513:3
	assign d_o[3] = (syndrome_o == 6'h07) ^ in[3];
	// Trace: design.sv:2514:3
	assign d_o[4] = (syndrome_o == 6'h2c) ^ in[4];
	// Trace: design.sv:2515:3
	assign d_o[5] = (syndrome_o == 6'h31) ^ in[5];
	// Trace: design.sv:2516:3
	assign d_o[6] = (syndrome_o == 6'h25) ^ in[6];
	// Trace: design.sv:2517:3
	assign d_o[7] = (syndrome_o == 6'h34) ^ in[7];
	// Trace: design.sv:2518:3
	assign d_o[8] = (syndrome_o == 6'h29) ^ in[8];
	// Trace: design.sv:2519:3
	assign d_o[9] = (syndrome_o == 6'h0e) ^ in[9];
	// Trace: design.sv:2520:3
	assign d_o[10] = (syndrome_o == 6'h1c) ^ in[10];
	// Trace: design.sv:2521:3
	assign d_o[11] = (syndrome_o == 6'h15) ^ in[11];
	// Trace: design.sv:2522:3
	assign d_o[12] = (syndrome_o == 6'h2a) ^ in[12];
	// Trace: design.sv:2523:3
	assign d_o[13] = (syndrome_o == 6'h1a) ^ in[13];
	// Trace: design.sv:2524:3
	assign d_o[14] = (syndrome_o == 6'h0b) ^ in[14];
	// Trace: design.sv:2525:3
	assign d_o[15] = (syndrome_o == 6'h16) ^ in[15];
	// Trace: design.sv:2528:3
	assign single_error = ^syndrome_o;
	// Trace: design.sv:2529:3
	assign err_o[0] = single_error;
	// Trace: design.sv:2530:3
	assign err_o[1] = ~single_error & |syndrome_o;
endmodule
module prim_secded_22_16_enc (
	in,
	out
);
	reg _sv2v_0;
	// Trace: design.sv:2540:3
	input [15:0] in;
	// Trace: design.sv:2541:3
	output reg [21:0] out;
	// Trace: design.sv:2544:3
	function automatic [21:0] sv2v_cast_22;
		input reg [21:0] inp;
		sv2v_cast_22 = inp;
	endfunction
	always @(*) begin : p_encode
		if (_sv2v_0)
			;
		// Trace: design.sv:2545:5
		out = sv2v_cast_22(in);
		// Trace: design.sv:2546:5
		out[16] = ^(out & 22'h00496e);
		// Trace: design.sv:2547:5
		out[17] = ^(out & 22'h00f20b);
		// Trace: design.sv:2548:5
		out[18] = ^(out & 22'h008ed8);
		// Trace: design.sv:2549:5
		out[19] = ^(out & 22'h007714);
		// Trace: design.sv:2550:5
		out[20] = ^(out & 22'h00aca5);
		// Trace: design.sv:2551:5
		out[21] = ^(out & 22'h0011f3);
	end
	initial _sv2v_0 = 0;
endmodule
module prim_secded_28_22_dec (
	in,
	d_o,
	syndrome_o,
	err_o
);
	// Trace: design.sv:2562:3
	input [27:0] in;
	// Trace: design.sv:2563:3
	output wire [21:0] d_o;
	// Trace: design.sv:2564:3
	output wire [5:0] syndrome_o;
	// Trace: design.sv:2565:3
	output wire [1:0] err_o;
	// Trace: design.sv:2568:3
	wire single_error;
	// Trace: design.sv:2571:3
	assign syndrome_o[0] = ^(in & 28'h07003ff);
	// Trace: design.sv:2572:3
	assign syndrome_o[1] = ^(in & 28'h090fc0f);
	// Trace: design.sv:2573:3
	assign syndrome_o[2] = ^(in & 28'h1271c71);
	// Trace: design.sv:2574:3
	assign syndrome_o[3] = ^(in & 28'h23b6592);
	// Trace: design.sv:2575:3
	assign syndrome_o[4] = ^(in & 28'h43daaa4);
	// Trace: design.sv:2576:3
	assign syndrome_o[5] = ^(in & 28'h83ed348);
	// Trace: design.sv:2579:3
	assign d_o[0] = (syndrome_o == 6'h07) ^ in[0];
	// Trace: design.sv:2580:3
	assign d_o[1] = (syndrome_o == 6'h0b) ^ in[1];
	// Trace: design.sv:2581:3
	assign d_o[2] = (syndrome_o == 6'h13) ^ in[2];
	// Trace: design.sv:2582:3
	assign d_o[3] = (syndrome_o == 6'h23) ^ in[3];
	// Trace: design.sv:2583:3
	assign d_o[4] = (syndrome_o == 6'h0d) ^ in[4];
	// Trace: design.sv:2584:3
	assign d_o[5] = (syndrome_o == 6'h15) ^ in[5];
	// Trace: design.sv:2585:3
	assign d_o[6] = (syndrome_o == 6'h25) ^ in[6];
	// Trace: design.sv:2586:3
	assign d_o[7] = (syndrome_o == 6'h19) ^ in[7];
	// Trace: design.sv:2587:3
	assign d_o[8] = (syndrome_o == 6'h29) ^ in[8];
	// Trace: design.sv:2588:3
	assign d_o[9] = (syndrome_o == 6'h31) ^ in[9];
	// Trace: design.sv:2589:3
	assign d_o[10] = (syndrome_o == 6'h0e) ^ in[10];
	// Trace: design.sv:2590:3
	assign d_o[11] = (syndrome_o == 6'h16) ^ in[11];
	// Trace: design.sv:2591:3
	assign d_o[12] = (syndrome_o == 6'h26) ^ in[12];
	// Trace: design.sv:2592:3
	assign d_o[13] = (syndrome_o == 6'h1a) ^ in[13];
	// Trace: design.sv:2593:3
	assign d_o[14] = (syndrome_o == 6'h2a) ^ in[14];
	// Trace: design.sv:2594:3
	assign d_o[15] = (syndrome_o == 6'h32) ^ in[15];
	// Trace: design.sv:2595:3
	assign d_o[16] = (syndrome_o == 6'h1c) ^ in[16];
	// Trace: design.sv:2596:3
	assign d_o[17] = (syndrome_o == 6'h2c) ^ in[17];
	// Trace: design.sv:2597:3
	assign d_o[18] = (syndrome_o == 6'h34) ^ in[18];
	// Trace: design.sv:2598:3
	assign d_o[19] = (syndrome_o == 6'h38) ^ in[19];
	// Trace: design.sv:2599:3
	assign d_o[20] = (syndrome_o == 6'h3b) ^ in[20];
	// Trace: design.sv:2600:3
	assign d_o[21] = (syndrome_o == 6'h3d) ^ in[21];
	// Trace: design.sv:2603:3
	assign single_error = ^syndrome_o;
	// Trace: design.sv:2604:3
	assign err_o[0] = single_error;
	// Trace: design.sv:2605:3
	assign err_o[1] = ~single_error & |syndrome_o;
endmodule
module prim_secded_28_22_enc (
	in,
	out
);
	reg _sv2v_0;
	// Trace: design.sv:2615:3
	input [21:0] in;
	// Trace: design.sv:2616:3
	output reg [27:0] out;
	// Trace: design.sv:2619:3
	function automatic [27:0] sv2v_cast_28;
		input reg [27:0] inp;
		sv2v_cast_28 = inp;
	endfunction
	always @(*) begin : p_encode
		if (_sv2v_0)
			;
		// Trace: design.sv:2620:5
		out = sv2v_cast_28(in);
		// Trace: design.sv:2621:5
		out[22] = ^(out & 28'h03003ff);
		// Trace: design.sv:2622:5
		out[23] = ^(out & 28'h010fc0f);
		// Trace: design.sv:2623:5
		out[24] = ^(out & 28'h0271c71);
		// Trace: design.sv:2624:5
		out[25] = ^(out & 28'h03b6592);
		// Trace: design.sv:2625:5
		out[26] = ^(out & 28'h03daaa4);
		// Trace: design.sv:2626:5
		out[27] = ^(out & 28'h03ed348);
	end
	initial _sv2v_0 = 0;
endmodule
module prim_secded_39_32_dec (
	in,
	d_o,
	syndrome_o,
	err_o
);
	// Trace: design.sv:2637:3
	input [38:0] in;
	// Trace: design.sv:2638:3
	output wire [31:0] d_o;
	// Trace: design.sv:2639:3
	output wire [6:0] syndrome_o;
	// Trace: design.sv:2640:3
	output wire [1:0] err_o;
	// Trace: design.sv:2643:3
	wire single_error;
	// Trace: design.sv:2646:3
	assign syndrome_o[0] = ^(in & 39'h012606bd25);
	// Trace: design.sv:2647:3
	assign syndrome_o[1] = ^(in & 39'h02deba8050);
	// Trace: design.sv:2648:3
	assign syndrome_o[2] = ^(in & 39'h04413d89aa);
	// Trace: design.sv:2649:3
	assign syndrome_o[3] = ^(in & 39'h0831234ed1);
	// Trace: design.sv:2650:3
	assign syndrome_o[4] = ^(in & 39'h10c2c1323b);
	// Trace: design.sv:2651:3
	assign syndrome_o[5] = ^(in & 39'h202dcc624c);
	// Trace: design.sv:2652:3
	assign syndrome_o[6] = ^(in & 39'h4098505586);
	// Trace: design.sv:2655:3
	assign d_o[0] = (syndrome_o == 7'h19) ^ in[0];
	// Trace: design.sv:2656:3
	assign d_o[1] = (syndrome_o == 7'h54) ^ in[1];
	// Trace: design.sv:2657:3
	assign d_o[2] = (syndrome_o == 7'h61) ^ in[2];
	// Trace: design.sv:2658:3
	assign d_o[3] = (syndrome_o == 7'h34) ^ in[3];
	// Trace: design.sv:2659:3
	assign d_o[4] = (syndrome_o == 7'h1a) ^ in[4];
	// Trace: design.sv:2660:3
	assign d_o[5] = (syndrome_o == 7'h15) ^ in[5];
	// Trace: design.sv:2661:3
	assign d_o[6] = (syndrome_o == 7'h2a) ^ in[6];
	// Trace: design.sv:2662:3
	assign d_o[7] = (syndrome_o == 7'h4c) ^ in[7];
	// Trace: design.sv:2663:3
	assign d_o[8] = (syndrome_o == 7'h45) ^ in[8];
	// Trace: design.sv:2664:3
	assign d_o[9] = (syndrome_o == 7'h38) ^ in[9];
	// Trace: design.sv:2665:3
	assign d_o[10] = (syndrome_o == 7'h49) ^ in[10];
	// Trace: design.sv:2666:3
	assign d_o[11] = (syndrome_o == 7'h0d) ^ in[11];
	// Trace: design.sv:2667:3
	assign d_o[12] = (syndrome_o == 7'h51) ^ in[12];
	// Trace: design.sv:2668:3
	assign d_o[13] = (syndrome_o == 7'h31) ^ in[13];
	// Trace: design.sv:2669:3
	assign d_o[14] = (syndrome_o == 7'h68) ^ in[14];
	// Trace: design.sv:2670:3
	assign d_o[15] = (syndrome_o == 7'h07) ^ in[15];
	// Trace: design.sv:2671:3
	assign d_o[16] = (syndrome_o == 7'h1c) ^ in[16];
	// Trace: design.sv:2672:3
	assign d_o[17] = (syndrome_o == 7'h0b) ^ in[17];
	// Trace: design.sv:2673:3
	assign d_o[18] = (syndrome_o == 7'h25) ^ in[18];
	// Trace: design.sv:2674:3
	assign d_o[19] = (syndrome_o == 7'h26) ^ in[19];
	// Trace: design.sv:2675:3
	assign d_o[20] = (syndrome_o == 7'h46) ^ in[20];
	// Trace: design.sv:2676:3
	assign d_o[21] = (syndrome_o == 7'h0e) ^ in[21];
	// Trace: design.sv:2677:3
	assign d_o[22] = (syndrome_o == 7'h70) ^ in[22];
	// Trace: design.sv:2678:3
	assign d_o[23] = (syndrome_o == 7'h32) ^ in[23];
	// Trace: design.sv:2679:3
	assign d_o[24] = (syndrome_o == 7'h2c) ^ in[24];
	// Trace: design.sv:2680:3
	assign d_o[25] = (syndrome_o == 7'h13) ^ in[25];
	// Trace: design.sv:2681:3
	assign d_o[26] = (syndrome_o == 7'h23) ^ in[26];
	// Trace: design.sv:2682:3
	assign d_o[27] = (syndrome_o == 7'h62) ^ in[27];
	// Trace: design.sv:2683:3
	assign d_o[28] = (syndrome_o == 7'h4a) ^ in[28];
	// Trace: design.sv:2684:3
	assign d_o[29] = (syndrome_o == 7'h29) ^ in[29];
	// Trace: design.sv:2685:3
	assign d_o[30] = (syndrome_o == 7'h16) ^ in[30];
	// Trace: design.sv:2686:3
	assign d_o[31] = (syndrome_o == 7'h52) ^ in[31];
	// Trace: design.sv:2689:3
	assign single_error = ^syndrome_o;
	// Trace: design.sv:2690:3
	assign err_o[0] = single_error;
	// Trace: design.sv:2691:3
	assign err_o[1] = ~single_error & |syndrome_o;
endmodule
module prim_secded_39_32_enc (
	in,
	out
);
	reg _sv2v_0;
	// Trace: design.sv:2701:3
	input [31:0] in;
	// Trace: design.sv:2702:3
	output reg [38:0] out;
	// Trace: design.sv:2705:3
	function automatic [38:0] sv2v_cast_39;
		input reg [38:0] inp;
		sv2v_cast_39 = inp;
	endfunction
	always @(*) begin : p_encode
		if (_sv2v_0)
			;
		// Trace: design.sv:2706:5
		out = sv2v_cast_39(in);
		// Trace: design.sv:2707:5
		out[32] = ^(out & 39'h002606bd25);
		// Trace: design.sv:2708:5
		out[33] = ^(out & 39'h00deba8050);
		// Trace: design.sv:2709:5
		out[34] = ^(out & 39'h00413d89aa);
		// Trace: design.sv:2710:5
		out[35] = ^(out & 39'h0031234ed1);
		// Trace: design.sv:2711:5
		out[36] = ^(out & 39'h00c2c1323b);
		// Trace: design.sv:2712:5
		out[37] = ^(out & 39'h002dcc624c);
		// Trace: design.sv:2713:5
		out[38] = ^(out & 39'h0098505586);
	end
	initial _sv2v_0 = 0;
endmodule
module prim_secded_64_57_dec (
	in,
	d_o,
	syndrome_o,
	err_o
);
	// Trace: design.sv:2724:3
	input [63:0] in;
	// Trace: design.sv:2725:3
	output wire [56:0] d_o;
	// Trace: design.sv:2726:3
	output wire [6:0] syndrome_o;
	// Trace: design.sv:2727:3
	output wire [1:0] err_o;
	// Trace: design.sv:2730:3
	wire single_error;
	// Trace: design.sv:2733:3
	assign syndrome_o[0] = ^(in & 64'h0303fff800007fff);
	// Trace: design.sv:2734:3
	assign syndrome_o[1] = ^(in & 64'h057c1ff801ff801f);
	// Trace: design.sv:2735:3
	assign syndrome_o[2] = ^(in & 64'h09bde1f87e0781e1);
	// Trace: design.sv:2736:3
	assign syndrome_o[3] = ^(in & 64'h11deee3b8e388e22);
	// Trace: design.sv:2737:3
	assign syndrome_o[4] = ^(in & 64'h21ef76cdb2c93244);
	// Trace: design.sv:2738:3
	assign syndrome_o[5] = ^(in & 64'h41f7bb56d5525488);
	// Trace: design.sv:2739:3
	assign syndrome_o[6] = ^(in & 64'h81fbdda769a46910);
	// Trace: design.sv:2742:3
	assign d_o[0] = (syndrome_o == 7'h07) ^ in[0];
	// Trace: design.sv:2743:3
	assign d_o[1] = (syndrome_o == 7'h0b) ^ in[1];
	// Trace: design.sv:2744:3
	assign d_o[2] = (syndrome_o == 7'h13) ^ in[2];
	// Trace: design.sv:2745:3
	assign d_o[3] = (syndrome_o == 7'h23) ^ in[3];
	// Trace: design.sv:2746:3
	assign d_o[4] = (syndrome_o == 7'h43) ^ in[4];
	// Trace: design.sv:2747:3
	assign d_o[5] = (syndrome_o == 7'h0d) ^ in[5];
	// Trace: design.sv:2748:3
	assign d_o[6] = (syndrome_o == 7'h15) ^ in[6];
	// Trace: design.sv:2749:3
	assign d_o[7] = (syndrome_o == 7'h25) ^ in[7];
	// Trace: design.sv:2750:3
	assign d_o[8] = (syndrome_o == 7'h45) ^ in[8];
	// Trace: design.sv:2751:3
	assign d_o[9] = (syndrome_o == 7'h19) ^ in[9];
	// Trace: design.sv:2752:3
	assign d_o[10] = (syndrome_o == 7'h29) ^ in[10];
	// Trace: design.sv:2753:3
	assign d_o[11] = (syndrome_o == 7'h49) ^ in[11];
	// Trace: design.sv:2754:3
	assign d_o[12] = (syndrome_o == 7'h31) ^ in[12];
	// Trace: design.sv:2755:3
	assign d_o[13] = (syndrome_o == 7'h51) ^ in[13];
	// Trace: design.sv:2756:3
	assign d_o[14] = (syndrome_o == 7'h61) ^ in[14];
	// Trace: design.sv:2757:3
	assign d_o[15] = (syndrome_o == 7'h0e) ^ in[15];
	// Trace: design.sv:2758:3
	assign d_o[16] = (syndrome_o == 7'h16) ^ in[16];
	// Trace: design.sv:2759:3
	assign d_o[17] = (syndrome_o == 7'h26) ^ in[17];
	// Trace: design.sv:2760:3
	assign d_o[18] = (syndrome_o == 7'h46) ^ in[18];
	// Trace: design.sv:2761:3
	assign d_o[19] = (syndrome_o == 7'h1a) ^ in[19];
	// Trace: design.sv:2762:3
	assign d_o[20] = (syndrome_o == 7'h2a) ^ in[20];
	// Trace: design.sv:2763:3
	assign d_o[21] = (syndrome_o == 7'h4a) ^ in[21];
	// Trace: design.sv:2764:3
	assign d_o[22] = (syndrome_o == 7'h32) ^ in[22];
	// Trace: design.sv:2765:3
	assign d_o[23] = (syndrome_o == 7'h52) ^ in[23];
	// Trace: design.sv:2766:3
	assign d_o[24] = (syndrome_o == 7'h62) ^ in[24];
	// Trace: design.sv:2767:3
	assign d_o[25] = (syndrome_o == 7'h1c) ^ in[25];
	// Trace: design.sv:2768:3
	assign d_o[26] = (syndrome_o == 7'h2c) ^ in[26];
	// Trace: design.sv:2769:3
	assign d_o[27] = (syndrome_o == 7'h4c) ^ in[27];
	// Trace: design.sv:2770:3
	assign d_o[28] = (syndrome_o == 7'h34) ^ in[28];
	// Trace: design.sv:2771:3
	assign d_o[29] = (syndrome_o == 7'h54) ^ in[29];
	// Trace: design.sv:2772:3
	assign d_o[30] = (syndrome_o == 7'h64) ^ in[30];
	// Trace: design.sv:2773:3
	assign d_o[31] = (syndrome_o == 7'h38) ^ in[31];
	// Trace: design.sv:2774:3
	assign d_o[32] = (syndrome_o == 7'h58) ^ in[32];
	// Trace: design.sv:2775:3
	assign d_o[33] = (syndrome_o == 7'h68) ^ in[33];
	// Trace: design.sv:2776:3
	assign d_o[34] = (syndrome_o == 7'h70) ^ in[34];
	// Trace: design.sv:2777:3
	assign d_o[35] = (syndrome_o == 7'h1f) ^ in[35];
	// Trace: design.sv:2778:3
	assign d_o[36] = (syndrome_o == 7'h2f) ^ in[36];
	// Trace: design.sv:2779:3
	assign d_o[37] = (syndrome_o == 7'h4f) ^ in[37];
	// Trace: design.sv:2780:3
	assign d_o[38] = (syndrome_o == 7'h37) ^ in[38];
	// Trace: design.sv:2781:3
	assign d_o[39] = (syndrome_o == 7'h57) ^ in[39];
	// Trace: design.sv:2782:3
	assign d_o[40] = (syndrome_o == 7'h67) ^ in[40];
	// Trace: design.sv:2783:3
	assign d_o[41] = (syndrome_o == 7'h3b) ^ in[41];
	// Trace: design.sv:2784:3
	assign d_o[42] = (syndrome_o == 7'h5b) ^ in[42];
	// Trace: design.sv:2785:3
	assign d_o[43] = (syndrome_o == 7'h6b) ^ in[43];
	// Trace: design.sv:2786:3
	assign d_o[44] = (syndrome_o == 7'h73) ^ in[44];
	// Trace: design.sv:2787:3
	assign d_o[45] = (syndrome_o == 7'h3d) ^ in[45];
	// Trace: design.sv:2788:3
	assign d_o[46] = (syndrome_o == 7'h5d) ^ in[46];
	// Trace: design.sv:2789:3
	assign d_o[47] = (syndrome_o == 7'h6d) ^ in[47];
	// Trace: design.sv:2790:3
	assign d_o[48] = (syndrome_o == 7'h75) ^ in[48];
	// Trace: design.sv:2791:3
	assign d_o[49] = (syndrome_o == 7'h79) ^ in[49];
	// Trace: design.sv:2792:3
	assign d_o[50] = (syndrome_o == 7'h3e) ^ in[50];
	// Trace: design.sv:2793:3
	assign d_o[51] = (syndrome_o == 7'h5e) ^ in[51];
	// Trace: design.sv:2794:3
	assign d_o[52] = (syndrome_o == 7'h6e) ^ in[52];
	// Trace: design.sv:2795:3
	assign d_o[53] = (syndrome_o == 7'h76) ^ in[53];
	// Trace: design.sv:2796:3
	assign d_o[54] = (syndrome_o == 7'h7a) ^ in[54];
	// Trace: design.sv:2797:3
	assign d_o[55] = (syndrome_o == 7'h7c) ^ in[55];
	// Trace: design.sv:2798:3
	assign d_o[56] = (syndrome_o == 7'h7f) ^ in[56];
	// Trace: design.sv:2801:3
	assign single_error = ^syndrome_o;
	// Trace: design.sv:2802:3
	assign err_o[0] = single_error;
	// Trace: design.sv:2803:3
	assign err_o[1] = ~single_error & |syndrome_o;
endmodule
module prim_secded_64_57_enc (
	in,
	out
);
	reg _sv2v_0;
	// Trace: design.sv:2813:3
	input [56:0] in;
	// Trace: design.sv:2814:3
	output reg [63:0] out;
	// Trace: design.sv:2817:3
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	always @(*) begin : p_encode
		if (_sv2v_0)
			;
		// Trace: design.sv:2818:5
		out = sv2v_cast_64(in);
		// Trace: design.sv:2819:5
		out[57] = ^(out & 64'h0103fff800007fff);
		// Trace: design.sv:2820:5
		out[58] = ^(out & 64'h017c1ff801ff801f);
		// Trace: design.sv:2821:5
		out[59] = ^(out & 64'h01bde1f87e0781e1);
		// Trace: design.sv:2822:5
		out[60] = ^(out & 64'h01deee3b8e388e22);
		// Trace: design.sv:2823:5
		out[61] = ^(out & 64'h01ef76cdb2c93244);
		// Trace: design.sv:2824:5
		out[62] = ^(out & 64'h01f7bb56d5525488);
		// Trace: design.sv:2825:5
		out[63] = ^(out & 64'h01fbdda769a46910);
	end
	initial _sv2v_0 = 0;
endmodule
module prim_secded_72_64_dec (
	in,
	d_o,
	syndrome_o,
	err_o
);
	// Trace: design.sv:2836:3
	input [71:0] in;
	// Trace: design.sv:2837:3
	output wire [63:0] d_o;
	// Trace: design.sv:2838:3
	output wire [7:0] syndrome_o;
	// Trace: design.sv:2839:3
	output wire [1:0] err_o;
	// Trace: design.sv:2842:3
	wire single_error;
	// Trace: design.sv:2845:3
	assign syndrome_o[0] = ^(in & 72'h01b9000000001fffff);
	// Trace: design.sv:2846:3
	assign syndrome_o[1] = ^(in & 72'h025e00000fffe0003f);
	// Trace: design.sv:2847:3
	assign syndrome_o[2] = ^(in & 72'h0467003ff003e007c1);
	// Trace: design.sv:2848:3
	assign syndrome_o[3] = ^(in & 72'h08cd0fc0f03c207842);
	// Trace: design.sv:2849:3
	assign syndrome_o[4] = ^(in & 72'h10b671c711c4438884);
	// Trace: design.sv:2850:3
	assign syndrome_o[5] = ^(in & 72'h20b5b65926488c9108);
	// Trace: design.sv:2851:3
	assign syndrome_o[6] = ^(in & 72'h40cbdaaa4a91152210);
	// Trace: design.sv:2852:3
	assign syndrome_o[7] = ^(in & 72'h807aed348d221a4420);
	// Trace: design.sv:2855:3
	assign d_o[0] = (syndrome_o == 8'h07) ^ in[0];
	// Trace: design.sv:2856:3
	assign d_o[1] = (syndrome_o == 8'h0b) ^ in[1];
	// Trace: design.sv:2857:3
	assign d_o[2] = (syndrome_o == 8'h13) ^ in[2];
	// Trace: design.sv:2858:3
	assign d_o[3] = (syndrome_o == 8'h23) ^ in[3];
	// Trace: design.sv:2859:3
	assign d_o[4] = (syndrome_o == 8'h43) ^ in[4];
	// Trace: design.sv:2860:3
	assign d_o[5] = (syndrome_o == 8'h83) ^ in[5];
	// Trace: design.sv:2861:3
	assign d_o[6] = (syndrome_o == 8'h0d) ^ in[6];
	// Trace: design.sv:2862:3
	assign d_o[7] = (syndrome_o == 8'h15) ^ in[7];
	// Trace: design.sv:2863:3
	assign d_o[8] = (syndrome_o == 8'h25) ^ in[8];
	// Trace: design.sv:2864:3
	assign d_o[9] = (syndrome_o == 8'h45) ^ in[9];
	// Trace: design.sv:2865:3
	assign d_o[10] = (syndrome_o == 8'h85) ^ in[10];
	// Trace: design.sv:2866:3
	assign d_o[11] = (syndrome_o == 8'h19) ^ in[11];
	// Trace: design.sv:2867:3
	assign d_o[12] = (syndrome_o == 8'h29) ^ in[12];
	// Trace: design.sv:2868:3
	assign d_o[13] = (syndrome_o == 8'h49) ^ in[13];
	// Trace: design.sv:2869:3
	assign d_o[14] = (syndrome_o == 8'h89) ^ in[14];
	// Trace: design.sv:2870:3
	assign d_o[15] = (syndrome_o == 8'h31) ^ in[15];
	// Trace: design.sv:2871:3
	assign d_o[16] = (syndrome_o == 8'h51) ^ in[16];
	// Trace: design.sv:2872:3
	assign d_o[17] = (syndrome_o == 8'h91) ^ in[17];
	// Trace: design.sv:2873:3
	assign d_o[18] = (syndrome_o == 8'h61) ^ in[18];
	// Trace: design.sv:2874:3
	assign d_o[19] = (syndrome_o == 8'ha1) ^ in[19];
	// Trace: design.sv:2875:3
	assign d_o[20] = (syndrome_o == 8'hc1) ^ in[20];
	// Trace: design.sv:2876:3
	assign d_o[21] = (syndrome_o == 8'h0e) ^ in[21];
	// Trace: design.sv:2877:3
	assign d_o[22] = (syndrome_o == 8'h16) ^ in[22];
	// Trace: design.sv:2878:3
	assign d_o[23] = (syndrome_o == 8'h26) ^ in[23];
	// Trace: design.sv:2879:3
	assign d_o[24] = (syndrome_o == 8'h46) ^ in[24];
	// Trace: design.sv:2880:3
	assign d_o[25] = (syndrome_o == 8'h86) ^ in[25];
	// Trace: design.sv:2881:3
	assign d_o[26] = (syndrome_o == 8'h1a) ^ in[26];
	// Trace: design.sv:2882:3
	assign d_o[27] = (syndrome_o == 8'h2a) ^ in[27];
	// Trace: design.sv:2883:3
	assign d_o[28] = (syndrome_o == 8'h4a) ^ in[28];
	// Trace: design.sv:2884:3
	assign d_o[29] = (syndrome_o == 8'h8a) ^ in[29];
	// Trace: design.sv:2885:3
	assign d_o[30] = (syndrome_o == 8'h32) ^ in[30];
	// Trace: design.sv:2886:3
	assign d_o[31] = (syndrome_o == 8'h52) ^ in[31];
	// Trace: design.sv:2887:3
	assign d_o[32] = (syndrome_o == 8'h92) ^ in[32];
	// Trace: design.sv:2888:3
	assign d_o[33] = (syndrome_o == 8'h62) ^ in[33];
	// Trace: design.sv:2889:3
	assign d_o[34] = (syndrome_o == 8'ha2) ^ in[34];
	// Trace: design.sv:2890:3
	assign d_o[35] = (syndrome_o == 8'hc2) ^ in[35];
	// Trace: design.sv:2891:3
	assign d_o[36] = (syndrome_o == 8'h1c) ^ in[36];
	// Trace: design.sv:2892:3
	assign d_o[37] = (syndrome_o == 8'h2c) ^ in[37];
	// Trace: design.sv:2893:3
	assign d_o[38] = (syndrome_o == 8'h4c) ^ in[38];
	// Trace: design.sv:2894:3
	assign d_o[39] = (syndrome_o == 8'h8c) ^ in[39];
	// Trace: design.sv:2895:3
	assign d_o[40] = (syndrome_o == 8'h34) ^ in[40];
	// Trace: design.sv:2896:3
	assign d_o[41] = (syndrome_o == 8'h54) ^ in[41];
	// Trace: design.sv:2897:3
	assign d_o[42] = (syndrome_o == 8'h94) ^ in[42];
	// Trace: design.sv:2898:3
	assign d_o[43] = (syndrome_o == 8'h64) ^ in[43];
	// Trace: design.sv:2899:3
	assign d_o[44] = (syndrome_o == 8'ha4) ^ in[44];
	// Trace: design.sv:2900:3
	assign d_o[45] = (syndrome_o == 8'hc4) ^ in[45];
	// Trace: design.sv:2901:3
	assign d_o[46] = (syndrome_o == 8'h38) ^ in[46];
	// Trace: design.sv:2902:3
	assign d_o[47] = (syndrome_o == 8'h58) ^ in[47];
	// Trace: design.sv:2903:3
	assign d_o[48] = (syndrome_o == 8'h98) ^ in[48];
	// Trace: design.sv:2904:3
	assign d_o[49] = (syndrome_o == 8'h68) ^ in[49];
	// Trace: design.sv:2905:3
	assign d_o[50] = (syndrome_o == 8'ha8) ^ in[50];
	// Trace: design.sv:2906:3
	assign d_o[51] = (syndrome_o == 8'hc8) ^ in[51];
	// Trace: design.sv:2907:3
	assign d_o[52] = (syndrome_o == 8'h70) ^ in[52];
	// Trace: design.sv:2908:3
	assign d_o[53] = (syndrome_o == 8'hb0) ^ in[53];
	// Trace: design.sv:2909:3
	assign d_o[54] = (syndrome_o == 8'hd0) ^ in[54];
	// Trace: design.sv:2910:3
	assign d_o[55] = (syndrome_o == 8'he0) ^ in[55];
	// Trace: design.sv:2911:3
	assign d_o[56] = (syndrome_o == 8'h6d) ^ in[56];
	// Trace: design.sv:2912:3
	assign d_o[57] = (syndrome_o == 8'hd6) ^ in[57];
	// Trace: design.sv:2913:3
	assign d_o[58] = (syndrome_o == 8'h3e) ^ in[58];
	// Trace: design.sv:2914:3
	assign d_o[59] = (syndrome_o == 8'hcb) ^ in[59];
	// Trace: design.sv:2915:3
	assign d_o[60] = (syndrome_o == 8'hb3) ^ in[60];
	// Trace: design.sv:2916:3
	assign d_o[61] = (syndrome_o == 8'hb5) ^ in[61];
	// Trace: design.sv:2917:3
	assign d_o[62] = (syndrome_o == 8'hce) ^ in[62];
	// Trace: design.sv:2918:3
	assign d_o[63] = (syndrome_o == 8'h79) ^ in[63];
	// Trace: design.sv:2921:3
	assign single_error = ^syndrome_o;
	// Trace: design.sv:2922:3
	assign err_o[0] = single_error;
	// Trace: design.sv:2923:3
	assign err_o[1] = ~single_error & |syndrome_o;
endmodule
module prim_secded_72_64_enc (
	in,
	out
);
	reg _sv2v_0;
	// Trace: design.sv:2933:3
	input [63:0] in;
	// Trace: design.sv:2934:3
	output reg [71:0] out;
	// Trace: design.sv:2937:3
	function automatic [71:0] sv2v_cast_72;
		input reg [71:0] inp;
		sv2v_cast_72 = inp;
	endfunction
	always @(*) begin : p_encode
		if (_sv2v_0)
			;
		// Trace: design.sv:2938:5
		out = sv2v_cast_72(in);
		// Trace: design.sv:2939:5
		out[64] = ^(out & 72'h00b9000000001fffff);
		// Trace: design.sv:2940:5
		out[65] = ^(out & 72'h005e00000fffe0003f);
		// Trace: design.sv:2941:5
		out[66] = ^(out & 72'h0067003ff003e007c1);
		// Trace: design.sv:2942:5
		out[67] = ^(out & 72'h00cd0fc0f03c207842);
		// Trace: design.sv:2943:5
		out[68] = ^(out & 72'h00b671c711c4438884);
		// Trace: design.sv:2944:5
		out[69] = ^(out & 72'h00b5b65926488c9108);
		// Trace: design.sv:2945:5
		out[70] = ^(out & 72'h00cbdaaa4a91152210);
		// Trace: design.sv:2946:5
		out[71] = ^(out & 72'h007aed348d221a4420);
	end
	initial _sv2v_0 = 0;
endmodule
module prim_secded_hamming_22_16_dec (
	in,
	d_o,
	syndrome_o,
	err_o
);
	// Trace: design.sv:2957:3
	input [21:0] in;
	// Trace: design.sv:2958:3
	output wire [15:0] d_o;
	// Trace: design.sv:2959:3
	output wire [5:0] syndrome_o;
	// Trace: design.sv:2960:3
	output wire [1:0] err_o;
	// Trace: design.sv:2965:3
	assign syndrome_o[0] = ^(in & 22'h01ad5b);
	// Trace: design.sv:2966:3
	assign syndrome_o[1] = ^(in & 22'h02366d);
	// Trace: design.sv:2967:3
	assign syndrome_o[2] = ^(in & 22'h04c78e);
	// Trace: design.sv:2968:3
	assign syndrome_o[3] = ^(in & 22'h0807f0);
	// Trace: design.sv:2969:3
	assign syndrome_o[4] = ^(in & 22'h10f800);
	// Trace: design.sv:2970:3
	assign syndrome_o[5] = ^(in & 22'h3fffff);
	// Trace: design.sv:2973:3
	assign d_o[0] = (syndrome_o == 6'h23) ^ in[0];
	// Trace: design.sv:2974:3
	assign d_o[1] = (syndrome_o == 6'h25) ^ in[1];
	// Trace: design.sv:2975:3
	assign d_o[2] = (syndrome_o == 6'h26) ^ in[2];
	// Trace: design.sv:2976:3
	assign d_o[3] = (syndrome_o == 6'h27) ^ in[3];
	// Trace: design.sv:2977:3
	assign d_o[4] = (syndrome_o == 6'h29) ^ in[4];
	// Trace: design.sv:2978:3
	assign d_o[5] = (syndrome_o == 6'h2a) ^ in[5];
	// Trace: design.sv:2979:3
	assign d_o[6] = (syndrome_o == 6'h2b) ^ in[6];
	// Trace: design.sv:2980:3
	assign d_o[7] = (syndrome_o == 6'h2c) ^ in[7];
	// Trace: design.sv:2981:3
	assign d_o[8] = (syndrome_o == 6'h2d) ^ in[8];
	// Trace: design.sv:2982:3
	assign d_o[9] = (syndrome_o == 6'h2e) ^ in[9];
	// Trace: design.sv:2983:3
	assign d_o[10] = (syndrome_o == 6'h2f) ^ in[10];
	// Trace: design.sv:2984:3
	assign d_o[11] = (syndrome_o == 6'h31) ^ in[11];
	// Trace: design.sv:2985:3
	assign d_o[12] = (syndrome_o == 6'h32) ^ in[12];
	// Trace: design.sv:2986:3
	assign d_o[13] = (syndrome_o == 6'h33) ^ in[13];
	// Trace: design.sv:2987:3
	assign d_o[14] = (syndrome_o == 6'h34) ^ in[14];
	// Trace: design.sv:2988:3
	assign d_o[15] = (syndrome_o == 6'h35) ^ in[15];
	// Trace: design.sv:2991:3
	assign err_o[0] = syndrome_o[5];
	// Trace: design.sv:2992:3
	assign err_o[1] = |syndrome_o[4:0] & ~syndrome_o[5];
endmodule
module prim_secded_hamming_22_16_enc (
	in,
	out
);
	reg _sv2v_0;
	// Trace: design.sv:3002:3
	input [15:0] in;
	// Trace: design.sv:3003:3
	output reg [21:0] out;
	// Trace: design.sv:3006:3
	function automatic [21:0] sv2v_cast_22;
		input reg [21:0] inp;
		sv2v_cast_22 = inp;
	endfunction
	always @(*) begin : p_encode
		if (_sv2v_0)
			;
		// Trace: design.sv:3007:5
		out = sv2v_cast_22(in);
		// Trace: design.sv:3008:5
		out[16] = ^(out & 22'h00ad5b);
		// Trace: design.sv:3009:5
		out[17] = ^(out & 22'h00366d);
		// Trace: design.sv:3010:5
		out[18] = ^(out & 22'h00c78e);
		// Trace: design.sv:3011:5
		out[19] = ^(out & 22'h0007f0);
		// Trace: design.sv:3012:5
		out[20] = ^(out & 22'h00f800);
		// Trace: design.sv:3013:5
		out[21] = ^(out & 22'h1fffff);
	end
	initial _sv2v_0 = 0;
endmodule
module prim_secded_hamming_39_32_dec (
	in,
	d_o,
	syndrome_o,
	err_o
);
	// Trace: design.sv:3024:3
	input [38:0] in;
	// Trace: design.sv:3025:3
	output wire [31:0] d_o;
	// Trace: design.sv:3026:3
	output wire [6:0] syndrome_o;
	// Trace: design.sv:3027:3
	output wire [1:0] err_o;
	// Trace: design.sv:3032:3
	assign syndrome_o[0] = ^(in & 39'h0156aaad5b);
	// Trace: design.sv:3033:3
	assign syndrome_o[1] = ^(in & 39'h029b33366d);
	// Trace: design.sv:3034:3
	assign syndrome_o[2] = ^(in & 39'h04e3c3c78e);
	// Trace: design.sv:3035:3
	assign syndrome_o[3] = ^(in & 39'h0803fc07f0);
	// Trace: design.sv:3036:3
	assign syndrome_o[4] = ^(in & 39'h1003fff800);
	// Trace: design.sv:3037:3
	assign syndrome_o[5] = ^(in & 39'h20fc000000);
	// Trace: design.sv:3038:3
	assign syndrome_o[6] = ^(in & 39'h7fffffffff);
	// Trace: design.sv:3041:3
	assign d_o[0] = (syndrome_o == 7'h43) ^ in[0];
	// Trace: design.sv:3042:3
	assign d_o[1] = (syndrome_o == 7'h45) ^ in[1];
	// Trace: design.sv:3043:3
	assign d_o[2] = (syndrome_o == 7'h46) ^ in[2];
	// Trace: design.sv:3044:3
	assign d_o[3] = (syndrome_o == 7'h47) ^ in[3];
	// Trace: design.sv:3045:3
	assign d_o[4] = (syndrome_o == 7'h49) ^ in[4];
	// Trace: design.sv:3046:3
	assign d_o[5] = (syndrome_o == 7'h4a) ^ in[5];
	// Trace: design.sv:3047:3
	assign d_o[6] = (syndrome_o == 7'h4b) ^ in[6];
	// Trace: design.sv:3048:3
	assign d_o[7] = (syndrome_o == 7'h4c) ^ in[7];
	// Trace: design.sv:3049:3
	assign d_o[8] = (syndrome_o == 7'h4d) ^ in[8];
	// Trace: design.sv:3050:3
	assign d_o[9] = (syndrome_o == 7'h4e) ^ in[9];
	// Trace: design.sv:3051:3
	assign d_o[10] = (syndrome_o == 7'h4f) ^ in[10];
	// Trace: design.sv:3052:3
	assign d_o[11] = (syndrome_o == 7'h51) ^ in[11];
	// Trace: design.sv:3053:3
	assign d_o[12] = (syndrome_o == 7'h52) ^ in[12];
	// Trace: design.sv:3054:3
	assign d_o[13] = (syndrome_o == 7'h53) ^ in[13];
	// Trace: design.sv:3055:3
	assign d_o[14] = (syndrome_o == 7'h54) ^ in[14];
	// Trace: design.sv:3056:3
	assign d_o[15] = (syndrome_o == 7'h55) ^ in[15];
	// Trace: design.sv:3057:3
	assign d_o[16] = (syndrome_o == 7'h56) ^ in[16];
	// Trace: design.sv:3058:3
	assign d_o[17] = (syndrome_o == 7'h57) ^ in[17];
	// Trace: design.sv:3059:3
	assign d_o[18] = (syndrome_o == 7'h58) ^ in[18];
	// Trace: design.sv:3060:3
	assign d_o[19] = (syndrome_o == 7'h59) ^ in[19];
	// Trace: design.sv:3061:3
	assign d_o[20] = (syndrome_o == 7'h5a) ^ in[20];
	// Trace: design.sv:3062:3
	assign d_o[21] = (syndrome_o == 7'h5b) ^ in[21];
	// Trace: design.sv:3063:3
	assign d_o[22] = (syndrome_o == 7'h5c) ^ in[22];
	// Trace: design.sv:3064:3
	assign d_o[23] = (syndrome_o == 7'h5d) ^ in[23];
	// Trace: design.sv:3065:3
	assign d_o[24] = (syndrome_o == 7'h5e) ^ in[24];
	// Trace: design.sv:3066:3
	assign d_o[25] = (syndrome_o == 7'h5f) ^ in[25];
	// Trace: design.sv:3067:3
	assign d_o[26] = (syndrome_o == 7'h61) ^ in[26];
	// Trace: design.sv:3068:3
	assign d_o[27] = (syndrome_o == 7'h62) ^ in[27];
	// Trace: design.sv:3069:3
	assign d_o[28] = (syndrome_o == 7'h63) ^ in[28];
	// Trace: design.sv:3070:3
	assign d_o[29] = (syndrome_o == 7'h64) ^ in[29];
	// Trace: design.sv:3071:3
	assign d_o[30] = (syndrome_o == 7'h65) ^ in[30];
	// Trace: design.sv:3072:3
	assign d_o[31] = (syndrome_o == 7'h66) ^ in[31];
	// Trace: design.sv:3075:3
	assign err_o[0] = syndrome_o[6];
	// Trace: design.sv:3076:3
	assign err_o[1] = |syndrome_o[5:0] & ~syndrome_o[6];
endmodule
module prim_secded_hamming_39_32_enc (
	in,
	out
);
	reg _sv2v_0;
	// Trace: design.sv:3086:3
	input [31:0] in;
	// Trace: design.sv:3087:3
	output reg [38:0] out;
	// Trace: design.sv:3090:3
	function automatic [38:0] sv2v_cast_39;
		input reg [38:0] inp;
		sv2v_cast_39 = inp;
	endfunction
	always @(*) begin : p_encode
		if (_sv2v_0)
			;
		// Trace: design.sv:3091:5
		out = sv2v_cast_39(in);
		// Trace: design.sv:3092:5
		out[32] = ^(out & 39'h0056aaad5b);
		// Trace: design.sv:3093:5
		out[33] = ^(out & 39'h009b33366d);
		// Trace: design.sv:3094:5
		out[34] = ^(out & 39'h00e3c3c78e);
		// Trace: design.sv:3095:5
		out[35] = ^(out & 39'h0003fc07f0);
		// Trace: design.sv:3096:5
		out[36] = ^(out & 39'h0003fff800);
		// Trace: design.sv:3097:5
		out[37] = ^(out & 39'h00fc000000);
		// Trace: design.sv:3098:5
		out[38] = ^(out & 39'h3fffffffff);
	end
	initial _sv2v_0 = 0;
endmodule
module prim_secded_hamming_72_64_dec (
	in,
	d_o,
	syndrome_o,
	err_o
);
	// Trace: design.sv:3109:3
	input [71:0] in;
	// Trace: design.sv:3110:3
	output wire [63:0] d_o;
	// Trace: design.sv:3111:3
	output wire [7:0] syndrome_o;
	// Trace: design.sv:3112:3
	output wire [1:0] err_o;
	// Trace: design.sv:3117:3
	assign syndrome_o[0] = ^(in & 72'h01ab55555556aaad5b);
	// Trace: design.sv:3118:3
	assign syndrome_o[1] = ^(in & 72'h02cd9999999b33366d);
	// Trace: design.sv:3119:3
	assign syndrome_o[2] = ^(in & 72'h04f1e1e1e1e3c3c78e);
	// Trace: design.sv:3120:3
	assign syndrome_o[3] = ^(in & 72'h0801fe01fe03fc07f0);
	// Trace: design.sv:3121:3
	assign syndrome_o[4] = ^(in & 72'h1001fffe0003fff800);
	// Trace: design.sv:3122:3
	assign syndrome_o[5] = ^(in & 72'h2001fffffffc000000);
	// Trace: design.sv:3123:3
	assign syndrome_o[6] = ^(in & 72'h40fe00000000000000);
	// Trace: design.sv:3124:3
	assign syndrome_o[7] = ^(in & 72'hffffffffffffffffff);
	// Trace: design.sv:3127:3
	assign d_o[0] = (syndrome_o == 8'h83) ^ in[0];
	// Trace: design.sv:3128:3
	assign d_o[1] = (syndrome_o == 8'h85) ^ in[1];
	// Trace: design.sv:3129:3
	assign d_o[2] = (syndrome_o == 8'h86) ^ in[2];
	// Trace: design.sv:3130:3
	assign d_o[3] = (syndrome_o == 8'h87) ^ in[3];
	// Trace: design.sv:3131:3
	assign d_o[4] = (syndrome_o == 8'h89) ^ in[4];
	// Trace: design.sv:3132:3
	assign d_o[5] = (syndrome_o == 8'h8a) ^ in[5];
	// Trace: design.sv:3133:3
	assign d_o[6] = (syndrome_o == 8'h8b) ^ in[6];
	// Trace: design.sv:3134:3
	assign d_o[7] = (syndrome_o == 8'h8c) ^ in[7];
	// Trace: design.sv:3135:3
	assign d_o[8] = (syndrome_o == 8'h8d) ^ in[8];
	// Trace: design.sv:3136:3
	assign d_o[9] = (syndrome_o == 8'h8e) ^ in[9];
	// Trace: design.sv:3137:3
	assign d_o[10] = (syndrome_o == 8'h8f) ^ in[10];
	// Trace: design.sv:3138:3
	assign d_o[11] = (syndrome_o == 8'h91) ^ in[11];
	// Trace: design.sv:3139:3
	assign d_o[12] = (syndrome_o == 8'h92) ^ in[12];
	// Trace: design.sv:3140:3
	assign d_o[13] = (syndrome_o == 8'h93) ^ in[13];
	// Trace: design.sv:3141:3
	assign d_o[14] = (syndrome_o == 8'h94) ^ in[14];
	// Trace: design.sv:3142:3
	assign d_o[15] = (syndrome_o == 8'h95) ^ in[15];
	// Trace: design.sv:3143:3
	assign d_o[16] = (syndrome_o == 8'h96) ^ in[16];
	// Trace: design.sv:3144:3
	assign d_o[17] = (syndrome_o == 8'h97) ^ in[17];
	// Trace: design.sv:3145:3
	assign d_o[18] = (syndrome_o == 8'h98) ^ in[18];
	// Trace: design.sv:3146:3
	assign d_o[19] = (syndrome_o == 8'h99) ^ in[19];
	// Trace: design.sv:3147:3
	assign d_o[20] = (syndrome_o == 8'h9a) ^ in[20];
	// Trace: design.sv:3148:3
	assign d_o[21] = (syndrome_o == 8'h9b) ^ in[21];
	// Trace: design.sv:3149:3
	assign d_o[22] = (syndrome_o == 8'h9c) ^ in[22];
	// Trace: design.sv:3150:3
	assign d_o[23] = (syndrome_o == 8'h9d) ^ in[23];
	// Trace: design.sv:3151:3
	assign d_o[24] = (syndrome_o == 8'h9e) ^ in[24];
	// Trace: design.sv:3152:3
	assign d_o[25] = (syndrome_o == 8'h9f) ^ in[25];
	// Trace: design.sv:3153:3
	assign d_o[26] = (syndrome_o == 8'ha1) ^ in[26];
	// Trace: design.sv:3154:3
	assign d_o[27] = (syndrome_o == 8'ha2) ^ in[27];
	// Trace: design.sv:3155:3
	assign d_o[28] = (syndrome_o == 8'ha3) ^ in[28];
	// Trace: design.sv:3156:3
	assign d_o[29] = (syndrome_o == 8'ha4) ^ in[29];
	// Trace: design.sv:3157:3
	assign d_o[30] = (syndrome_o == 8'ha5) ^ in[30];
	// Trace: design.sv:3158:3
	assign d_o[31] = (syndrome_o == 8'ha6) ^ in[31];
	// Trace: design.sv:3159:3
	assign d_o[32] = (syndrome_o == 8'ha7) ^ in[32];
	// Trace: design.sv:3160:3
	assign d_o[33] = (syndrome_o == 8'ha8) ^ in[33];
	// Trace: design.sv:3161:3
	assign d_o[34] = (syndrome_o == 8'ha9) ^ in[34];
	// Trace: design.sv:3162:3
	assign d_o[35] = (syndrome_o == 8'haa) ^ in[35];
	// Trace: design.sv:3163:3
	assign d_o[36] = (syndrome_o == 8'hab) ^ in[36];
	// Trace: design.sv:3164:3
	assign d_o[37] = (syndrome_o == 8'hac) ^ in[37];
	// Trace: design.sv:3165:3
	assign d_o[38] = (syndrome_o == 8'had) ^ in[38];
	// Trace: design.sv:3166:3
	assign d_o[39] = (syndrome_o == 8'hae) ^ in[39];
	// Trace: design.sv:3167:3
	assign d_o[40] = (syndrome_o == 8'haf) ^ in[40];
	// Trace: design.sv:3168:3
	assign d_o[41] = (syndrome_o == 8'hb0) ^ in[41];
	// Trace: design.sv:3169:3
	assign d_o[42] = (syndrome_o == 8'hb1) ^ in[42];
	// Trace: design.sv:3170:3
	assign d_o[43] = (syndrome_o == 8'hb2) ^ in[43];
	// Trace: design.sv:3171:3
	assign d_o[44] = (syndrome_o == 8'hb3) ^ in[44];
	// Trace: design.sv:3172:3
	assign d_o[45] = (syndrome_o == 8'hb4) ^ in[45];
	// Trace: design.sv:3173:3
	assign d_o[46] = (syndrome_o == 8'hb5) ^ in[46];
	// Trace: design.sv:3174:3
	assign d_o[47] = (syndrome_o == 8'hb6) ^ in[47];
	// Trace: design.sv:3175:3
	assign d_o[48] = (syndrome_o == 8'hb7) ^ in[48];
	// Trace: design.sv:3176:3
	assign d_o[49] = (syndrome_o == 8'hb8) ^ in[49];
	// Trace: design.sv:3177:3
	assign d_o[50] = (syndrome_o == 8'hb9) ^ in[50];
	// Trace: design.sv:3178:3
	assign d_o[51] = (syndrome_o == 8'hba) ^ in[51];
	// Trace: design.sv:3179:3
	assign d_o[52] = (syndrome_o == 8'hbb) ^ in[52];
	// Trace: design.sv:3180:3
	assign d_o[53] = (syndrome_o == 8'hbc) ^ in[53];
	// Trace: design.sv:3181:3
	assign d_o[54] = (syndrome_o == 8'hbd) ^ in[54];
	// Trace: design.sv:3182:3
	assign d_o[55] = (syndrome_o == 8'hbe) ^ in[55];
	// Trace: design.sv:3183:3
	assign d_o[56] = (syndrome_o == 8'hbf) ^ in[56];
	// Trace: design.sv:3184:3
	assign d_o[57] = (syndrome_o == 8'hc1) ^ in[57];
	// Trace: design.sv:3185:3
	assign d_o[58] = (syndrome_o == 8'hc2) ^ in[58];
	// Trace: design.sv:3186:3
	assign d_o[59] = (syndrome_o == 8'hc3) ^ in[59];
	// Trace: design.sv:3187:3
	assign d_o[60] = (syndrome_o == 8'hc4) ^ in[60];
	// Trace: design.sv:3188:3
	assign d_o[61] = (syndrome_o == 8'hc5) ^ in[61];
	// Trace: design.sv:3189:3
	assign d_o[62] = (syndrome_o == 8'hc6) ^ in[62];
	// Trace: design.sv:3190:3
	assign d_o[63] = (syndrome_o == 8'hc7) ^ in[63];
	// Trace: design.sv:3193:3
	assign err_o[0] = syndrome_o[7];
	// Trace: design.sv:3194:3
	assign err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
endmodule
module prim_secded_hamming_72_64_enc (
	in,
	out
);
	reg _sv2v_0;
	// Trace: design.sv:3204:3
	input [63:0] in;
	// Trace: design.sv:3205:3
	output reg [71:0] out;
	// Trace: design.sv:3208:3
	function automatic [71:0] sv2v_cast_72;
		input reg [71:0] inp;
		sv2v_cast_72 = inp;
	endfunction
	always @(*) begin : p_encode
		if (_sv2v_0)
			;
		// Trace: design.sv:3209:5
		out = sv2v_cast_72(in);
		// Trace: design.sv:3210:5
		out[64] = ^(out & 72'h00ab55555556aaad5b);
		// Trace: design.sv:3211:5
		out[65] = ^(out & 72'h00cd9999999b33366d);
		// Trace: design.sv:3212:5
		out[66] = ^(out & 72'h00f1e1e1e1e3c3c78e);
		// Trace: design.sv:3213:5
		out[67] = ^(out & 72'h0001fe01fe03fc07f0);
		// Trace: design.sv:3214:5
		out[68] = ^(out & 72'h0001fffe0003fff800);
		// Trace: design.sv:3215:5
		out[69] = ^(out & 72'h0001fffffffc000000);
		// Trace: design.sv:3216:5
		out[70] = ^(out & 72'h00fe00000000000000);
		// Trace: design.sv:3217:5
		out[71] = ^(out & 72'h7fffffffffffffffff);
	end
	initial _sv2v_0 = 0;
endmodule
module prim_subreg_arb (
	we,
	wd,
	de,
	d,
	q,
	wr_en,
	wr_data
);
	// Trace: design.sv:3228:13
	parameter signed [31:0] DW = 32;
	// Trace: design.sv:3229:17
	parameter SWACCESS = "RW";
	// Trace: design.sv:3233:3
	input we;
	// Trace: design.sv:3234:3
	input [DW - 1:0] wd;
	// Trace: design.sv:3237:3
	input de;
	// Trace: design.sv:3238:3
	input [DW - 1:0] d;
	// Trace: design.sv:3241:3
	input [DW - 1:0] q;
	// Trace: design.sv:3244:3
	output wire wr_en;
	// Trace: design.sv:3245:3
	output wire [DW - 1:0] wr_data;
	// Trace: design.sv:3248:3
	generate
		if ((SWACCESS == "RW") || (SWACCESS == "WO")) begin : gen_w
			// Trace: design.sv:3249:5
			assign wr_en = we | de;
			// Trace: design.sv:3250:5
			assign wr_data = (we == 1'b1 ? wd : d);
			// Trace: design.sv:3252:5
			wire [DW - 1:0] unused_q;
			// Trace: design.sv:3253:5
			assign unused_q = q;
		end
		else if (SWACCESS == "RO") begin : gen_ro
			// Trace: design.sv:3255:5
			assign wr_en = de;
			// Trace: design.sv:3256:5
			assign wr_data = d;
			// Trace: design.sv:3258:5
			wire unused_we;
			// Trace: design.sv:3259:5
			wire [DW - 1:0] unused_wd;
			// Trace: design.sv:3260:5
			wire [DW - 1:0] unused_q;
			// Trace: design.sv:3261:5
			assign unused_we = we;
			// Trace: design.sv:3262:5
			assign unused_wd = wd;
			// Trace: design.sv:3263:5
			assign unused_q = q;
		end
		else if (SWACCESS == "W1S") begin : gen_w1s
			// Trace: design.sv:3268:5
			assign wr_en = we | de;
			// Trace: design.sv:3269:5
			assign wr_data = (de ? d : q) | (we ? wd : {DW {1'sb0}});
		end
		else if (SWACCESS == "W1C") begin : gen_w1c
			// Trace: design.sv:3274:5
			assign wr_en = we | de;
			// Trace: design.sv:3275:5
			assign wr_data = (de ? d : q) & (we ? ~wd : {DW {1'sb1}});
		end
		else if (SWACCESS == "W0C") begin : gen_w0c
			// Trace: design.sv:3277:5
			assign wr_en = we | de;
			// Trace: design.sv:3278:5
			assign wr_data = (de ? d : q) & (we ? wd : {DW {1'sb1}});
		end
		else if (SWACCESS == "RC") begin : gen_rc
			// Trace: design.sv:3282:5
			assign wr_en = we | de;
			// Trace: design.sv:3283:5
			assign wr_data = (de ? d : q) & (we ? {DW {1'sb0}} : {DW {1'sb1}});
			// Trace: design.sv:3285:5
			wire [DW - 1:0] unused_wd;
			// Trace: design.sv:3286:5
			assign unused_wd = wd;
		end
		else begin : gen_hw
			// Trace: design.sv:3288:5
			assign wr_en = de;
			// Trace: design.sv:3289:5
			assign wr_data = d;
			// Trace: design.sv:3291:5
			wire unused_we;
			// Trace: design.sv:3292:5
			wire [DW - 1:0] unused_wd;
			// Trace: design.sv:3293:5
			wire [DW - 1:0] unused_q;
			// Trace: design.sv:3294:5
			assign unused_we = we;
			// Trace: design.sv:3295:5
			assign unused_wd = wd;
			// Trace: design.sv:3296:5
			assign unused_q = q;
		end
	endgenerate
endmodule
module prim_subreg (
	clk_i,
	rst_ni,
	we,
	wd,
	de,
	d,
	qe,
	q,
	qs
);
	// Trace: design.sv:3307:13
	parameter signed [31:0] DW = 32;
	// Trace: design.sv:3308:28
	parameter SWACCESS = "RW";
	// Trace: design.sv:3309:13
	parameter [DW - 1:0] RESVAL = 1'sb0;
	// Trace: design.sv:3311:3
	input clk_i;
	// Trace: design.sv:3312:3
	input rst_ni;
	// Trace: design.sv:3316:3
	input we;
	// Trace: design.sv:3317:3
	input [DW - 1:0] wd;
	// Trace: design.sv:3320:3
	input de;
	// Trace: design.sv:3321:3
	input [DW - 1:0] d;
	// Trace: design.sv:3324:3
	output reg qe;
	// Trace: design.sv:3325:3
	output reg [DW - 1:0] q;
	// Trace: design.sv:3326:3
	output wire [DW - 1:0] qs;
	// Trace: design.sv:3329:3
	wire wr_en;
	// Trace: design.sv:3330:3
	wire [DW - 1:0] wr_data;
	// Trace: design.sv:3332:3
	prim_subreg_arb #(
		.DW(DW),
		.SWACCESS(SWACCESS)
	) wr_en_data_arb(
		.we(we),
		.wd(wd),
		.de(de),
		.d(d),
		.q(q),
		.wr_en(wr_en),
		.wr_data(wr_data)
	);
	// Trace: design.sv:3345:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:3346:5
		if (!rst_ni)
			// Trace: design.sv:3347:7
			qe <= 1'b0;
		else
			// Trace: design.sv:3349:7
			qe <= we;
	// Trace: design.sv:3353:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:3354:5
		if (!rst_ni)
			// Trace: design.sv:3355:7
			q <= RESVAL;
		else if (wr_en)
			// Trace: design.sv:3357:7
			q <= wr_data;
	// Trace: design.sv:3361:3
	assign qs = q;
endmodule
module prim_subreg_ext (
	re,
	we,
	wd,
	d,
	qe,
	qre,
	q,
	qs
);
	// Trace: design.sv:3371:13
	parameter [31:0] DW = 32;
	// Trace: design.sv:3373:3
	input re;
	// Trace: design.sv:3374:3
	input we;
	// Trace: design.sv:3375:3
	input [DW - 1:0] wd;
	// Trace: design.sv:3377:3
	input [DW - 1:0] d;
	// Trace: design.sv:3380:3
	output wire qe;
	// Trace: design.sv:3381:3
	output wire qre;
	// Trace: design.sv:3382:3
	output wire [DW - 1:0] q;
	// Trace: design.sv:3383:3
	output wire [DW - 1:0] qs;
	// Trace: design.sv:3386:3
	assign qs = d;
	// Trace: design.sv:3387:3
	assign q = wd;
	// Trace: design.sv:3388:3
	assign qe = we;
	// Trace: design.sv:3389:3
	assign qre = re;
endmodule
module prim_subreg_shadow (
	clk_i,
	rst_ni,
	re,
	we,
	wd,
	de,
	d,
	qe,
	q,
	qs,
	err_update,
	err_storage
);
	// Trace: design.sv:3399:13
	parameter signed [31:0] DW = 32;
	// Trace: design.sv:3400:28
	parameter SWACCESS = "RW";
	// Trace: design.sv:3401:13
	parameter [DW - 1:0] RESVAL = 1'sb0;
	// Trace: design.sv:3403:3
	input clk_i;
	// Trace: design.sv:3404:3
	input rst_ni;
	// Trace: design.sv:3408:3
	input re;
	// Trace: design.sv:3410:3
	input we;
	// Trace: design.sv:3411:3
	input [DW - 1:0] wd;
	// Trace: design.sv:3414:3
	input de;
	// Trace: design.sv:3415:3
	input [DW - 1:0] d;
	// Trace: design.sv:3418:3
	output wire qe;
	// Trace: design.sv:3419:3
	output wire [DW - 1:0] q;
	// Trace: design.sv:3420:3
	output wire [DW - 1:0] qs;
	// Trace: design.sv:3423:3
	output wire err_update;
	// Trace: design.sv:3424:3
	output wire err_storage;
	// Trace: design.sv:3428:3
	wire phase_clear;
	// Trace: design.sv:3429:3
	reg phase_q;
	// Trace: design.sv:3430:3
	wire staged_we;
	wire shadow_we;
	wire committed_we;
	// Trace: design.sv:3431:3
	wire staged_de;
	wire shadow_de;
	wire committed_de;
	// Trace: design.sv:3434:3
	wire staged_qe;
	wire shadow_qe;
	wire committed_qe;
	// Trace: design.sv:3435:3
	wire [DW - 1:0] staged_q;
	wire [DW - 1:0] shadow_q;
	wire [DW - 1:0] committed_q;
	// Trace: design.sv:3436:3
	wire [DW - 1:0] committed_qs;
	// Trace: design.sv:3440:3
	wire wr_en;
	// Trace: design.sv:3441:3
	wire [DW - 1:0] wr_data;
	// Trace: design.sv:3443:3
	prim_subreg_arb #(
		.DW(DW),
		.SWACCESS(SWACCESS)
	) wr_en_data_arb(
		.we(we),
		.wd(wd),
		.de(de),
		.d(d),
		.q(q),
		.wr_en(wr_en),
		.wr_data(wr_data)
	);
	// Trace: design.sv:3459:3
	assign phase_clear = (SWACCESS == "RO" ? 1'b0 : re);
	// Trace: design.sv:3464:3
	always @(posedge clk_i or negedge rst_ni) begin : phase_reg
		// Trace: design.sv:3465:5
		if (!rst_ni)
			// Trace: design.sv:3466:7
			phase_q <= 1'b0;
		else if (wr_en)
			// Trace: design.sv:3468:7
			phase_q <= ~phase_q;
		else if (phase_clear)
			// Trace: design.sv:3470:7
			phase_q <= 1'b0;
	end
	// Trace: design.sv:3477:3
	assign staged_we = we & ~phase_q;
	// Trace: design.sv:3478:3
	assign staged_de = de & ~phase_q;
	// Trace: design.sv:3479:3
	prim_subreg #(
		.DW(DW),
		.SWACCESS(SWACCESS),
		.RESVAL(~RESVAL)
	) staged_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(staged_we),
		.wd(~wd),
		.de(staged_de),
		.d(~d),
		.qe(staged_qe),
		.q(staged_q),
		.qs()
	);
	// Trace: design.sv:3500:3
	assign shadow_we = (we & phase_q) & ~err_update;
	// Trace: design.sv:3501:3
	assign shadow_de = (de & phase_q) & ~err_update;
	// Trace: design.sv:3502:3
	prim_subreg #(
		.DW(DW),
		.SWACCESS(SWACCESS),
		.RESVAL(~RESVAL)
	) shadow_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(shadow_we),
		.wd(staged_q),
		.de(shadow_de),
		.d(staged_q),
		.qe(shadow_qe),
		.q(shadow_q),
		.qs()
	);
	// Trace: design.sv:3521:3
	assign committed_we = shadow_we;
	// Trace: design.sv:3522:3
	assign committed_de = shadow_de;
	// Trace: design.sv:3523:3
	prim_subreg #(
		.DW(DW),
		.SWACCESS(SWACCESS),
		.RESVAL(RESVAL)
	) committed_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(committed_we),
		.wd(wd),
		.de(committed_de),
		.d(d),
		.qe(committed_qe),
		.q(committed_q),
		.qs(committed_qs)
	);
	// Trace: design.sv:3540:3
	assign err_update = (~staged_q != wr_data ? phase_q & wr_en : 1'b0);
	// Trace: design.sv:3541:3
	assign err_storage = ~shadow_q != committed_q;
	// Trace: design.sv:3544:3
	assign qe = (staged_qe | shadow_qe) | committed_qe;
	// Trace: design.sv:3545:3
	assign q = committed_q;
	// Trace: design.sv:3546:3
	assign qs = committed_qs;
endmodule
// removed package "prim_util_pkg"
// removed package "cv32e40p_apu_core_pkg"
// removed package "cv32e40p_fpu_pkg"
// removed package "cv32e40p_pkg"
module cv32e40p_alu (
	clk,
	rst_n,
	enable_i,
	operator_i,
	operand_a_i,
	operand_b_i,
	operand_c_i,
	vector_mode_i,
	bmask_a_i,
	bmask_b_i,
	imm_vec_ext_i,
	is_clpx_i,
	is_subrot_i,
	clpx_shift_i,
	result_o,
	comparison_result_o,
	ready_o,
	ex_ready_i
);
	reg _sv2v_0;
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:4581:5
	input wire clk;
	// Trace: design.sv:4582:5
	input wire rst_n;
	// Trace: design.sv:4583:5
	input wire enable_i;
	// Trace: design.sv:4584:5
	localparam cv32e40p_pkg_ALU_OP_WIDTH = 7;
	// removed localparam type cv32e40p_pkg_alu_opcode_e
	input wire [6:0] operator_i;
	// Trace: design.sv:4585:5
	input wire [31:0] operand_a_i;
	// Trace: design.sv:4586:5
	input wire [31:0] operand_b_i;
	// Trace: design.sv:4587:5
	input wire [31:0] operand_c_i;
	// Trace: design.sv:4589:5
	input wire [1:0] vector_mode_i;
	// Trace: design.sv:4590:5
	input wire [4:0] bmask_a_i;
	// Trace: design.sv:4591:5
	input wire [4:0] bmask_b_i;
	// Trace: design.sv:4592:5
	input wire [1:0] imm_vec_ext_i;
	// Trace: design.sv:4594:5
	input wire is_clpx_i;
	// Trace: design.sv:4595:5
	input wire is_subrot_i;
	// Trace: design.sv:4596:5
	input wire [1:0] clpx_shift_i;
	// Trace: design.sv:4598:5
	output reg [31:0] result_o;
	// Trace: design.sv:4599:5
	output wire comparison_result_o;
	// Trace: design.sv:4601:5
	output wire ready_o;
	// Trace: design.sv:4602:5
	input wire ex_ready_i;
	// Trace: design.sv:4605:3
	wire [31:0] operand_a_rev;
	// Trace: design.sv:4606:3
	wire [31:0] operand_a_neg;
	// Trace: design.sv:4607:3
	wire [31:0] operand_a_neg_rev;
	// Trace: design.sv:4609:3
	assign operand_a_neg = ~operand_a_i;
	// Trace: design.sv:4612:3
	// Trace: design.sv:4613:5
	genvar _gv_k_1;
	generate
		for (_gv_k_1 = 0; _gv_k_1 < 32; _gv_k_1 = _gv_k_1 + 1) begin : gen_operand_a_rev
			localparam k = _gv_k_1;
			// Trace: design.sv:4615:7
			assign operand_a_rev[k] = operand_a_i[31 - k];
		end
	endgenerate
	// Trace: design.sv:4620:3
	// Trace: design.sv:4621:5
	genvar _gv_m_1;
	generate
		for (_gv_m_1 = 0; _gv_m_1 < 32; _gv_m_1 = _gv_m_1 + 1) begin : gen_operand_a_neg_rev
			localparam m = _gv_m_1;
			// Trace: design.sv:4623:7
			assign operand_a_neg_rev[m] = operand_a_neg[31 - m];
		end
	endgenerate
	// Trace: design.sv:4627:3
	wire [31:0] operand_b_neg;
	// Trace: design.sv:4629:3
	assign operand_b_neg = ~operand_b_i;
	// Trace: design.sv:4632:3
	wire [5:0] div_shift;
	// Trace: design.sv:4633:3
	wire div_valid;
	// Trace: design.sv:4634:3
	wire [31:0] bmask;
	// Trace: design.sv:4645:3
	wire adder_op_b_negate;
	// Trace: design.sv:4646:3
	wire [31:0] adder_op_a;
	wire [31:0] adder_op_b;
	// Trace: design.sv:4647:3
	reg [35:0] adder_in_a;
	reg [35:0] adder_in_b;
	// Trace: design.sv:4648:3
	wire [31:0] adder_result;
	// Trace: design.sv:4649:3
	wire [36:0] adder_result_expanded;
	// Trace: design.sv:4652:3
	function automatic [6:0] sv2v_cast_C07C4;
		input reg [6:0] inp;
		sv2v_cast_C07C4 = inp;
	endfunction
	assign adder_op_b_negate = ((((operator_i == sv2v_cast_C07C4(7'b0011001)) || (operator_i == sv2v_cast_C07C4(7'b0011101))) || (operator_i == sv2v_cast_C07C4(7'b0011011))) || (operator_i == sv2v_cast_C07C4(7'b0011111))) || is_subrot_i;
	// Trace: design.sv:4656:3
	assign adder_op_a = (operator_i == sv2v_cast_C07C4(7'b0010100) ? operand_a_neg : (is_subrot_i ? {operand_b_i[15:0], operand_a_i[31:16]} : operand_a_i));
	// Trace: design.sv:4661:3
	assign adder_op_b = (adder_op_b_negate ? (is_subrot_i ? ~{operand_a_i[15:0], operand_b_i[31:16]} : operand_b_neg) : operand_b_i);
	// Trace: design.sv:4666:3
	localparam cv32e40p_pkg_VEC_MODE16 = 2'b10;
	localparam cv32e40p_pkg_VEC_MODE8 = 2'b11;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:4667:5
		adder_in_a[0] = 1'b1;
		// Trace: design.sv:4668:5
		adder_in_a[8:1] = adder_op_a[7:0];
		// Trace: design.sv:4669:5
		adder_in_a[9] = 1'b1;
		// Trace: design.sv:4670:5
		adder_in_a[17:10] = adder_op_a[15:8];
		// Trace: design.sv:4671:5
		adder_in_a[18] = 1'b1;
		// Trace: design.sv:4672:5
		adder_in_a[26:19] = adder_op_a[23:16];
		// Trace: design.sv:4673:5
		adder_in_a[27] = 1'b1;
		// Trace: design.sv:4674:5
		adder_in_a[35:28] = adder_op_a[31:24];
		// Trace: design.sv:4676:5
		adder_in_b[0] = 1'b0;
		// Trace: design.sv:4677:5
		adder_in_b[8:1] = adder_op_b[7:0];
		// Trace: design.sv:4678:5
		adder_in_b[9] = 1'b0;
		// Trace: design.sv:4679:5
		adder_in_b[17:10] = adder_op_b[15:8];
		// Trace: design.sv:4680:5
		adder_in_b[18] = 1'b0;
		// Trace: design.sv:4681:5
		adder_in_b[26:19] = adder_op_b[23:16];
		// Trace: design.sv:4682:5
		adder_in_b[27] = 1'b0;
		// Trace: design.sv:4683:5
		adder_in_b[35:28] = adder_op_b[31:24];
		// Trace: design.sv:4685:5
		if (adder_op_b_negate || ((operator_i == sv2v_cast_C07C4(7'b0010100)) || (operator_i == sv2v_cast_C07C4(7'b0010110)))) begin
			// Trace: design.sv:4687:7
			adder_in_b[0] = 1'b1;
			// Trace: design.sv:4689:7
			case (vector_mode_i)
				cv32e40p_pkg_VEC_MODE16:
					// Trace: design.sv:4691:11
					adder_in_b[18] = 1'b1;
				cv32e40p_pkg_VEC_MODE8: begin
					// Trace: design.sv:4695:11
					adder_in_b[9] = 1'b1;
					// Trace: design.sv:4696:11
					adder_in_b[18] = 1'b1;
					// Trace: design.sv:4697:11
					adder_in_b[27] = 1'b1;
				end
			endcase
		end
		else
			// Trace: design.sv:4703:7
			case (vector_mode_i)
				cv32e40p_pkg_VEC_MODE16:
					// Trace: design.sv:4705:11
					adder_in_a[18] = 1'b0;
				cv32e40p_pkg_VEC_MODE8: begin
					// Trace: design.sv:4709:11
					adder_in_a[9] = 1'b0;
					// Trace: design.sv:4710:11
					adder_in_a[18] = 1'b0;
					// Trace: design.sv:4711:11
					adder_in_a[27] = 1'b0;
				end
			endcase
	end
	// Trace: design.sv:4718:3
	assign adder_result_expanded = $signed(adder_in_a) + $signed(adder_in_b);
	// Trace: design.sv:4719:3
	assign adder_result = {adder_result_expanded[35:28], adder_result_expanded[26:19], adder_result_expanded[17:10], adder_result_expanded[8:1]};
	// Trace: design.sv:4728:3
	wire [31:0] adder_round_value;
	// Trace: design.sv:4729:3
	wire [31:0] adder_round_result;
	// Trace: design.sv:4731:3
	assign adder_round_value = ((((operator_i == sv2v_cast_C07C4(7'b0011100)) || (operator_i == sv2v_cast_C07C4(7'b0011101))) || (operator_i == sv2v_cast_C07C4(7'b0011110))) || (operator_i == sv2v_cast_C07C4(7'b0011111)) ? {1'b0, bmask[31:1]} : {32 {1'sb0}});
	// Trace: design.sv:4736:3
	assign adder_round_result = adder_result + adder_round_value;
	// Trace: design.sv:4748:3
	wire shift_left;
	// Trace: design.sv:4749:3
	wire shift_use_round;
	// Trace: design.sv:4750:3
	wire shift_arithmetic;
	// Trace: design.sv:4752:3
	reg [31:0] shift_amt_left;
	// Trace: design.sv:4753:3
	wire [31:0] shift_amt;
	// Trace: design.sv:4754:3
	wire [31:0] shift_amt_int;
	// Trace: design.sv:4755:3
	wire [31:0] shift_amt_norm;
	// Trace: design.sv:4756:3
	wire [31:0] shift_op_a;
	// Trace: design.sv:4757:3
	wire [31:0] shift_result;
	// Trace: design.sv:4758:3
	reg [31:0] shift_right_result;
	// Trace: design.sv:4759:3
	wire [31:0] shift_left_result;
	// Trace: design.sv:4760:3
	wire [15:0] clpx_shift_ex;
	// Trace: design.sv:4763:3
	assign shift_amt = (div_valid ? div_shift : operand_b_i);
	// Trace: design.sv:4766:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:4767:5
		case (vector_mode_i)
			cv32e40p_pkg_VEC_MODE16: begin
				// Trace: design.sv:4769:9
				shift_amt_left[15:0] = shift_amt[31:16];
				// Trace: design.sv:4770:9
				shift_amt_left[31:16] = shift_amt[15:0];
			end
			cv32e40p_pkg_VEC_MODE8: begin
				// Trace: design.sv:4774:9
				shift_amt_left[7:0] = shift_amt[31:24];
				// Trace: design.sv:4775:9
				shift_amt_left[15:8] = shift_amt[23:16];
				// Trace: design.sv:4776:9
				shift_amt_left[23:16] = shift_amt[15:8];
				// Trace: design.sv:4777:9
				shift_amt_left[31:24] = shift_amt[7:0];
			end
			default:
				// Trace: design.sv:4782:9
				shift_amt_left[31:0] = shift_amt[31:0];
		endcase
	end
	// Trace: design.sv:4788:3
	assign shift_left = ((((((((operator_i == sv2v_cast_C07C4(7'b0100111)) || (operator_i == sv2v_cast_C07C4(7'b0101010))) || (operator_i == sv2v_cast_C07C4(7'b0110111))) || (operator_i == sv2v_cast_C07C4(7'b0110101))) || (operator_i == sv2v_cast_C07C4(7'b0110001))) || (operator_i == sv2v_cast_C07C4(7'b0110000))) || (operator_i == sv2v_cast_C07C4(7'b0110011))) || (operator_i == sv2v_cast_C07C4(7'b0110010))) || (operator_i == sv2v_cast_C07C4(7'b1001001));
	// Trace: design.sv:4794:3
	assign shift_use_round = (((((((operator_i == sv2v_cast_C07C4(7'b0011000)) || (operator_i == sv2v_cast_C07C4(7'b0011001))) || (operator_i == sv2v_cast_C07C4(7'b0011100))) || (operator_i == sv2v_cast_C07C4(7'b0011101))) || (operator_i == sv2v_cast_C07C4(7'b0011010))) || (operator_i == sv2v_cast_C07C4(7'b0011011))) || (operator_i == sv2v_cast_C07C4(7'b0011110))) || (operator_i == sv2v_cast_C07C4(7'b0011111));
	// Trace: design.sv:4799:3
	assign shift_arithmetic = (((((operator_i == sv2v_cast_C07C4(7'b0100100)) || (operator_i == sv2v_cast_C07C4(7'b0101000))) || (operator_i == sv2v_cast_C07C4(7'b0011000))) || (operator_i == sv2v_cast_C07C4(7'b0011001))) || (operator_i == sv2v_cast_C07C4(7'b0011100))) || (operator_i == sv2v_cast_C07C4(7'b0011101));
	// Trace: design.sv:4804:3
	assign shift_op_a = (shift_left ? operand_a_rev : (shift_use_round ? adder_round_result : operand_a_i));
	// Trace: design.sv:4806:3
	assign shift_amt_int = (shift_use_round ? shift_amt_norm : (shift_left ? shift_amt_left : shift_amt));
	// Trace: design.sv:4809:3
	assign shift_amt_norm = (is_clpx_i ? {clpx_shift_ex, clpx_shift_ex} : {4 {3'b000, bmask_b_i}});
	// Trace: design.sv:4811:3
	assign clpx_shift_ex = $unsigned(clpx_shift_i);
	// Trace: design.sv:4814:3
	wire [63:0] shift_op_a_32;
	// Trace: design.sv:4816:3
	assign shift_op_a_32 = (operator_i == sv2v_cast_C07C4(7'b0100110) ? {shift_op_a, shift_op_a} : $signed({{32 {shift_arithmetic & shift_op_a[31]}}, shift_op_a}));
	// Trace: design.sv:4822:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:4823:5
		case (vector_mode_i)
			cv32e40p_pkg_VEC_MODE16: begin
				// Trace: design.sv:4825:9
				shift_right_result[31:16] = $signed({shift_arithmetic & shift_op_a[31], shift_op_a[31:16]}) >>> shift_amt_int[19:16];
				// Trace: design.sv:4828:9
				shift_right_result[15:0] = $signed({shift_arithmetic & shift_op_a[15], shift_op_a[15:0]}) >>> shift_amt_int[3:0];
			end
			cv32e40p_pkg_VEC_MODE8: begin
				// Trace: design.sv:4834:9
				shift_right_result[31:24] = $signed({shift_arithmetic & shift_op_a[31], shift_op_a[31:24]}) >>> shift_amt_int[26:24];
				// Trace: design.sv:4837:9
				shift_right_result[23:16] = $signed({shift_arithmetic & shift_op_a[23], shift_op_a[23:16]}) >>> shift_amt_int[18:16];
				// Trace: design.sv:4840:9
				shift_right_result[15:8] = $signed({shift_arithmetic & shift_op_a[15], shift_op_a[15:8]}) >>> shift_amt_int[10:8];
				// Trace: design.sv:4843:9
				shift_right_result[7:0] = $signed({shift_arithmetic & shift_op_a[7], shift_op_a[7:0]}) >>> shift_amt_int[2:0];
			end
			default:
				// Trace: design.sv:4850:9
				shift_right_result = shift_op_a_32 >> shift_amt_int[4:0];
		endcase
	end
	// Trace: design.sv:4857:3
	genvar _gv_j_1;
	// Trace: design.sv:4858:3
	generate
		for (_gv_j_1 = 0; _gv_j_1 < 32; _gv_j_1 = _gv_j_1 + 1) begin : gen_shift_left_result
			localparam j = _gv_j_1;
			// Trace: design.sv:4860:7
			assign shift_left_result[j] = shift_right_result[31 - j];
		end
	endgenerate
	// Trace: design.sv:4864:3
	assign shift_result = (shift_left ? shift_left_result : shift_right_result);
	// Trace: design.sv:4876:3
	reg [3:0] is_equal;
	// Trace: design.sv:4877:3
	reg [3:0] is_greater;
	// Trace: design.sv:4880:3
	reg [3:0] cmp_signed;
	// Trace: design.sv:4881:3
	wire [3:0] is_equal_vec;
	// Trace: design.sv:4882:3
	wire [3:0] is_greater_vec;
	// Trace: design.sv:4883:3
	reg [31:0] operand_b_eq;
	// Trace: design.sv:4884:3
	wire is_equal_clip;
	// Trace: design.sv:4888:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:4889:5
		operand_b_eq = operand_b_neg;
		// Trace: design.sv:4890:5
		if (operator_i == sv2v_cast_C07C4(7'b0010111))
			// Trace: design.sv:4890:34
			operand_b_eq = 1'sb0;
		else
			// Trace: design.sv:4891:10
			operand_b_eq = operand_b_neg;
	end
	// Trace: design.sv:4893:3
	assign is_equal_clip = operand_a_i == operand_b_eq;
	// Trace: design.sv:4895:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:4896:5
		cmp_signed = 4'b0000;
		// Trace: design.sv:4898:5
		(* full_case, parallel_case *)
		case (operator_i)
			sv2v_cast_C07C4(7'b0001000), sv2v_cast_C07C4(7'b0001010), sv2v_cast_C07C4(7'b0000000), sv2v_cast_C07C4(7'b0000100), sv2v_cast_C07C4(7'b0000010), sv2v_cast_C07C4(7'b0000110), sv2v_cast_C07C4(7'b0010000), sv2v_cast_C07C4(7'b0010010), sv2v_cast_C07C4(7'b0010100), sv2v_cast_C07C4(7'b0010110), sv2v_cast_C07C4(7'b0010111):
				// Trace: design.sv:4910:9
				case (vector_mode_i)
					cv32e40p_pkg_VEC_MODE8:
						// Trace: design.sv:4911:23
						cmp_signed[3:0] = 4'b1111;
					cv32e40p_pkg_VEC_MODE16:
						// Trace: design.sv:4912:23
						cmp_signed[3:0] = 4'b1010;
					default:
						// Trace: design.sv:4913:23
						cmp_signed[3:0] = 4'b1000;
				endcase
			default:
				;
		endcase
	end
	// Trace: design.sv:4923:3
	genvar _gv_i_1;
	// Trace: design.sv:4924:3
	generate
		for (_gv_i_1 = 0; _gv_i_1 < 4; _gv_i_1 = _gv_i_1 + 1) begin : gen_is_vec
			localparam i = _gv_i_1;
			// Trace: design.sv:4926:7
			assign is_equal_vec[i] = operand_a_i[(8 * i) + 7:8 * i] == operand_b_i[(8 * i) + 7:i * 8];
			// Trace: design.sv:4927:7
			assign is_greater_vec[i] = $signed({operand_a_i[(8 * i) + 7] & cmp_signed[i], operand_a_i[(8 * i) + 7:8 * i]}) > $signed({operand_b_i[(8 * i) + 7] & cmp_signed[i], operand_b_i[(8 * i) + 7:i * 8]});
		end
	endgenerate
	// Trace: design.sv:4937:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:4939:5
		is_equal[3:0] = {4 {((is_equal_vec[3] & is_equal_vec[2]) & is_equal_vec[1]) & is_equal_vec[0]}};
		// Trace: design.sv:4940:5
		is_greater[3:0] = {4 {is_greater_vec[3] | (is_equal_vec[3] & (is_greater_vec[2] | (is_equal_vec[2] & (is_greater_vec[1] | (is_equal_vec[1] & is_greater_vec[0])))))}};
		// Trace: design.sv:4944:5
		case (vector_mode_i)
			cv32e40p_pkg_VEC_MODE16: begin
				// Trace: design.sv:4946:9
				is_equal[1:0] = {2 {is_equal_vec[0] & is_equal_vec[1]}};
				// Trace: design.sv:4947:9
				is_equal[3:2] = {2 {is_equal_vec[2] & is_equal_vec[3]}};
				// Trace: design.sv:4948:9
				is_greater[1:0] = {2 {is_greater_vec[1] | (is_equal_vec[1] & is_greater_vec[0])}};
				// Trace: design.sv:4949:9
				is_greater[3:2] = {2 {is_greater_vec[3] | (is_equal_vec[3] & is_greater_vec[2])}};
			end
			cv32e40p_pkg_VEC_MODE8: begin
				// Trace: design.sv:4953:9
				is_equal[3:0] = is_equal_vec[3:0];
				// Trace: design.sv:4954:9
				is_greater[3:0] = is_greater_vec[3:0];
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:4962:3
	reg [3:0] cmp_result;
	// Trace: design.sv:4964:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:4965:5
		cmp_result = is_equal;
		// Trace: design.sv:4966:5
		(* full_case, parallel_case *)
		case (operator_i)
			sv2v_cast_C07C4(7'b0001100):
				// Trace: design.sv:4967:47
				cmp_result = is_equal;
			sv2v_cast_C07C4(7'b0001101):
				// Trace: design.sv:4968:47
				cmp_result = ~is_equal;
			sv2v_cast_C07C4(7'b0001000), sv2v_cast_C07C4(7'b0001001):
				// Trace: design.sv:4969:47
				cmp_result = is_greater;
			sv2v_cast_C07C4(7'b0001010), sv2v_cast_C07C4(7'b0001011):
				// Trace: design.sv:4970:47
				cmp_result = is_greater | is_equal;
			sv2v_cast_C07C4(7'b0000000), sv2v_cast_C07C4(7'b0000010), sv2v_cast_C07C4(7'b0000001), sv2v_cast_C07C4(7'b0000011):
				// Trace: design.sv:4971:47
				cmp_result = ~(is_greater | is_equal);
			sv2v_cast_C07C4(7'b0000110), sv2v_cast_C07C4(7'b0000111), sv2v_cast_C07C4(7'b0000100), sv2v_cast_C07C4(7'b0000101):
				// Trace: design.sv:4972:47
				cmp_result = ~is_greater;
			default:
				;
		endcase
	end
	// Trace: design.sv:4977:3
	assign comparison_result_o = cmp_result[3];
	// Trace: design.sv:4981:3
	wire [31:0] result_minmax;
	// Trace: design.sv:4982:3
	wire [3:0] sel_minmax;
	// Trace: design.sv:4983:3
	wire do_min;
	// Trace: design.sv:4984:3
	wire [31:0] minmax_b;
	// Trace: design.sv:4986:3
	assign minmax_b = (operator_i == sv2v_cast_C07C4(7'b0010100) ? adder_result : operand_b_i);
	// Trace: design.sv:4988:3
	assign do_min = (((operator_i == sv2v_cast_C07C4(7'b0010000)) || (operator_i == sv2v_cast_C07C4(7'b0010001))) || (operator_i == sv2v_cast_C07C4(7'b0010110))) || (operator_i == sv2v_cast_C07C4(7'b0010111));
	// Trace: design.sv:4991:3
	assign sel_minmax[3:0] = is_greater ^ {4 {do_min}};
	// Trace: design.sv:4993:3
	assign result_minmax[31:24] = (sel_minmax[3] == 1'b1 ? operand_a_i[31:24] : minmax_b[31:24]);
	// Trace: design.sv:4994:3
	assign result_minmax[23:16] = (sel_minmax[2] == 1'b1 ? operand_a_i[23:16] : minmax_b[23:16]);
	// Trace: design.sv:4995:3
	assign result_minmax[15:8] = (sel_minmax[1] == 1'b1 ? operand_a_i[15:8] : minmax_b[15:8]);
	// Trace: design.sv:4996:3
	assign result_minmax[7:0] = (sel_minmax[0] == 1'b1 ? operand_a_i[7:0] : minmax_b[7:0]);
	// Trace: design.sv:5001:3
	reg [31:0] clip_result;
	// Trace: design.sv:5003:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:5004:5
		clip_result = result_minmax;
		// Trace: design.sv:5005:5
		if (operator_i == sv2v_cast_C07C4(7'b0010111)) begin
			begin
				// Trace: design.sv:5006:7
				if (operand_a_i[31] || is_equal_clip)
					// Trace: design.sv:5007:9
					clip_result = 1'sb0;
				else
					// Trace: design.sv:5009:9
					clip_result = result_minmax;
			end
		end
		else
			// Trace: design.sv:5013:7
			if (adder_result_expanded[36] || is_equal_clip)
				// Trace: design.sv:5014:9
				clip_result = operand_b_neg;
			else
				// Trace: design.sv:5016:9
				clip_result = result_minmax;
	end
	// Trace: design.sv:5031:3
	reg [7:0] shuffle_byte_sel;
	// Trace: design.sv:5032:3
	reg [3:0] shuffle_reg_sel;
	// Trace: design.sv:5033:3
	reg [1:0] shuffle_reg1_sel;
	// Trace: design.sv:5034:3
	reg [1:0] shuffle_reg0_sel;
	// Trace: design.sv:5035:3
	reg [3:0] shuffle_through;
	// Trace: design.sv:5037:3
	wire [31:0] shuffle_r1;
	wire [31:0] shuffle_r0;
	// Trace: design.sv:5038:3
	wire [31:0] shuffle_r1_in;
	wire [31:0] shuffle_r0_in;
	// Trace: design.sv:5039:3
	wire [31:0] shuffle_result;
	// Trace: design.sv:5040:3
	wire [31:0] pack_result;
	// Trace: design.sv:5043:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:5044:5
		shuffle_reg_sel = 1'sb0;
		// Trace: design.sv:5045:5
		shuffle_reg1_sel = 2'b01;
		// Trace: design.sv:5046:5
		shuffle_reg0_sel = 2'b10;
		// Trace: design.sv:5047:5
		shuffle_through = 1'sb1;
		// Trace: design.sv:5049:5
		(* full_case, parallel_case *)
		case (operator_i)
			sv2v_cast_C07C4(7'b0111111), sv2v_cast_C07C4(7'b0111110): begin
				// Trace: design.sv:5051:9
				if (operator_i == sv2v_cast_C07C4(7'b0111110))
					// Trace: design.sv:5051:37
					shuffle_reg1_sel = 2'b11;
				if (vector_mode_i == cv32e40p_pkg_VEC_MODE8) begin
					// Trace: design.sv:5054:11
					shuffle_reg_sel[3:1] = 3'b111;
					// Trace: design.sv:5055:11
					shuffle_reg_sel[0] = 1'b0;
				end
				else begin
					// Trace: design.sv:5057:11
					shuffle_reg_sel[3:2] = 2'b11;
					// Trace: design.sv:5058:11
					shuffle_reg_sel[1:0] = 2'b00;
				end
			end
			sv2v_cast_C07C4(7'b0111000): begin
				// Trace: design.sv:5063:9
				shuffle_reg1_sel = 2'b00;
				// Trace: design.sv:5065:9
				if (vector_mode_i == cv32e40p_pkg_VEC_MODE8) begin
					// Trace: design.sv:5066:11
					shuffle_through = 4'b0011;
					// Trace: design.sv:5067:11
					shuffle_reg_sel = 4'b0001;
				end
				else
					// Trace: design.sv:5069:11
					shuffle_reg_sel = 4'b0011;
			end
			sv2v_cast_C07C4(7'b0111001): begin
				// Trace: design.sv:5074:9
				shuffle_reg1_sel = 2'b00;
				// Trace: design.sv:5076:9
				if (vector_mode_i == cv32e40p_pkg_VEC_MODE8) begin
					// Trace: design.sv:5077:11
					shuffle_through = 4'b1100;
					// Trace: design.sv:5078:11
					shuffle_reg_sel = 4'b0100;
				end
				else
					// Trace: design.sv:5080:11
					shuffle_reg_sel = 4'b0011;
			end
			sv2v_cast_C07C4(7'b0111011):
				// Trace: design.sv:5085:9
				(* full_case, parallel_case *)
				case (vector_mode_i)
					cv32e40p_pkg_VEC_MODE8: begin
						// Trace: design.sv:5087:13
						shuffle_reg_sel[3] = ~operand_b_i[26];
						// Trace: design.sv:5088:13
						shuffle_reg_sel[2] = ~operand_b_i[18];
						// Trace: design.sv:5089:13
						shuffle_reg_sel[1] = ~operand_b_i[10];
						// Trace: design.sv:5090:13
						shuffle_reg_sel[0] = ~operand_b_i[2];
					end
					cv32e40p_pkg_VEC_MODE16: begin
						// Trace: design.sv:5094:13
						shuffle_reg_sel[3] = ~operand_b_i[17];
						// Trace: design.sv:5095:13
						shuffle_reg_sel[2] = ~operand_b_i[17];
						// Trace: design.sv:5096:13
						shuffle_reg_sel[1] = ~operand_b_i[1];
						// Trace: design.sv:5097:13
						shuffle_reg_sel[0] = ~operand_b_i[1];
					end
					default:
						;
				endcase
			sv2v_cast_C07C4(7'b0101101):
				// Trace: design.sv:5104:9
				(* full_case, parallel_case *)
				case (vector_mode_i)
					cv32e40p_pkg_VEC_MODE8: begin
						// Trace: design.sv:5106:13
						shuffle_reg0_sel = 2'b00;
						// Trace: design.sv:5107:13
						(* full_case, parallel_case *)
						case (imm_vec_ext_i)
							2'b00:
								// Trace: design.sv:5109:17
								shuffle_reg_sel[3:0] = 4'b1110;
							2'b01:
								// Trace: design.sv:5112:17
								shuffle_reg_sel[3:0] = 4'b1101;
							2'b10:
								// Trace: design.sv:5115:17
								shuffle_reg_sel[3:0] = 4'b1011;
							2'b11:
								// Trace: design.sv:5118:17
								shuffle_reg_sel[3:0] = 4'b0111;
						endcase
					end
					cv32e40p_pkg_VEC_MODE16: begin
						// Trace: design.sv:5123:13
						shuffle_reg0_sel = 2'b01;
						// Trace: design.sv:5124:13
						shuffle_reg_sel[3] = ~imm_vec_ext_i[0];
						// Trace: design.sv:5125:13
						shuffle_reg_sel[2] = ~imm_vec_ext_i[0];
						// Trace: design.sv:5126:13
						shuffle_reg_sel[1] = imm_vec_ext_i[0];
						// Trace: design.sv:5127:13
						shuffle_reg_sel[0] = imm_vec_ext_i[0];
					end
					default:
						;
				endcase
			default:
				;
		endcase
	end
	// Trace: design.sv:5137:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:5138:5
		shuffle_byte_sel = 1'sb0;
		// Trace: design.sv:5141:5
		(* full_case, parallel_case *)
		case (operator_i)
			sv2v_cast_C07C4(7'b0111110), sv2v_cast_C07C4(7'b0111111):
				// Trace: design.sv:5143:9
				(* full_case, parallel_case *)
				case (vector_mode_i)
					cv32e40p_pkg_VEC_MODE8: begin
						// Trace: design.sv:5145:13
						shuffle_byte_sel[6+:2] = imm_vec_ext_i[1:0];
						// Trace: design.sv:5146:13
						shuffle_byte_sel[4+:2] = imm_vec_ext_i[1:0];
						// Trace: design.sv:5147:13
						shuffle_byte_sel[2+:2] = imm_vec_ext_i[1:0];
						// Trace: design.sv:5148:13
						shuffle_byte_sel[0+:2] = imm_vec_ext_i[1:0];
					end
					cv32e40p_pkg_VEC_MODE16: begin
						// Trace: design.sv:5152:13
						shuffle_byte_sel[6+:2] = {imm_vec_ext_i[0], 1'b1};
						// Trace: design.sv:5153:13
						shuffle_byte_sel[4+:2] = {imm_vec_ext_i[0], 1'b1};
						// Trace: design.sv:5154:13
						shuffle_byte_sel[2+:2] = {imm_vec_ext_i[0], 1'b1};
						// Trace: design.sv:5155:13
						shuffle_byte_sel[0+:2] = {imm_vec_ext_i[0], 1'b0};
					end
					default:
						;
				endcase
			sv2v_cast_C07C4(7'b0111000):
				// Trace: design.sv:5163:9
				(* full_case, parallel_case *)
				case (vector_mode_i)
					cv32e40p_pkg_VEC_MODE8: begin
						// Trace: design.sv:5165:13
						shuffle_byte_sel[6+:2] = 2'b00;
						// Trace: design.sv:5166:13
						shuffle_byte_sel[4+:2] = 2'b00;
						// Trace: design.sv:5167:13
						shuffle_byte_sel[2+:2] = 2'b00;
						// Trace: design.sv:5168:13
						shuffle_byte_sel[0+:2] = 2'b00;
					end
					cv32e40p_pkg_VEC_MODE16: begin
						// Trace: design.sv:5172:13
						shuffle_byte_sel[6+:2] = 2'b01;
						// Trace: design.sv:5173:13
						shuffle_byte_sel[4+:2] = 2'b00;
						// Trace: design.sv:5174:13
						shuffle_byte_sel[2+:2] = 2'b01;
						// Trace: design.sv:5175:13
						shuffle_byte_sel[0+:2] = 2'b00;
					end
					default:
						;
				endcase
			sv2v_cast_C07C4(7'b0111001):
				// Trace: design.sv:5183:9
				(* full_case, parallel_case *)
				case (vector_mode_i)
					cv32e40p_pkg_VEC_MODE8: begin
						// Trace: design.sv:5185:13
						shuffle_byte_sel[6+:2] = 2'b00;
						// Trace: design.sv:5186:13
						shuffle_byte_sel[4+:2] = 2'b00;
						// Trace: design.sv:5187:13
						shuffle_byte_sel[2+:2] = 2'b00;
						// Trace: design.sv:5188:13
						shuffle_byte_sel[0+:2] = 2'b00;
					end
					cv32e40p_pkg_VEC_MODE16: begin
						// Trace: design.sv:5192:13
						shuffle_byte_sel[6+:2] = 2'b11;
						// Trace: design.sv:5193:13
						shuffle_byte_sel[4+:2] = 2'b10;
						// Trace: design.sv:5194:13
						shuffle_byte_sel[2+:2] = 2'b11;
						// Trace: design.sv:5195:13
						shuffle_byte_sel[0+:2] = 2'b10;
					end
					default:
						;
				endcase
			sv2v_cast_C07C4(7'b0111011), sv2v_cast_C07C4(7'b0111010):
				// Trace: design.sv:5203:9
				(* full_case, parallel_case *)
				case (vector_mode_i)
					cv32e40p_pkg_VEC_MODE8: begin
						// Trace: design.sv:5205:13
						shuffle_byte_sel[6+:2] = operand_b_i[25:24];
						// Trace: design.sv:5206:13
						shuffle_byte_sel[4+:2] = operand_b_i[17:16];
						// Trace: design.sv:5207:13
						shuffle_byte_sel[2+:2] = operand_b_i[9:8];
						// Trace: design.sv:5208:13
						shuffle_byte_sel[0+:2] = operand_b_i[1:0];
					end
					cv32e40p_pkg_VEC_MODE16: begin
						// Trace: design.sv:5212:13
						shuffle_byte_sel[6+:2] = {operand_b_i[16], 1'b1};
						// Trace: design.sv:5213:13
						shuffle_byte_sel[4+:2] = {operand_b_i[16], 1'b0};
						// Trace: design.sv:5214:13
						shuffle_byte_sel[2+:2] = {operand_b_i[0], 1'b1};
						// Trace: design.sv:5215:13
						shuffle_byte_sel[0+:2] = {operand_b_i[0], 1'b0};
					end
					default:
						;
				endcase
			sv2v_cast_C07C4(7'b0101101): begin
				// Trace: design.sv:5222:9
				shuffle_byte_sel[6+:2] = 2'b11;
				// Trace: design.sv:5223:9
				shuffle_byte_sel[4+:2] = 2'b10;
				// Trace: design.sv:5224:9
				shuffle_byte_sel[2+:2] = 2'b01;
				// Trace: design.sv:5225:9
				shuffle_byte_sel[0+:2] = 2'b00;
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:5232:3
	assign shuffle_r0_in = (shuffle_reg0_sel[1] ? operand_a_i : (shuffle_reg0_sel[0] ? {2 {operand_a_i[15:0]}} : {4 {operand_a_i[7:0]}}));
	// Trace: design.sv:5236:3
	assign shuffle_r1_in = (shuffle_reg1_sel[1] ? {{8 {operand_a_i[31]}}, {8 {operand_a_i[23]}}, {8 {operand_a_i[15]}}, {8 {operand_a_i[7]}}} : (shuffle_reg1_sel[0] ? operand_c_i : operand_b_i));
	// Trace: design.sv:5240:3
	assign shuffle_r0[31:24] = (shuffle_byte_sel[7] ? (shuffle_byte_sel[6] ? shuffle_r0_in[31:24] : shuffle_r0_in[23:16]) : (shuffle_byte_sel[6] ? shuffle_r0_in[15:8] : shuffle_r0_in[7:0]));
	// Trace: design.sv:5243:3
	assign shuffle_r0[23:16] = (shuffle_byte_sel[5] ? (shuffle_byte_sel[4] ? shuffle_r0_in[31:24] : shuffle_r0_in[23:16]) : (shuffle_byte_sel[4] ? shuffle_r0_in[15:8] : shuffle_r0_in[7:0]));
	// Trace: design.sv:5246:3
	assign shuffle_r0[15:8] = (shuffle_byte_sel[3] ? (shuffle_byte_sel[2] ? shuffle_r0_in[31:24] : shuffle_r0_in[23:16]) : (shuffle_byte_sel[2] ? shuffle_r0_in[15:8] : shuffle_r0_in[7:0]));
	// Trace: design.sv:5249:3
	assign shuffle_r0[7:0] = (shuffle_byte_sel[1] ? (shuffle_byte_sel[0] ? shuffle_r0_in[31:24] : shuffle_r0_in[23:16]) : (shuffle_byte_sel[0] ? shuffle_r0_in[15:8] : shuffle_r0_in[7:0]));
	// Trace: design.sv:5253:3
	assign shuffle_r1[31:24] = (shuffle_byte_sel[7] ? (shuffle_byte_sel[6] ? shuffle_r1_in[31:24] : shuffle_r1_in[23:16]) : (shuffle_byte_sel[6] ? shuffle_r1_in[15:8] : shuffle_r1_in[7:0]));
	// Trace: design.sv:5256:3
	assign shuffle_r1[23:16] = (shuffle_byte_sel[5] ? (shuffle_byte_sel[4] ? shuffle_r1_in[31:24] : shuffle_r1_in[23:16]) : (shuffle_byte_sel[4] ? shuffle_r1_in[15:8] : shuffle_r1_in[7:0]));
	// Trace: design.sv:5259:3
	assign shuffle_r1[15:8] = (shuffle_byte_sel[3] ? (shuffle_byte_sel[2] ? shuffle_r1_in[31:24] : shuffle_r1_in[23:16]) : (shuffle_byte_sel[2] ? shuffle_r1_in[15:8] : shuffle_r1_in[7:0]));
	// Trace: design.sv:5262:3
	assign shuffle_r1[7:0] = (shuffle_byte_sel[1] ? (shuffle_byte_sel[0] ? shuffle_r1_in[31:24] : shuffle_r1_in[23:16]) : (shuffle_byte_sel[0] ? shuffle_r1_in[15:8] : shuffle_r1_in[7:0]));
	// Trace: design.sv:5266:3
	assign shuffle_result[31:24] = (shuffle_reg_sel[3] ? shuffle_r1[31:24] : shuffle_r0[31:24]);
	// Trace: design.sv:5267:3
	assign shuffle_result[23:16] = (shuffle_reg_sel[2] ? shuffle_r1[23:16] : shuffle_r0[23:16]);
	// Trace: design.sv:5268:3
	assign shuffle_result[15:8] = (shuffle_reg_sel[1] ? shuffle_r1[15:8] : shuffle_r0[15:8]);
	// Trace: design.sv:5269:3
	assign shuffle_result[7:0] = (shuffle_reg_sel[0] ? shuffle_r1[7:0] : shuffle_r0[7:0]);
	// Trace: design.sv:5271:3
	assign pack_result[31:24] = (shuffle_through[3] ? shuffle_result[31:24] : operand_c_i[31:24]);
	// Trace: design.sv:5272:3
	assign pack_result[23:16] = (shuffle_through[2] ? shuffle_result[23:16] : operand_c_i[23:16]);
	// Trace: design.sv:5273:3
	assign pack_result[15:8] = (shuffle_through[1] ? shuffle_result[15:8] : operand_c_i[15:8]);
	// Trace: design.sv:5274:3
	assign pack_result[7:0] = (shuffle_through[0] ? shuffle_result[7:0] : operand_c_i[7:0]);
	// Trace: design.sv:5286:3
	reg [31:0] ff_input;
	// Trace: design.sv:5287:3
	wire [5:0] cnt_result;
	// Trace: design.sv:5288:3
	wire [5:0] clb_result;
	// Trace: design.sv:5289:3
	wire [4:0] ff1_result;
	// Trace: design.sv:5290:3
	wire ff_no_one;
	// Trace: design.sv:5291:3
	wire [4:0] fl1_result;
	// Trace: design.sv:5292:3
	reg [5:0] bitop_result;
	// Trace: design.sv:5294:3
	cv32e40p_popcnt popcnt_i(
		.in_i(operand_a_i),
		.result_o(cnt_result)
	);
	// Trace: design.sv:5299:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:5300:5
		ff_input = 1'sb0;
		// Trace: design.sv:5302:5
		case (operator_i)
			sv2v_cast_C07C4(7'b0110110):
				// Trace: design.sv:5303:16
				ff_input = operand_a_i;
			sv2v_cast_C07C4(7'b0110000), sv2v_cast_C07C4(7'b0110010), sv2v_cast_C07C4(7'b0110111):
				// Trace: design.sv:5305:36
				ff_input = operand_a_rev;
			sv2v_cast_C07C4(7'b0110001), sv2v_cast_C07C4(7'b0110011), sv2v_cast_C07C4(7'b0110101):
				// Trace: design.sv:5308:9
				if (operand_a_i[31])
					// Trace: design.sv:5308:30
					ff_input = operand_a_neg_rev;
				else
					// Trace: design.sv:5309:14
					ff_input = operand_a_rev;
		endcase
	end
	// Trace: design.sv:5314:3
	cv32e40p_ff_one ff_one_i(
		.in_i(ff_input),
		.first_one_o(ff1_result),
		.no_ones_o(ff_no_one)
	);
	// Trace: design.sv:5322:3
	assign fl1_result = 5'd31 - ff1_result;
	// Trace: design.sv:5323:3
	assign clb_result = ff1_result - 5'd1;
	// Trace: design.sv:5325:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:5326:5
		bitop_result = 1'sb0;
		// Trace: design.sv:5327:5
		case (operator_i)
			sv2v_cast_C07C4(7'b0110110):
				// Trace: design.sv:5328:16
				bitop_result = (ff_no_one ? 6'd32 : {1'b0, ff1_result});
			sv2v_cast_C07C4(7'b0110111):
				// Trace: design.sv:5329:16
				bitop_result = (ff_no_one ? 6'd32 : {1'b0, fl1_result});
			sv2v_cast_C07C4(7'b0110100):
				// Trace: design.sv:5330:16
				bitop_result = cnt_result;
			sv2v_cast_C07C4(7'b0110101):
				// Trace: design.sv:5332:9
				if (ff_no_one) begin
					begin
						// Trace: design.sv:5333:11
						if (operand_a_i[31])
							// Trace: design.sv:5333:32
							bitop_result = 6'd31;
						else
							// Trace: design.sv:5334:16
							bitop_result = 1'sb0;
					end
				end
				else
					// Trace: design.sv:5336:11
					bitop_result = clb_result;
			default:
				;
		endcase
	end
	// Trace: design.sv:5353:3
	wire extract_is_signed;
	// Trace: design.sv:5354:3
	wire extract_sign;
	// Trace: design.sv:5355:3
	wire [31:0] bmask_first;
	wire [31:0] bmask_inv;
	// Trace: design.sv:5356:3
	wire [31:0] bextins_and;
	// Trace: design.sv:5357:3
	wire [31:0] bextins_result;
	wire [31:0] bclr_result;
	wire [31:0] bset_result;
	// Trace: design.sv:5362:3
	assign bmask_first = 32'hfffffffe << bmask_a_i;
	// Trace: design.sv:5363:3
	assign bmask = ~bmask_first << bmask_b_i;
	// Trace: design.sv:5364:3
	assign bmask_inv = ~bmask;
	// Trace: design.sv:5366:3
	assign bextins_and = (operator_i == sv2v_cast_C07C4(7'b0101010) ? operand_c_i : {32 {extract_sign}});
	// Trace: design.sv:5368:3
	assign extract_is_signed = operator_i == sv2v_cast_C07C4(7'b0101000);
	// Trace: design.sv:5369:3
	assign extract_sign = extract_is_signed & shift_result[bmask_a_i];
	// Trace: design.sv:5371:3
	assign bextins_result = (bmask & shift_result) | (bextins_and & bmask_inv);
	// Trace: design.sv:5373:3
	assign bclr_result = operand_a_i & bmask_inv;
	// Trace: design.sv:5374:3
	assign bset_result = operand_a_i | bmask;
	// Trace: design.sv:5386:3
	wire [31:0] radix_2_rev;
	// Trace: design.sv:5387:3
	wire [31:0] radix_4_rev;
	// Trace: design.sv:5388:3
	wire [31:0] radix_8_rev;
	// Trace: design.sv:5389:3
	reg [31:0] reverse_result;
	// Trace: design.sv:5390:3
	wire [1:0] radix_mux_sel;
	// Trace: design.sv:5392:3
	assign radix_mux_sel = bmask_a_i[1:0];
	// Trace: design.sv:5394:3
	generate
		for (_gv_j_1 = 0; _gv_j_1 < 32; _gv_j_1 = _gv_j_1 + 1) begin : gen_radix_2_rev
			localparam j = _gv_j_1;
			// Trace: design.sv:5397:7
			assign radix_2_rev[j] = shift_result[31 - j];
		end
		for (_gv_j_1 = 0; _gv_j_1 < 16; _gv_j_1 = _gv_j_1 + 1) begin : gen_radix_4_rev
			localparam j = _gv_j_1;
			// Trace: design.sv:5401:7
			assign radix_4_rev[(2 * j) + 1:2 * j] = shift_result[31 - (j * 2):(31 - (j * 2)) - 1];
		end
		for (_gv_j_1 = 0; _gv_j_1 < 10; _gv_j_1 = _gv_j_1 + 1) begin : gen_radix_8_rev
			localparam j = _gv_j_1;
			// Trace: design.sv:5405:7
			assign radix_8_rev[(3 * j) + 2:3 * j] = shift_result[31 - (j * 3):(31 - (j * 3)) - 2];
		end
	endgenerate
	// Trace: design.sv:5407:5
	assign radix_8_rev[31:30] = 2'b00;
	// Trace: design.sv:5410:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:5411:5
		reverse_result = 1'sb0;
		// Trace: design.sv:5413:5
		(* full_case, parallel_case *)
		case (radix_mux_sel)
			2'b00:
				// Trace: design.sv:5414:14
				reverse_result = radix_2_rev;
			2'b01:
				// Trace: design.sv:5415:14
				reverse_result = radix_4_rev;
			2'b10:
				// Trace: design.sv:5416:14
				reverse_result = radix_8_rev;
			default:
				// Trace: design.sv:5418:16
				reverse_result = radix_2_rev;
		endcase
	end
	// Trace: design.sv:5431:3
	wire [31:0] result_div;
	// Trace: design.sv:5432:3
	wire div_ready;
	// Trace: design.sv:5433:3
	wire div_signed;
	// Trace: design.sv:5434:3
	wire div_op_a_signed;
	// Trace: design.sv:5435:3
	wire [5:0] div_shift_int;
	// Trace: design.sv:5437:3
	assign div_signed = operator_i[0];
	// Trace: design.sv:5439:3
	assign div_op_a_signed = operand_a_i[31] & div_signed;
	// Trace: design.sv:5441:3
	assign div_shift_int = (ff_no_one ? 6'd31 : clb_result);
	// Trace: design.sv:5442:3
	assign div_shift = div_shift_int + (div_op_a_signed ? 6'd0 : 6'd1);
	// Trace: design.sv:5444:3
	assign div_valid = enable_i & ((((operator_i == sv2v_cast_C07C4(7'b0110001)) || (operator_i == sv2v_cast_C07C4(7'b0110000))) || (operator_i == sv2v_cast_C07C4(7'b0110011))) || (operator_i == sv2v_cast_C07C4(7'b0110010)));
	// Trace: design.sv:5448:3
	cv32e40p_alu_div alu_div_i(
		.Clk_CI(clk),
		.Rst_RBI(rst_n),
		.OpA_DI(operand_b_i),
		.OpB_DI(shift_left_result),
		.OpBShift_DI(div_shift),
		.OpBIsZero_SI(cnt_result == 0),
		.OpBSign_SI(div_op_a_signed),
		.OpCode_SI(operator_i[1:0]),
		.Res_DO(result_div),
		.InVld_SI(div_valid),
		.OutRdy_SI(ex_ready_i),
		.OutVld_SO(div_ready)
	);
	// Trace: design.sv:5478:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:5479:5
		result_o = 1'sb0;
		// Trace: design.sv:5481:5
		(* full_case, parallel_case *)
		case (operator_i)
			sv2v_cast_C07C4(7'b0010101):
				// Trace: design.sv:5483:16
				result_o = operand_a_i & operand_b_i;
			sv2v_cast_C07C4(7'b0101110):
				// Trace: design.sv:5484:16
				result_o = operand_a_i | operand_b_i;
			sv2v_cast_C07C4(7'b0101111):
				// Trace: design.sv:5485:16
				result_o = operand_a_i ^ operand_b_i;
			sv2v_cast_C07C4(7'b0011000), sv2v_cast_C07C4(7'b0011100), sv2v_cast_C07C4(7'b0011010), sv2v_cast_C07C4(7'b0011110), sv2v_cast_C07C4(7'b0011001), sv2v_cast_C07C4(7'b0011101), sv2v_cast_C07C4(7'b0011011), sv2v_cast_C07C4(7'b0011111), sv2v_cast_C07C4(7'b0100111), sv2v_cast_C07C4(7'b0100101), sv2v_cast_C07C4(7'b0100100), sv2v_cast_C07C4(7'b0100110):
				// Trace: design.sv:5493:7
				result_o = shift_result;
			sv2v_cast_C07C4(7'b0101010), sv2v_cast_C07C4(7'b0101000), sv2v_cast_C07C4(7'b0101001):
				// Trace: design.sv:5496:38
				result_o = bextins_result;
			sv2v_cast_C07C4(7'b0101011):
				// Trace: design.sv:5498:17
				result_o = bclr_result;
			sv2v_cast_C07C4(7'b0101100):
				// Trace: design.sv:5499:17
				result_o = bset_result;
			sv2v_cast_C07C4(7'b1001001):
				// Trace: design.sv:5502:17
				result_o = reverse_result;
			sv2v_cast_C07C4(7'b0111010), sv2v_cast_C07C4(7'b0111011), sv2v_cast_C07C4(7'b0111000), sv2v_cast_C07C4(7'b0111001), sv2v_cast_C07C4(7'b0111111), sv2v_cast_C07C4(7'b0111110), sv2v_cast_C07C4(7'b0101101):
				// Trace: design.sv:5505:78
				result_o = pack_result;
			sv2v_cast_C07C4(7'b0010000), sv2v_cast_C07C4(7'b0010001), sv2v_cast_C07C4(7'b0010010), sv2v_cast_C07C4(7'b0010011):
				// Trace: design.sv:5508:45
				result_o = result_minmax;
			sv2v_cast_C07C4(7'b0010100):
				// Trace: design.sv:5511:16
				result_o = (is_clpx_i ? {adder_result[31:16], operand_a_i[15:0]} : result_minmax);
			sv2v_cast_C07C4(7'b0010110), sv2v_cast_C07C4(7'b0010111):
				// Trace: design.sv:5513:28
				result_o = clip_result;
			sv2v_cast_C07C4(7'b0001100), sv2v_cast_C07C4(7'b0001101), sv2v_cast_C07C4(7'b0001001), sv2v_cast_C07C4(7'b0001011), sv2v_cast_C07C4(7'b0000001), sv2v_cast_C07C4(7'b0000101), sv2v_cast_C07C4(7'b0001000), sv2v_cast_C07C4(7'b0001010), sv2v_cast_C07C4(7'b0000000), sv2v_cast_C07C4(7'b0000100): begin
				// Trace: design.sv:5517:9
				result_o[31:24] = {8 {cmp_result[3]}};
				// Trace: design.sv:5518:9
				result_o[23:16] = {8 {cmp_result[2]}};
				// Trace: design.sv:5519:9
				result_o[15:8] = {8 {cmp_result[1]}};
				// Trace: design.sv:5520:9
				result_o[7:0] = {8 {cmp_result[0]}};
			end
			sv2v_cast_C07C4(7'b0000010), sv2v_cast_C07C4(7'b0000011), sv2v_cast_C07C4(7'b0000110), sv2v_cast_C07C4(7'b0000111):
				// Trace: design.sv:5523:49
				result_o = {31'b0000000000000000000000000000000, comparison_result_o};
			sv2v_cast_C07C4(7'b0110110), sv2v_cast_C07C4(7'b0110111), sv2v_cast_C07C4(7'b0110101), sv2v_cast_C07C4(7'b0110100):
				// Trace: design.sv:5525:43
				result_o = {26'h0000000, bitop_result[5:0]};
			sv2v_cast_C07C4(7'b0110001), sv2v_cast_C07C4(7'b0110000), sv2v_cast_C07C4(7'b0110011), sv2v_cast_C07C4(7'b0110010):
				// Trace: design.sv:5528:45
				result_o = result_div;
			default:
				;
		endcase
	end
	// Trace: design.sv:5534:3
	assign ready_o = div_ready;
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_alu_div (
	Clk_CI,
	Rst_RBI,
	OpA_DI,
	OpB_DI,
	OpBShift_DI,
	OpBIsZero_SI,
	OpBSign_SI,
	OpCode_SI,
	InVld_SI,
	OutRdy_SI,
	OutVld_SO,
	Res_DO
);
	reg _sv2v_0;
	// Trace: design.sv:5563:15
	parameter C_WIDTH = 32;
	// Trace: design.sv:5564:15
	parameter C_LOG_WIDTH = 6;
	// Trace: design.sv:5566:5
	input wire Clk_CI;
	// Trace: design.sv:5567:5
	input wire Rst_RBI;
	// Trace: design.sv:5569:5
	input wire [C_WIDTH - 1:0] OpA_DI;
	// Trace: design.sv:5570:5
	input wire [C_WIDTH - 1:0] OpB_DI;
	// Trace: design.sv:5571:5
	input wire [C_LOG_WIDTH - 1:0] OpBShift_DI;
	// Trace: design.sv:5572:5
	input wire OpBIsZero_SI;
	// Trace: design.sv:5574:5
	input wire OpBSign_SI;
	// Trace: design.sv:5575:5
	input wire [1:0] OpCode_SI;
	// Trace: design.sv:5577:5
	input wire InVld_SI;
	// Trace: design.sv:5579:5
	input wire OutRdy_SI;
	// Trace: design.sv:5580:5
	output reg OutVld_SO;
	// Trace: design.sv:5581:5
	output wire [C_WIDTH - 1:0] Res_DO;
	// Trace: design.sv:5588:3
	reg [C_WIDTH - 1:0] ResReg_DP;
	wire [C_WIDTH - 1:0] ResReg_DN;
	// Trace: design.sv:5589:3
	wire [C_WIDTH - 1:0] ResReg_DP_rev;
	// Trace: design.sv:5590:3
	reg [C_WIDTH - 1:0] AReg_DP;
	wire [C_WIDTH - 1:0] AReg_DN;
	// Trace: design.sv:5591:3
	reg [C_WIDTH - 1:0] BReg_DP;
	wire [C_WIDTH - 1:0] BReg_DN;
	// Trace: design.sv:5593:3
	wire RemSel_SN;
	reg RemSel_SP;
	// Trace: design.sv:5594:3
	wire CompInv_SN;
	reg CompInv_SP;
	// Trace: design.sv:5595:3
	wire ResInv_SN;
	reg ResInv_SP;
	// Trace: design.sv:5597:3
	wire [C_WIDTH - 1:0] AddMux_D;
	// Trace: design.sv:5598:3
	wire [C_WIDTH - 1:0] AddOut_D;
	// Trace: design.sv:5599:3
	wire [C_WIDTH - 1:0] AddTmp_D;
	// Trace: design.sv:5600:3
	wire [C_WIDTH - 1:0] BMux_D;
	// Trace: design.sv:5601:3
	wire [C_WIDTH - 1:0] OutMux_D;
	// Trace: design.sv:5603:3
	reg [C_LOG_WIDTH - 1:0] Cnt_DP;
	wire [C_LOG_WIDTH - 1:0] Cnt_DN;
	// Trace: design.sv:5604:3
	wire CntZero_S;
	// Trace: design.sv:5606:3
	reg ARegEn_S;
	reg BRegEn_S;
	reg ResRegEn_S;
	wire ABComp_S;
	wire PmSel_S;
	reg LoadEn_S;
	// Trace: design.sv:5608:3
	reg [1:0] State_SN;
	reg [1:0] State_SP;
	// Trace: design.sv:5620:3
	assign PmSel_S = LoadEn_S & ~(OpCode_SI[0] & (OpA_DI[C_WIDTH - 1] ^ OpBSign_SI));
	// Trace: design.sv:5623:3
	assign AddMux_D = (LoadEn_S ? OpA_DI : BReg_DP);
	// Trace: design.sv:5626:3
	assign BMux_D = (LoadEn_S ? OpB_DI : {CompInv_SP, BReg_DP[C_WIDTH - 1:1]});
	// Trace: design.sv:5628:3
	genvar _gv_index_1;
	// Trace: design.sv:5629:3
	generate
		for (_gv_index_1 = 0; _gv_index_1 < C_WIDTH; _gv_index_1 = _gv_index_1 + 1) begin : gen_bit_swapping
			localparam index = _gv_index_1;
			// Trace: design.sv:5631:7
			assign ResReg_DP_rev[index] = ResReg_DP[(C_WIDTH - 1) - index];
		end
	endgenerate
	// Trace: design.sv:5635:3
	assign OutMux_D = (RemSel_SP ? AReg_DP : ResReg_DP_rev);
	// Trace: design.sv:5638:3
	assign Res_DO = (ResInv_SP ? -$signed(OutMux_D) : OutMux_D);
	// Trace: design.sv:5641:3
	assign ABComp_S = ((AReg_DP == BReg_DP) | ((AReg_DP > BReg_DP) ^ CompInv_SP)) & (|AReg_DP | OpBIsZero_SI);
	// Trace: design.sv:5644:3
	assign AddTmp_D = (LoadEn_S ? 0 : AReg_DP);
	// Trace: design.sv:5645:3
	assign AddOut_D = (PmSel_S ? AddTmp_D + AddMux_D : AddTmp_D - $signed(AddMux_D));
	// Trace: design.sv:5651:3
	assign Cnt_DN = (LoadEn_S ? OpBShift_DI : (~CntZero_S ? Cnt_DP - 1 : Cnt_DP));
	// Trace: design.sv:5653:3
	assign CntZero_S = ~(|Cnt_DP);
	// Trace: design.sv:5659:3
	always @(*) begin : p_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:5661:5
		State_SN = State_SP;
		// Trace: design.sv:5663:5
		OutVld_SO = 1'b0;
		// Trace: design.sv:5665:5
		LoadEn_S = 1'b0;
		// Trace: design.sv:5667:5
		ARegEn_S = 1'b0;
		// Trace: design.sv:5668:5
		BRegEn_S = 1'b0;
		// Trace: design.sv:5669:5
		ResRegEn_S = 1'b0;
		// Trace: design.sv:5671:5
		case (State_SP)
			2'd0: begin
				// Trace: design.sv:5674:9
				OutVld_SO = 1'b1;
				// Trace: design.sv:5676:9
				if (InVld_SI) begin
					// Trace: design.sv:5677:11
					OutVld_SO = 1'b0;
					// Trace: design.sv:5678:11
					ARegEn_S = 1'b1;
					// Trace: design.sv:5679:11
					BRegEn_S = 1'b1;
					// Trace: design.sv:5680:11
					LoadEn_S = 1'b1;
					// Trace: design.sv:5681:11
					State_SN = 2'd1;
				end
			end
			2'd1: begin
				// Trace: design.sv:5687:9
				ARegEn_S = ABComp_S;
				// Trace: design.sv:5688:9
				BRegEn_S = 1'b1;
				// Trace: design.sv:5689:9
				ResRegEn_S = 1'b1;
				// Trace: design.sv:5693:9
				if (CntZero_S)
					// Trace: design.sv:5694:11
					State_SN = 2'd2;
			end
			2'd2: begin
				// Trace: design.sv:5699:9
				OutVld_SO = 1'b1;
				// Trace: design.sv:5701:9
				if (OutRdy_SI)
					// Trace: design.sv:5702:11
					State_SN = 2'd0;
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:5717:3
	assign RemSel_SN = (LoadEn_S ? OpCode_SI[1] : RemSel_SP);
	// Trace: design.sv:5718:3
	assign CompInv_SN = (LoadEn_S ? OpBSign_SI : CompInv_SP);
	// Trace: design.sv:5719:3
	assign ResInv_SN = (LoadEn_S ? ((~OpBIsZero_SI | OpCode_SI[1]) & OpCode_SI[0]) & (OpA_DI[C_WIDTH - 1] ^ OpBSign_SI) : ResInv_SP);
	// Trace: design.sv:5723:3
	assign AReg_DN = (ARegEn_S ? AddOut_D : AReg_DP);
	// Trace: design.sv:5724:3
	assign BReg_DN = (BRegEn_S ? BMux_D : BReg_DP);
	// Trace: design.sv:5725:3
	assign ResReg_DN = (LoadEn_S ? {C_WIDTH {1'sb0}} : (ResRegEn_S ? {ABComp_S, ResReg_DP[C_WIDTH - 1:1]} : ResReg_DP));
	// Trace: design.sv:5729:3
	always @(posedge Clk_CI or negedge Rst_RBI) begin : p_regs
		// Trace: design.sv:5730:5
		if (~Rst_RBI) begin
			// Trace: design.sv:5731:7
			State_SP <= 2'd0;
			// Trace: design.sv:5732:7
			AReg_DP <= 1'sb0;
			// Trace: design.sv:5733:7
			BReg_DP <= 1'sb0;
			// Trace: design.sv:5734:7
			ResReg_DP <= 1'sb0;
			// Trace: design.sv:5735:7
			Cnt_DP <= 1'sb0;
			// Trace: design.sv:5736:7
			RemSel_SP <= 1'b0;
			// Trace: design.sv:5737:7
			CompInv_SP <= 1'b0;
			// Trace: design.sv:5738:7
			ResInv_SP <= 1'b0;
		end
		else begin
			// Trace: design.sv:5740:7
			State_SP <= State_SN;
			// Trace: design.sv:5741:7
			AReg_DP <= AReg_DN;
			// Trace: design.sv:5742:7
			BReg_DP <= BReg_DN;
			// Trace: design.sv:5743:7
			ResReg_DP <= ResReg_DN;
			// Trace: design.sv:5744:7
			Cnt_DP <= Cnt_DN;
			// Trace: design.sv:5745:7
			RemSel_SP <= RemSel_SN;
			// Trace: design.sv:5746:7
			CompInv_SP <= CompInv_SN;
			// Trace: design.sv:5747:7
			ResInv_SP <= ResInv_SN;
		end
	end
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_ff_one (
	in_i,
	first_one_o,
	no_ones_o
);
	// Trace: design.sv:5788:15
	parameter LEN = 32;
	// Trace: design.sv:5790:5
	input wire [LEN - 1:0] in_i;
	// Trace: design.sv:5792:5
	output wire [$clog2(LEN) - 1:0] first_one_o;
	// Trace: design.sv:5793:5
	output wire no_ones_o;
	// Trace: design.sv:5796:3
	localparam NUM_LEVELS = $clog2(LEN);
	// Trace: design.sv:5798:3
	wire [(LEN * NUM_LEVELS) - 1:0] index_lut;
	// Trace: design.sv:5799:3
	wire [(2 ** NUM_LEVELS) - 1:0] sel_nodes;
	// Trace: design.sv:5800:3
	wire [((2 ** NUM_LEVELS) * NUM_LEVELS) - 1:0] index_nodes;
	// Trace: design.sv:5807:3
	// Trace: design.sv:5808:5
	genvar _gv_j_2;
	generate
		for (_gv_j_2 = 0; _gv_j_2 < LEN; _gv_j_2 = _gv_j_2 + 1) begin : gen_index_lut
			localparam j = _gv_j_2;
			// Trace: design.sv:5810:7
			assign index_lut[j * NUM_LEVELS+:NUM_LEVELS] = $unsigned(j);
		end
	endgenerate
	// Trace: design.sv:5814:3
	// Trace: design.sv:5815:5
	genvar _gv_k_2;
	// Trace: design.sv:5816:5
	genvar _gv_l_1;
	// Trace: design.sv:5817:5
	genvar _gv_level_1;
	generate
		for (_gv_level_1 = 0; _gv_level_1 < NUM_LEVELS; _gv_level_1 = _gv_level_1 + 1) begin : gen_tree
			localparam level = _gv_level_1;
			if (level < (NUM_LEVELS - 1)) begin : gen_non_root_level
				for (_gv_l_1 = 0; _gv_l_1 < (2 ** level); _gv_l_1 = _gv_l_1 + 1) begin : gen_node
					localparam l = _gv_l_1;
					// Trace: design.sv:5822:11
					assign sel_nodes[((2 ** level) - 1) + l] = sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] | sel_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) + 1];
					// Trace: design.sv:5823:11
					assign index_nodes[(((2 ** level) - 1) + l) * NUM_LEVELS+:NUM_LEVELS] = (sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] == 1'b1 ? index_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) * NUM_LEVELS+:NUM_LEVELS] : index_nodes[((((2 ** (level + 1)) - 1) + (l * 2)) + 1) * NUM_LEVELS+:NUM_LEVELS]);
				end
			end
			if (level == (NUM_LEVELS - 1)) begin : gen_root_level
				for (_gv_k_2 = 0; _gv_k_2 < (2 ** level); _gv_k_2 = _gv_k_2 + 1) begin : gen_node
					localparam k = _gv_k_2;
					if ((k * 2) < (LEN - 1)) begin : gen_two
						// Trace: design.sv:5832:13
						assign sel_nodes[((2 ** level) - 1) + k] = in_i[k * 2] | in_i[(k * 2) + 1];
						// Trace: design.sv:5833:13
						assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = (in_i[k * 2] == 1'b1 ? index_lut[(k * 2) * NUM_LEVELS+:NUM_LEVELS] : index_lut[((k * 2) + 1) * NUM_LEVELS+:NUM_LEVELS]);
					end
					if ((k * 2) == (LEN - 1)) begin : gen_one
						// Trace: design.sv:5837:13
						assign sel_nodes[((2 ** level) - 1) + k] = in_i[k * 2];
						// Trace: design.sv:5838:13
						assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = index_lut[(k * 2) * NUM_LEVELS+:NUM_LEVELS];
					end
					if ((k * 2) > (LEN - 1)) begin : gen_out_of_range
						// Trace: design.sv:5842:13
						assign sel_nodes[((2 ** level) - 1) + k] = 1'b0;
						// Trace: design.sv:5843:13
						assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = 1'sb0;
					end
				end
			end
		end
	endgenerate
	// Trace: design.sv:5855:3
	assign first_one_o = index_nodes[0+:NUM_LEVELS];
	// Trace: design.sv:5856:3
	assign no_ones_o = ~sel_nodes[0];
endmodule
module cv32e40p_popcnt (
	in_i,
	result_o
);
	// Trace: design.sv:5884:5
	input wire [31:0] in_i;
	// Trace: design.sv:5885:5
	output wire [5:0] result_o;
	// Trace: design.sv:5888:3
	wire [31:0] cnt_l1;
	// Trace: design.sv:5889:3
	wire [23:0] cnt_l2;
	// Trace: design.sv:5890:3
	wire [15:0] cnt_l3;
	// Trace: design.sv:5891:3
	wire [9:0] cnt_l4;
	// Trace: design.sv:5893:3
	genvar _gv_l_2;
	genvar _gv_m_2;
	genvar _gv_n_1;
	genvar _gv_p_1;
	// Trace: design.sv:5894:3
	generate
		for (_gv_l_2 = 0; _gv_l_2 < 16; _gv_l_2 = _gv_l_2 + 1) begin : gen_cnt_l1
			localparam l = _gv_l_2;
			// Trace: design.sv:5896:7
			assign cnt_l1[l * 2+:2] = {1'b0, in_i[2 * l]} + {1'b0, in_i[(2 * l) + 1]};
		end
	endgenerate
	// Trace: design.sv:5900:3
	generate
		for (_gv_m_2 = 0; _gv_m_2 < 8; _gv_m_2 = _gv_m_2 + 1) begin : gen_cnt_l2
			localparam m = _gv_m_2;
			// Trace: design.sv:5902:7
			assign cnt_l2[m * 3+:3] = {1'b0, cnt_l1[(2 * m) * 2+:2]} + {1'b0, cnt_l1[((2 * m) + 1) * 2+:2]};
		end
	endgenerate
	// Trace: design.sv:5906:3
	generate
		for (_gv_n_1 = 0; _gv_n_1 < 4; _gv_n_1 = _gv_n_1 + 1) begin : gen_cnt_l3
			localparam n = _gv_n_1;
			// Trace: design.sv:5908:7
			assign cnt_l3[n * 4+:4] = {1'b0, cnt_l2[(2 * n) * 3+:3]} + {1'b0, cnt_l2[((2 * n) + 1) * 3+:3]};
		end
	endgenerate
	// Trace: design.sv:5912:3
	generate
		for (_gv_p_1 = 0; _gv_p_1 < 2; _gv_p_1 = _gv_p_1 + 1) begin : gen_cnt_l4
			localparam p = _gv_p_1;
			// Trace: design.sv:5914:7
			assign cnt_l4[p * 5+:5] = {1'b0, cnt_l3[(2 * p) * 4+:4]} + {1'b0, cnt_l3[((2 * p) + 1) * 4+:4]};
		end
	endgenerate
	// Trace: design.sv:5918:3
	assign result_o = {1'b0, cnt_l4[0+:5]} + {1'b0, cnt_l4[5+:5]};
endmodule
module cv32e40p_compressed_decoder (
	instr_i,
	instr_o,
	is_compressed_o,
	illegal_instr_o
);
	reg _sv2v_0;
	// Trace: design.sv:5948:15
	parameter FPU = 0;
	// Trace: design.sv:5950:5
	input wire [31:0] instr_i;
	// Trace: design.sv:5951:5
	output reg [31:0] instr_o;
	// Trace: design.sv:5952:5
	output wire is_compressed_o;
	// Trace: design.sv:5953:5
	output reg illegal_instr_o;
	// Trace: design.sv:5956:3
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:5967:3
	localparam cv32e40p_pkg_OPCODE_BRANCH = 7'h63;
	localparam cv32e40p_pkg_OPCODE_JAL = 7'h6f;
	localparam cv32e40p_pkg_OPCODE_JALR = 7'h67;
	localparam cv32e40p_pkg_OPCODE_LOAD = 7'h03;
	localparam cv32e40p_pkg_OPCODE_LOAD_FP = 7'h07;
	localparam cv32e40p_pkg_OPCODE_LUI = 7'h37;
	localparam cv32e40p_pkg_OPCODE_OP = 7'h33;
	localparam cv32e40p_pkg_OPCODE_OPIMM = 7'h13;
	localparam cv32e40p_pkg_OPCODE_STORE = 7'h23;
	localparam cv32e40p_pkg_OPCODE_STORE_FP = 7'h27;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:5968:5
		illegal_instr_o = 1'b0;
		// Trace: design.sv:5969:5
		instr_o = 1'sb0;
		// Trace: design.sv:5971:5
		(* full_case, parallel_case *)
		case (instr_i[1:0])
			2'b00:
				// Trace: design.sv:5974:9
				(* full_case, parallel_case *)
				case (instr_i[15:13])
					3'b000: begin
						// Trace: design.sv:5977:13
						instr_o = {2'b00, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], cv32e40p_pkg_OPCODE_OPIMM};
						// Trace: design.sv:5990:13
						if (instr_i[12:5] == 8'b00000000)
							// Trace: design.sv:5990:40
							illegal_instr_o = 1'b1;
					end
					3'b001:
						// Trace: design.sv:5995:13
						if (FPU == 1)
							// Trace: design.sv:5996:15
							instr_o = {4'b0000, instr_i[6:5], instr_i[12:10], 5'b00001, instr_i[9:7], 5'b01101, instr_i[4:2], cv32e40p_pkg_OPCODE_LOAD_FP};
						else
							// Trace: design.sv:6008:18
							illegal_instr_o = 1'b1;
					3'b010:
						// Trace: design.sv:6013:13
						instr_o = {5'b00000, instr_i[5], instr_i[12:10], instr_i[6], 4'b0001, instr_i[9:7], 5'b01001, instr_i[4:2], cv32e40p_pkg_OPCODE_LOAD};
					3'b011:
						// Trace: design.sv:6030:13
						if (FPU == 1)
							// Trace: design.sv:6031:15
							instr_o = {5'b00000, instr_i[5], instr_i[12:10], instr_i[6], 4'b0001, instr_i[9:7], 5'b01001, instr_i[4:2], cv32e40p_pkg_OPCODE_LOAD_FP};
						else
							// Trace: design.sv:6044:18
							illegal_instr_o = 1'b1;
					3'b101:
						// Trace: design.sv:6049:13
						if (FPU == 1)
							// Trace: design.sv:6050:15
							instr_o = {4'b0000, instr_i[6:5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b011, instr_i[11:10], 3'b000, cv32e40p_pkg_OPCODE_STORE_FP};
						else
							// Trace: design.sv:6063:18
							illegal_instr_o = 1'b1;
					3'b110:
						// Trace: design.sv:6068:13
						instr_o = {5'b00000, instr_i[5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b010, instr_i[11:10], instr_i[6], 2'b00, cv32e40p_pkg_OPCODE_STORE};
					3'b111:
						// Trace: design.sv:6086:13
						if (FPU == 1)
							// Trace: design.sv:6087:15
							instr_o = {5'b00000, instr_i[5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b010, instr_i[11:10], instr_i[6], 2'b00, cv32e40p_pkg_OPCODE_STORE_FP};
						else
							// Trace: design.sv:6101:18
							illegal_instr_o = 1'b1;
					default:
						// Trace: design.sv:6104:13
						illegal_instr_o = 1'b1;
				endcase
			2'b01:
				// Trace: design.sv:6112:9
				(* full_case, parallel_case *)
				case (instr_i[15:13])
					3'b000:
						// Trace: design.sv:6116:13
						instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], cv32e40p_pkg_OPCODE_OPIMM};
					3'b001, 3'b101:
						// Trace: design.sv:6130:13
						instr_o = {instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], {9 {instr_i[12]}}, 4'b0000, ~instr_i[15], cv32e40p_pkg_OPCODE_JAL};
					3'b010:
						// Trace: design.sv:6147:13
						if (instr_i[11:7] == 5'b00000)
							// Trace: design.sv:6149:15
							instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 8'b00000000, instr_i[11:7], cv32e40p_pkg_OPCODE_OPIMM};
						else
							// Trace: design.sv:6154:15
							instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 8'b00000000, instr_i[11:7], cv32e40p_pkg_OPCODE_OPIMM};
					3'b011:
						// Trace: design.sv:6161:13
						if ({instr_i[12], instr_i[6:2]} == 6'b000000)
							// Trace: design.sv:6162:15
							illegal_instr_o = 1'b1;
						else
							// Trace: design.sv:6164:15
							if (instr_i[11:7] == 5'h02)
								// Trace: design.sv:6166:17
								instr_o = {{3 {instr_i[12]}}, instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 17'h00202, cv32e40p_pkg_OPCODE_OPIMM};
							else if (instr_i[11:7] == 5'b00000)
								// Trace: design.sv:6180:17
								instr_o = {{15 {instr_i[12]}}, instr_i[6:2], instr_i[11:7], cv32e40p_pkg_OPCODE_LUI};
							else
								// Trace: design.sv:6183:17
								instr_o = {{15 {instr_i[12]}}, instr_i[6:2], instr_i[11:7], cv32e40p_pkg_OPCODE_LUI};
					3'b100:
						// Trace: design.sv:6189:13
						(* full_case, parallel_case *)
						case (instr_i[11:10])
							2'b00, 2'b01:
								// Trace: design.sv:6193:17
								if (instr_i[12] == 1'b1) begin
									// Trace: design.sv:6195:19
									instr_o = {1'b0, instr_i[10], 5'b00000, instr_i[6:2], 2'b01, instr_i[9:7], 5'b10101, instr_i[9:7], cv32e40p_pkg_OPCODE_OPIMM};
									// Trace: design.sv:6207:19
									illegal_instr_o = 1'b1;
								end
								else
									// Trace: design.sv:6209:19
									if (instr_i[6:2] == 5'b00000)
										// Trace: design.sv:6211:21
										instr_o = {1'b0, instr_i[10], 5'b00000, instr_i[6:2], 2'b01, instr_i[9:7], 5'b10101, instr_i[9:7], cv32e40p_pkg_OPCODE_OPIMM};
									else
										// Trace: design.sv:6224:21
										instr_o = {1'b0, instr_i[10], 5'b00000, instr_i[6:2], 2'b01, instr_i[9:7], 5'b10101, instr_i[9:7], cv32e40p_pkg_OPCODE_OPIMM};
							2'b10:
								// Trace: design.sv:6242:17
								instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 2'b01, instr_i[9:7], 5'b11101, instr_i[9:7], cv32e40p_pkg_OPCODE_OPIMM};
							2'b11:
								// Trace: design.sv:6256:17
								(* full_case, parallel_case *)
								case ({instr_i[12], instr_i[6:5]})
									3'b000:
										// Trace: design.sv:6261:21
										instr_o = {9'b010000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b00001, instr_i[9:7], cv32e40p_pkg_OPCODE_OP};
									3'b001:
										// Trace: design.sv:6277:21
										instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b10001, instr_i[9:7], cv32e40p_pkg_OPCODE_OP};
									3'b010:
										// Trace: design.sv:6292:21
										instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b11001, instr_i[9:7], cv32e40p_pkg_OPCODE_OP};
									3'b011:
										// Trace: design.sv:6307:21
										instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b11101, instr_i[9:7], cv32e40p_pkg_OPCODE_OP};
									3'b100, 3'b101, 3'b110, 3'b111:
										// Trace: design.sv:6323:21
										illegal_instr_o = 1'b1;
								endcase
						endcase
					3'b110, 3'b111:
						// Trace: design.sv:6333:13
						instr_o = {{4 {instr_i[12]}}, instr_i[6:5], instr_i[2], 7'b0000001, instr_i[9:7], 2'b00, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], cv32e40p_pkg_OPCODE_BRANCH};
				endcase
			2'b10:
				// Trace: design.sv:6353:9
				(* full_case, parallel_case *)
				case (instr_i[15:13])
					3'b000:
						// Trace: design.sv:6355:13
						if (instr_i[12] == 1'b1) begin
							// Trace: design.sv:6357:15
							instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b001, instr_i[11:7], cv32e40p_pkg_OPCODE_OPIMM};
							// Trace: design.sv:6358:15
							illegal_instr_o = 1'b1;
						end
						else
							// Trace: design.sv:6360:15
							if ((instr_i[6:2] == 5'b00000) || (instr_i[11:7] == 5'b00000))
								// Trace: design.sv:6362:17
								instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b001, instr_i[11:7], cv32e40p_pkg_OPCODE_OPIMM};
							else
								// Trace: design.sv:6365:17
								instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b001, instr_i[11:7], cv32e40p_pkg_OPCODE_OPIMM};
					3'b001:
						// Trace: design.sv:6372:13
						if (FPU == 1)
							// Trace: design.sv:6373:15
							instr_o = {3'b000, instr_i[4:2], instr_i[12], instr_i[6:5], 11'h013, instr_i[11:7], cv32e40p_pkg_OPCODE_LOAD_FP};
						else
							// Trace: design.sv:6384:18
							illegal_instr_o = 1'b1;
					3'b010: begin
						// Trace: design.sv:6389:13
						instr_o = {4'b0000, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], cv32e40p_pkg_OPCODE_LOAD};
						// Trace: design.sv:6400:13
						if (instr_i[11:7] == 5'b00000)
							// Trace: design.sv:6400:40
							illegal_instr_o = 1'b1;
					end
					3'b011:
						// Trace: design.sv:6405:13
						if (FPU == 1)
							// Trace: design.sv:6406:15
							instr_o = {4'b0000, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], cv32e40p_pkg_OPCODE_LOAD_FP};
						else
							// Trace: design.sv:6417:18
							illegal_instr_o = 1'b1;
					3'b100:
						// Trace: design.sv:6421:13
						if (instr_i[12] == 1'b0) begin
							begin
								// Trace: design.sv:6422:15
								if (instr_i[6:2] == 5'b00000) begin
									// Trace: design.sv:6424:17
									instr_o = {12'b000000000000, instr_i[11:7], 8'b00000000, cv32e40p_pkg_OPCODE_JALR};
									// Trace: design.sv:6426:17
									if (instr_i[11:7] == 5'b00000)
										// Trace: design.sv:6426:44
										illegal_instr_o = 1'b1;
								end
								else
									// Trace: design.sv:6428:17
									if (instr_i[11:7] == 5'b00000)
										// Trace: design.sv:6430:19
										instr_o = {7'b0000000, instr_i[6:2], 8'b00000000, instr_i[11:7], cv32e40p_pkg_OPCODE_OP};
									else
										// Trace: design.sv:6433:19
										instr_o = {7'b0000000, instr_i[6:2], 8'b00000000, instr_i[11:7], cv32e40p_pkg_OPCODE_OP};
							end
						end
						else
							// Trace: design.sv:6437:15
							if (instr_i[6:2] == 5'b00000) begin
								begin
									// Trace: design.sv:6438:17
									if (instr_i[11:7] == 5'b00000)
										// Trace: design.sv:6440:19
										instr_o = 32'h00100073;
									else
										// Trace: design.sv:6443:19
										instr_o = {12'b000000000000, instr_i[11:7], 8'b00000001, cv32e40p_pkg_OPCODE_JALR};
								end
							end
							else
								// Trace: design.sv:6446:17
								if (instr_i[11:7] == 5'b00000)
									// Trace: design.sv:6448:19
									instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], cv32e40p_pkg_OPCODE_OP};
								else
									// Trace: design.sv:6451:19
									instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], cv32e40p_pkg_OPCODE_OP};
					3'b101:
						// Trace: design.sv:6459:13
						if (FPU == 1)
							// Trace: design.sv:6460:15
							instr_o = {3'b000, instr_i[9:7], instr_i[12], instr_i[6:2], 8'h13, instr_i[11:10], 3'b000, cv32e40p_pkg_OPCODE_STORE_FP};
						else
							// Trace: design.sv:6471:18
							illegal_instr_o = 1'b1;
					3'b110:
						// Trace: design.sv:6475:13
						instr_o = {4'b0000, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 2'b00, cv32e40p_pkg_OPCODE_STORE};
					3'b111:
						// Trace: design.sv:6490:13
						if (FPU == 1)
							// Trace: design.sv:6491:15
							instr_o = {4'b0000, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 2'b00, cv32e40p_pkg_OPCODE_STORE_FP};
						else
							// Trace: design.sv:6502:18
							illegal_instr_o = 1'b1;
				endcase
			default:
				// Trace: design.sv:6509:9
				instr_o = instr_i;
		endcase
	end
	// Trace: design.sv:6514:3
	assign is_compressed_o = instr_i[1:0] != 2'b11;
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_controller (
	clk,
	clk_ungated_i,
	rst_n,
	fetch_enable_i,
	ctrl_busy_o,
	is_decoding_o,
	is_fetch_failed_i,
	deassert_we_o,
	illegal_insn_i,
	ecall_insn_i,
	mret_insn_i,
	uret_insn_i,
	dret_insn_i,
	mret_dec_i,
	uret_dec_i,
	dret_dec_i,
	wfi_i,
	ebrk_insn_i,
	fencei_insn_i,
	csr_status_i,
	hwlp_mask_o,
	instr_valid_i,
	instr_req_o,
	pc_set_o,
	pc_mux_o,
	exc_pc_mux_o,
	trap_addr_mux_o,
	pc_id_i,
	is_compressed_i,
	hwlp_start_addr_i,
	hwlp_end_addr_i,
	hwlp_counter_i,
	hwlp_dec_cnt_o,
	hwlp_jump_o,
	hwlp_targ_addr_o,
	data_req_ex_i,
	data_we_ex_i,
	data_misaligned_i,
	data_load_event_i,
	data_err_i,
	data_err_ack_o,
	mult_multicycle_i,
	apu_en_i,
	apu_read_dep_i,
	apu_write_dep_i,
	apu_stall_o,
	branch_taken_ex_i,
	ctrl_transfer_insn_in_id_i,
	ctrl_transfer_insn_in_dec_i,
	irq_req_ctrl_i,
	irq_sec_ctrl_i,
	irq_id_ctrl_i,
	irq_wu_ctrl_i,
	current_priv_lvl_i,
	irq_ack_o,
	irq_id_o,
	exc_cause_o,
	debug_mode_o,
	debug_cause_o,
	debug_csr_save_o,
	debug_req_i,
	debug_single_step_i,
	debug_ebreakm_i,
	debug_ebreaku_i,
	trigger_match_i,
	debug_p_elw_no_sleep_o,
	debug_wfi_no_sleep_o,
	debug_havereset_o,
	debug_running_o,
	debug_halted_o,
	wake_from_sleep_o,
	csr_save_if_o,
	csr_save_id_o,
	csr_save_ex_o,
	csr_cause_o,
	csr_irq_sec_o,
	csr_restore_mret_id_o,
	csr_restore_uret_id_o,
	csr_restore_dret_id_o,
	csr_save_cause_o,
	regfile_we_id_i,
	regfile_alu_waddr_id_i,
	regfile_we_ex_i,
	regfile_waddr_ex_i,
	regfile_we_wb_i,
	regfile_alu_we_fw_i,
	operand_a_fw_mux_sel_o,
	operand_b_fw_mux_sel_o,
	operand_c_fw_mux_sel_o,
	reg_d_ex_is_reg_a_i,
	reg_d_ex_is_reg_b_i,
	reg_d_ex_is_reg_c_i,
	reg_d_wb_is_reg_a_i,
	reg_d_wb_is_reg_b_i,
	reg_d_wb_is_reg_c_i,
	reg_d_alu_is_reg_a_i,
	reg_d_alu_is_reg_b_i,
	reg_d_alu_is_reg_c_i,
	halt_if_o,
	halt_id_o,
	misaligned_stall_o,
	jr_stall_o,
	load_stall_o,
	id_ready_i,
	id_valid_i,
	ex_valid_i,
	wb_ready_i,
	perf_pipeline_stall_o
);
	reg _sv2v_0;
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:6549:13
	parameter PULP_CLUSTER = 0;
	// Trace: design.sv:6550:13
	parameter PULP_XPULP = 1;
	// Trace: design.sv:6553:3
	input wire clk;
	// Trace: design.sv:6554:3
	input wire clk_ungated_i;
	// Trace: design.sv:6555:3
	input wire rst_n;
	// Trace: design.sv:6557:3
	input wire fetch_enable_i;
	// Trace: design.sv:6558:3
	output reg ctrl_busy_o;
	// Trace: design.sv:6559:3
	output reg is_decoding_o;
	// Trace: design.sv:6560:3
	input wire is_fetch_failed_i;
	// Trace: design.sv:6563:3
	output reg deassert_we_o;
	// Trace: design.sv:6565:3
	input wire illegal_insn_i;
	// Trace: design.sv:6566:3
	input wire ecall_insn_i;
	// Trace: design.sv:6567:3
	input wire mret_insn_i;
	// Trace: design.sv:6568:3
	input wire uret_insn_i;
	// Trace: design.sv:6570:3
	input wire dret_insn_i;
	// Trace: design.sv:6572:3
	input wire mret_dec_i;
	// Trace: design.sv:6573:3
	input wire uret_dec_i;
	// Trace: design.sv:6574:3
	input wire dret_dec_i;
	// Trace: design.sv:6576:3
	input wire wfi_i;
	// Trace: design.sv:6577:3
	input wire ebrk_insn_i;
	// Trace: design.sv:6578:3
	input wire fencei_insn_i;
	// Trace: design.sv:6579:3
	input wire csr_status_i;
	// Trace: design.sv:6581:3
	output reg hwlp_mask_o;
	// Trace: design.sv:6584:3
	input wire instr_valid_i;
	// Trace: design.sv:6587:3
	output reg instr_req_o;
	// Trace: design.sv:6590:3
	output reg pc_set_o;
	// Trace: design.sv:6591:3
	output reg [3:0] pc_mux_o;
	// Trace: design.sv:6592:3
	output reg [2:0] exc_pc_mux_o;
	// Trace: design.sv:6593:3
	output reg [1:0] trap_addr_mux_o;
	// Trace: design.sv:6596:3
	input wire [31:0] pc_id_i;
	// Trace: design.sv:6597:3
	input wire is_compressed_i;
	// Trace: design.sv:6600:3
	input wire [63:0] hwlp_start_addr_i;
	// Trace: design.sv:6601:3
	input wire [63:0] hwlp_end_addr_i;
	// Trace: design.sv:6602:3
	input wire [63:0] hwlp_counter_i;
	// Trace: design.sv:6605:3
	output reg [1:0] hwlp_dec_cnt_o;
	// Trace: design.sv:6607:3
	output wire hwlp_jump_o;
	// Trace: design.sv:6608:3
	output reg [31:0] hwlp_targ_addr_o;
	// Trace: design.sv:6611:3
	input wire data_req_ex_i;
	// Trace: design.sv:6612:3
	input wire data_we_ex_i;
	// Trace: design.sv:6613:3
	input wire data_misaligned_i;
	// Trace: design.sv:6614:3
	input wire data_load_event_i;
	// Trace: design.sv:6615:3
	input wire data_err_i;
	// Trace: design.sv:6616:3
	output reg data_err_ack_o;
	// Trace: design.sv:6619:3
	input wire mult_multicycle_i;
	// Trace: design.sv:6622:3
	input wire apu_en_i;
	// Trace: design.sv:6623:3
	input wire apu_read_dep_i;
	// Trace: design.sv:6624:3
	input wire apu_write_dep_i;
	// Trace: design.sv:6626:3
	output wire apu_stall_o;
	// Trace: design.sv:6629:3
	input wire branch_taken_ex_i;
	// Trace: design.sv:6630:3
	input wire [1:0] ctrl_transfer_insn_in_id_i;
	// Trace: design.sv:6631:3
	input wire [1:0] ctrl_transfer_insn_in_dec_i;
	// Trace: design.sv:6634:3
	input wire irq_req_ctrl_i;
	// Trace: design.sv:6635:3
	input wire irq_sec_ctrl_i;
	// Trace: design.sv:6636:3
	input wire [4:0] irq_id_ctrl_i;
	// Trace: design.sv:6637:3
	input wire irq_wu_ctrl_i;
	// Trace: design.sv:6638:3
	// removed localparam type cv32e40p_pkg_PrivLvl_t
	input wire [1:0] current_priv_lvl_i;
	// Trace: design.sv:6640:3
	output reg irq_ack_o;
	// Trace: design.sv:6641:3
	output reg [4:0] irq_id_o;
	// Trace: design.sv:6643:3
	output reg [4:0] exc_cause_o;
	// Trace: design.sv:6646:3
	output wire debug_mode_o;
	// Trace: design.sv:6647:3
	output reg [2:0] debug_cause_o;
	// Trace: design.sv:6648:3
	output reg debug_csr_save_o;
	// Trace: design.sv:6649:3
	input wire debug_req_i;
	// Trace: design.sv:6650:3
	input wire debug_single_step_i;
	// Trace: design.sv:6651:3
	input wire debug_ebreakm_i;
	// Trace: design.sv:6652:3
	input wire debug_ebreaku_i;
	// Trace: design.sv:6653:3
	input wire trigger_match_i;
	// Trace: design.sv:6654:3
	output wire debug_p_elw_no_sleep_o;
	// Trace: design.sv:6655:3
	output wire debug_wfi_no_sleep_o;
	// Trace: design.sv:6656:3
	output wire debug_havereset_o;
	// Trace: design.sv:6657:3
	output wire debug_running_o;
	// Trace: design.sv:6658:3
	output wire debug_halted_o;
	// Trace: design.sv:6661:3
	output wire wake_from_sleep_o;
	// Trace: design.sv:6663:3
	output reg csr_save_if_o;
	// Trace: design.sv:6664:3
	output reg csr_save_id_o;
	// Trace: design.sv:6665:3
	output reg csr_save_ex_o;
	// Trace: design.sv:6666:3
	output reg [5:0] csr_cause_o;
	// Trace: design.sv:6667:3
	output reg csr_irq_sec_o;
	// Trace: design.sv:6668:3
	output reg csr_restore_mret_id_o;
	// Trace: design.sv:6669:3
	output reg csr_restore_uret_id_o;
	// Trace: design.sv:6671:3
	output reg csr_restore_dret_id_o;
	// Trace: design.sv:6673:3
	output reg csr_save_cause_o;
	// Trace: design.sv:6677:3
	input wire regfile_we_id_i;
	// Trace: design.sv:6678:3
	input wire [5:0] regfile_alu_waddr_id_i;
	// Trace: design.sv:6681:3
	input wire regfile_we_ex_i;
	// Trace: design.sv:6682:3
	input wire [5:0] regfile_waddr_ex_i;
	// Trace: design.sv:6683:3
	input wire regfile_we_wb_i;
	// Trace: design.sv:6684:3
	input wire regfile_alu_we_fw_i;
	// Trace: design.sv:6687:3
	output reg [1:0] operand_a_fw_mux_sel_o;
	// Trace: design.sv:6688:3
	output reg [1:0] operand_b_fw_mux_sel_o;
	// Trace: design.sv:6689:3
	output reg [1:0] operand_c_fw_mux_sel_o;
	// Trace: design.sv:6692:3
	input wire reg_d_ex_is_reg_a_i;
	// Trace: design.sv:6693:3
	input wire reg_d_ex_is_reg_b_i;
	// Trace: design.sv:6694:3
	input wire reg_d_ex_is_reg_c_i;
	// Trace: design.sv:6695:3
	input wire reg_d_wb_is_reg_a_i;
	// Trace: design.sv:6696:3
	input wire reg_d_wb_is_reg_b_i;
	// Trace: design.sv:6697:3
	input wire reg_d_wb_is_reg_c_i;
	// Trace: design.sv:6698:3
	input wire reg_d_alu_is_reg_a_i;
	// Trace: design.sv:6699:3
	input wire reg_d_alu_is_reg_b_i;
	// Trace: design.sv:6700:3
	input wire reg_d_alu_is_reg_c_i;
	// Trace: design.sv:6703:3
	output reg halt_if_o;
	// Trace: design.sv:6704:3
	output reg halt_id_o;
	// Trace: design.sv:6706:3
	output wire misaligned_stall_o;
	// Trace: design.sv:6707:3
	output reg jr_stall_o;
	// Trace: design.sv:6708:3
	output reg load_stall_o;
	// Trace: design.sv:6710:3
	input wire id_ready_i;
	// Trace: design.sv:6711:3
	input wire id_valid_i;
	// Trace: design.sv:6713:3
	input wire ex_valid_i;
	// Trace: design.sv:6715:3
	input wire wb_ready_i;
	// Trace: design.sv:6718:3
	output reg perf_pipeline_stall_o;
	// Trace: design.sv:6722:3
	// removed localparam type cv32e40p_pkg_ctrl_state_e
	reg [4:0] ctrl_fsm_cs;
	reg [4:0] ctrl_fsm_ns;
	// Trace: design.sv:6725:3
	// removed localparam type cv32e40p_pkg_debug_state_e
	reg [2:0] debug_fsm_cs;
	reg [2:0] debug_fsm_ns;
	// Trace: design.sv:6727:3
	reg jump_done;
	reg jump_done_q;
	reg jump_in_dec;
	reg branch_in_id_dec;
	reg branch_in_id;
	// Trace: design.sv:6729:3
	reg data_err_q;
	// Trace: design.sv:6731:3
	reg debug_mode_q;
	reg debug_mode_n;
	// Trace: design.sv:6732:3
	reg ebrk_force_debug_mode;
	// Trace: design.sv:6733:3
	reg is_hwlp_illegal;
	wire is_hwlp_body;
	// Trace: design.sv:6734:3
	reg illegal_insn_q;
	reg illegal_insn_n;
	// Trace: design.sv:6735:3
	reg debug_req_entry_q;
	reg debug_req_entry_n;
	// Trace: design.sv:6736:3
	reg debug_force_wakeup_q;
	reg debug_force_wakeup_n;
	// Trace: design.sv:6738:3
	wire hwlp_end0_eq_pc;
	// Trace: design.sv:6739:3
	wire hwlp_end1_eq_pc;
	// Trace: design.sv:6740:3
	wire hwlp_counter0_gt_1;
	// Trace: design.sv:6741:3
	wire hwlp_counter1_gt_1;
	// Trace: design.sv:6742:3
	wire hwlp_end0_eq_pc_plus4;
	// Trace: design.sv:6743:3
	wire hwlp_end1_eq_pc_plus4;
	// Trace: design.sv:6744:3
	wire hwlp_start0_leq_pc;
	// Trace: design.sv:6745:3
	wire hwlp_start1_leq_pc;
	// Trace: design.sv:6746:3
	wire hwlp_end0_geq_pc;
	// Trace: design.sv:6747:3
	wire hwlp_end1_geq_pc;
	// Trace: design.sv:6749:3
	reg hwlp_end_4_id_d;
	reg hwlp_end_4_id_q;
	// Trace: design.sv:6751:3
	reg debug_req_q;
	// Trace: design.sv:6752:3
	wire debug_req_pending;
	// Trace: design.sv:6755:3
	wire wfi_active;
	// Trace: design.sv:6767:3
	localparam cv32e40p_pkg_BRANCH_COND = 2'b11;
	localparam cv32e40p_pkg_BRANCH_JAL = 2'b01;
	localparam cv32e40p_pkg_BRANCH_JALR = 2'b10;
	localparam cv32e40p_pkg_DBG_CAUSE_EBREAK = 3'h1;
	localparam cv32e40p_pkg_DBG_CAUSE_HALTREQ = 3'h3;
	localparam cv32e40p_pkg_DBG_CAUSE_STEP = 3'h4;
	localparam cv32e40p_pkg_DBG_CAUSE_TRIGGER = 3'h2;
	localparam cv32e40p_pkg_EXC_CAUSE_BREAKPOINT = 5'h03;
	localparam cv32e40p_pkg_EXC_CAUSE_ECALL_MMODE = 5'h0b;
	localparam cv32e40p_pkg_EXC_CAUSE_ECALL_UMODE = 5'h08;
	localparam cv32e40p_pkg_EXC_CAUSE_ILLEGAL_INSN = 5'h02;
	localparam cv32e40p_pkg_EXC_CAUSE_INSTR_FAULT = 5'h01;
	localparam cv32e40p_pkg_EXC_CAUSE_LOAD_FAULT = 5'h05;
	localparam cv32e40p_pkg_EXC_CAUSE_STORE_FAULT = 5'h07;
	localparam cv32e40p_pkg_EXC_PC_DBD = 3'b010;
	localparam cv32e40p_pkg_EXC_PC_DBE = 3'b011;
	localparam cv32e40p_pkg_EXC_PC_EXCEPTION = 3'b000;
	localparam cv32e40p_pkg_EXC_PC_IRQ = 3'b001;
	localparam cv32e40p_pkg_PC_BOOT = 4'b0000;
	localparam cv32e40p_pkg_PC_BRANCH = 4'b0011;
	localparam cv32e40p_pkg_PC_DRET = 4'b0111;
	localparam cv32e40p_pkg_PC_EXCEPTION = 4'b0100;
	localparam cv32e40p_pkg_PC_FENCEI = 4'b0001;
	localparam cv32e40p_pkg_PC_HWLOOP = 4'b1000;
	localparam cv32e40p_pkg_PC_JUMP = 4'b0010;
	localparam cv32e40p_pkg_PC_MRET = 4'b0101;
	localparam cv32e40p_pkg_PC_URET = 4'b0110;
	localparam cv32e40p_pkg_TRAP_MACHINE = 2'b00;
	localparam cv32e40p_pkg_TRAP_USER = 2'b01;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:6771:5
		instr_req_o = 1'b1;
		// Trace: design.sv:6773:5
		data_err_ack_o = 1'b0;
		// Trace: design.sv:6775:5
		csr_save_if_o = 1'b0;
		// Trace: design.sv:6776:5
		csr_save_id_o = 1'b0;
		// Trace: design.sv:6777:5
		csr_save_ex_o = 1'b0;
		// Trace: design.sv:6778:5
		csr_restore_mret_id_o = 1'b0;
		// Trace: design.sv:6779:5
		csr_restore_uret_id_o = 1'b0;
		// Trace: design.sv:6781:5
		csr_restore_dret_id_o = 1'b0;
		// Trace: design.sv:6783:5
		csr_save_cause_o = 1'b0;
		// Trace: design.sv:6785:5
		exc_cause_o = 1'sb0;
		// Trace: design.sv:6786:5
		exc_pc_mux_o = cv32e40p_pkg_EXC_PC_IRQ;
		// Trace: design.sv:6787:5
		trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
		// Trace: design.sv:6789:5
		csr_cause_o = 1'sb0;
		// Trace: design.sv:6790:5
		csr_irq_sec_o = 1'b0;
		// Trace: design.sv:6792:5
		pc_mux_o = cv32e40p_pkg_PC_BOOT;
		// Trace: design.sv:6793:5
		pc_set_o = 1'b0;
		// Trace: design.sv:6794:5
		jump_done = jump_done_q;
		// Trace: design.sv:6796:5
		ctrl_fsm_ns = ctrl_fsm_cs;
		// Trace: design.sv:6798:5
		ctrl_busy_o = 1'b1;
		// Trace: design.sv:6800:5
		halt_if_o = 1'b0;
		// Trace: design.sv:6801:5
		halt_id_o = 1'b0;
		// Trace: design.sv:6802:5
		is_decoding_o = 1'b0;
		// Trace: design.sv:6803:5
		irq_ack_o = 1'b0;
		// Trace: design.sv:6804:5
		irq_id_o = 5'b00000;
		// Trace: design.sv:6806:5
		jump_in_dec = (ctrl_transfer_insn_in_dec_i == cv32e40p_pkg_BRANCH_JALR) || (ctrl_transfer_insn_in_dec_i == cv32e40p_pkg_BRANCH_JAL);
		// Trace: design.sv:6808:5
		branch_in_id = ctrl_transfer_insn_in_id_i == cv32e40p_pkg_BRANCH_COND;
		// Trace: design.sv:6809:5
		branch_in_id_dec = ctrl_transfer_insn_in_dec_i == cv32e40p_pkg_BRANCH_COND;
		// Trace: design.sv:6811:5
		ebrk_force_debug_mode = (debug_ebreakm_i && (current_priv_lvl_i == 2'b11)) || (debug_ebreaku_i && (current_priv_lvl_i == 2'b00));
		// Trace: design.sv:6813:5
		debug_csr_save_o = 1'b0;
		// Trace: design.sv:6814:5
		debug_cause_o = cv32e40p_pkg_DBG_CAUSE_EBREAK;
		// Trace: design.sv:6815:5
		debug_mode_n = debug_mode_q;
		// Trace: design.sv:6817:5
		illegal_insn_n = illegal_insn_q;
		// Trace: design.sv:6826:5
		debug_req_entry_n = debug_req_entry_q;
		// Trace: design.sv:6828:5
		debug_force_wakeup_n = debug_force_wakeup_q;
		// Trace: design.sv:6830:5
		perf_pipeline_stall_o = 1'b0;
		// Trace: design.sv:6832:5
		hwlp_mask_o = 1'b0;
		// Trace: design.sv:6834:5
		is_hwlp_illegal = 1'b0;
		// Trace: design.sv:6836:5
		hwlp_dec_cnt_o = 1'sb0;
		// Trace: design.sv:6837:5
		hwlp_end_4_id_d = 1'b0;
		// Trace: design.sv:6842:5
		hwlp_targ_addr_o = ((hwlp_start1_leq_pc && hwlp_end1_geq_pc) && !(hwlp_start0_leq_pc && hwlp_end0_geq_pc) ? hwlp_start_addr_i[32+:32] : hwlp_start_addr_i[0+:32]);
		// Trace: design.sv:6844:5
		(* full_case, parallel_case *)
		case (ctrl_fsm_cs)
			5'd0: begin
				// Trace: design.sv:6848:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:6849:9
				instr_req_o = 1'b0;
				// Trace: design.sv:6850:9
				if (fetch_enable_i == 1'b1)
					// Trace: design.sv:6852:11
					ctrl_fsm_ns = 5'd1;
			end
			5'd1: begin
				// Trace: design.sv:6859:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:6860:9
				instr_req_o = 1'b1;
				// Trace: design.sv:6861:9
				pc_mux_o = cv32e40p_pkg_PC_BOOT;
				// Trace: design.sv:6862:9
				pc_set_o = 1'b1;
				// Trace: design.sv:6863:9
				if (debug_req_pending) begin
					// Trace: design.sv:6864:13
					ctrl_fsm_ns = 5'd12;
					// Trace: design.sv:6865:13
					debug_force_wakeup_n = 1'b1;
				end
				else
					// Trace: design.sv:6867:13
					ctrl_fsm_ns = 5'd4;
			end
			5'd3: begin
				// Trace: design.sv:6873:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:6874:9
				ctrl_busy_o = 1'b0;
				// Trace: design.sv:6875:9
				instr_req_o = 1'b0;
				// Trace: design.sv:6876:9
				halt_if_o = 1'b1;
				// Trace: design.sv:6877:9
				halt_id_o = 1'b1;
				// Trace: design.sv:6878:9
				ctrl_fsm_ns = 5'd2;
			end
			5'd2: begin
				// Trace: design.sv:6886:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:6887:9
				instr_req_o = 1'b0;
				// Trace: design.sv:6888:9
				halt_if_o = 1'b1;
				// Trace: design.sv:6889:9
				halt_id_o = 1'b1;
				// Trace: design.sv:6893:9
				if (wake_from_sleep_o) begin
					begin
						// Trace: design.sv:6894:11
						if (debug_req_pending) begin
							// Trace: design.sv:6895:15
							ctrl_fsm_ns = 5'd12;
							// Trace: design.sv:6896:15
							debug_force_wakeup_n = 1'b1;
						end
						else
							// Trace: design.sv:6898:15
							ctrl_fsm_ns = 5'd4;
					end
				end
				else
					// Trace: design.sv:6901:11
					ctrl_busy_o = 1'b0;
			end
			5'd4: begin
				// Trace: design.sv:6907:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:6910:9
				ctrl_fsm_ns = 5'd5;
				// Trace: design.sv:6913:9
				if (irq_req_ctrl_i && ~(debug_req_pending || debug_mode_q)) begin
					// Trace: design.sv:6919:11
					halt_if_o = 1'b1;
					// Trace: design.sv:6920:11
					halt_id_o = 1'b1;
					// Trace: design.sv:6922:11
					pc_set_o = 1'b1;
					// Trace: design.sv:6923:11
					pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
					// Trace: design.sv:6924:11
					exc_pc_mux_o = cv32e40p_pkg_EXC_PC_IRQ;
					// Trace: design.sv:6925:11
					exc_cause_o = irq_id_ctrl_i;
					// Trace: design.sv:6926:11
					csr_irq_sec_o = irq_sec_ctrl_i;
					// Trace: design.sv:6929:11
					irq_ack_o = 1'b1;
					// Trace: design.sv:6930:11
					irq_id_o = irq_id_ctrl_i;
					// Trace: design.sv:6932:11
					if (irq_sec_ctrl_i)
						// Trace: design.sv:6933:13
						trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
					else
						// Trace: design.sv:6935:13
						trap_addr_mux_o = (current_priv_lvl_i == 2'b00 ? cv32e40p_pkg_TRAP_USER : cv32e40p_pkg_TRAP_MACHINE);
					// Trace: design.sv:6937:11
					csr_save_cause_o = 1'b1;
					// Trace: design.sv:6938:11
					csr_cause_o = {1'b1, irq_id_ctrl_i};
					// Trace: design.sv:6939:11
					csr_save_if_o = 1'b1;
				end
			end
			5'd5:
				// Trace: design.sv:6946:11
				if (branch_taken_ex_i) begin
					// Trace: design.sv:6950:13
					is_decoding_o = 1'b0;
					// Trace: design.sv:6952:13
					pc_mux_o = cv32e40p_pkg_PC_BRANCH;
					// Trace: design.sv:6953:13
					pc_set_o = 1'b1;
				end
				else if (data_err_i) begin
					// Trace: design.sv:6965:13
					is_decoding_o = 1'b0;
					// Trace: design.sv:6966:13
					halt_if_o = 1'b1;
					// Trace: design.sv:6967:13
					halt_id_o = 1'b1;
					// Trace: design.sv:6968:13
					csr_save_ex_o = 1'b1;
					// Trace: design.sv:6969:13
					csr_save_cause_o = 1'b1;
					// Trace: design.sv:6970:13
					data_err_ack_o = 1'b1;
					// Trace: design.sv:6973:13
					csr_cause_o = {1'b0, (data_we_ex_i ? cv32e40p_pkg_EXC_CAUSE_STORE_FAULT : cv32e40p_pkg_EXC_CAUSE_LOAD_FAULT)};
					// Trace: design.sv:6974:13
					ctrl_fsm_ns = 5'd9;
				end
				else if (is_fetch_failed_i) begin
					// Trace: design.sv:6983:13
					is_decoding_o = 1'b0;
					// Trace: design.sv:6984:13
					halt_id_o = 1'b1;
					// Trace: design.sv:6985:13
					halt_if_o = 1'b1;
					// Trace: design.sv:6986:13
					csr_save_if_o = 1'b1;
					// Trace: design.sv:6987:13
					csr_save_cause_o = !debug_mode_q;
					// Trace: design.sv:6991:13
					csr_cause_o = {1'b0, cv32e40p_pkg_EXC_CAUSE_INSTR_FAULT};
					// Trace: design.sv:6992:13
					ctrl_fsm_ns = 5'd9;
				end
				else if (instr_valid_i) begin : blk_decode_level1
					// Trace: design.sv:7002:13
					is_decoding_o = 1'b1;
					// Trace: design.sv:7003:13
					illegal_insn_n = 1'b0;
					// Trace: design.sv:7005:13
					if ((debug_req_pending || trigger_match_i) & ~debug_mode_q) begin
						// Trace: design.sv:7008:17
						halt_if_o = 1'b1;
						// Trace: design.sv:7009:17
						halt_id_o = 1'b1;
						// Trace: design.sv:7010:17
						ctrl_fsm_ns = 5'd13;
						// Trace: design.sv:7011:17
						debug_req_entry_n = 1'b1;
					end
					else if (irq_req_ctrl_i && ~debug_mode_q) begin
						// Trace: design.sv:7016:17
						hwlp_mask_o = (PULP_XPULP ? 1'b1 : 1'b0);
						// Trace: design.sv:7018:17
						is_decoding_o = 1'b0;
						// Trace: design.sv:7019:17
						halt_if_o = 1'b1;
						// Trace: design.sv:7020:17
						halt_id_o = 1'b1;
						// Trace: design.sv:7022:17
						pc_set_o = 1'b1;
						// Trace: design.sv:7023:17
						pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
						// Trace: design.sv:7024:17
						exc_pc_mux_o = cv32e40p_pkg_EXC_PC_IRQ;
						// Trace: design.sv:7025:17
						exc_cause_o = irq_id_ctrl_i;
						// Trace: design.sv:7026:17
						csr_irq_sec_o = irq_sec_ctrl_i;
						// Trace: design.sv:7029:17
						irq_ack_o = 1'b1;
						// Trace: design.sv:7030:17
						irq_id_o = irq_id_ctrl_i;
						// Trace: design.sv:7032:17
						if (irq_sec_ctrl_i)
							// Trace: design.sv:7033:19
							trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
						else
							// Trace: design.sv:7035:19
							trap_addr_mux_o = (current_priv_lvl_i == 2'b00 ? cv32e40p_pkg_TRAP_USER : cv32e40p_pkg_TRAP_MACHINE);
						// Trace: design.sv:7037:17
						csr_save_cause_o = 1'b1;
						// Trace: design.sv:7038:17
						csr_cause_o = {1'b1, irq_id_ctrl_i};
						// Trace: design.sv:7039:17
						csr_save_id_o = 1'b1;
					end
					else begin
						// Trace: design.sv:7044:17
						is_hwlp_illegal = is_hwlp_body & (((((((jump_in_dec || branch_in_id_dec) || mret_insn_i) || uret_insn_i) || dret_insn_i) || is_compressed_i) || fencei_insn_i) || wfi_active);
						// Trace: design.sv:7046:17
						if (illegal_insn_i || is_hwlp_illegal) begin
							// Trace: design.sv:7048:19
							halt_if_o = 1'b1;
							// Trace: design.sv:7049:19
							halt_id_o = 1'b0;
							// Trace: design.sv:7050:19
							ctrl_fsm_ns = (id_ready_i ? 5'd8 : 5'd5);
							// Trace: design.sv:7051:19
							illegal_insn_n = 1'b1;
						end
						else
							// Trace: design.sv:7056:19
							(* full_case, parallel_case *)
							case (1'b1)
								jump_in_dec: begin
									// Trace: design.sv:7063:23
									pc_mux_o = cv32e40p_pkg_PC_JUMP;
									// Trace: design.sv:7065:23
									if (~jr_stall_o && ~jump_done_q) begin
										// Trace: design.sv:7066:25
										pc_set_o = 1'b1;
										// Trace: design.sv:7067:25
										jump_done = 1'b1;
									end
								end
								ebrk_insn_i: begin
									// Trace: design.sv:7072:23
									halt_if_o = 1'b1;
									// Trace: design.sv:7073:23
									halt_id_o = 1'b0;
									// Trace: design.sv:7075:23
									if (debug_mode_q)
										// Trace: design.sv:7077:25
										ctrl_fsm_ns = 5'd13;
									else if (ebrk_force_debug_mode)
										// Trace: design.sv:7081:25
										ctrl_fsm_ns = 5'd13;
									else
										// Trace: design.sv:7084:25
										ctrl_fsm_ns = (id_ready_i ? 5'd8 : 5'd5);
								end
								wfi_active: begin
									// Trace: design.sv:7090:23
									halt_if_o = 1'b1;
									// Trace: design.sv:7091:23
									halt_id_o = 1'b0;
									// Trace: design.sv:7092:23
									ctrl_fsm_ns = (id_ready_i ? 5'd8 : 5'd5);
								end
								ecall_insn_i: begin
									// Trace: design.sv:7096:23
									halt_if_o = 1'b1;
									// Trace: design.sv:7097:23
									halt_id_o = 1'b0;
									// Trace: design.sv:7098:23
									ctrl_fsm_ns = (id_ready_i ? 5'd8 : 5'd5);
								end
								fencei_insn_i: begin
									// Trace: design.sv:7102:23
									halt_if_o = 1'b1;
									// Trace: design.sv:7103:23
									halt_id_o = 1'b0;
									// Trace: design.sv:7104:23
									ctrl_fsm_ns = (id_ready_i ? 5'd8 : 5'd5);
								end
								(mret_insn_i | uret_insn_i) | dret_insn_i: begin
									// Trace: design.sv:7108:23
									halt_if_o = 1'b1;
									// Trace: design.sv:7109:23
									halt_id_o = 1'b0;
									// Trace: design.sv:7110:23
									ctrl_fsm_ns = (id_ready_i ? 5'd8 : 5'd5);
								end
								csr_status_i: begin
									// Trace: design.sv:7114:23
									halt_if_o = 1'b1;
									// Trace: design.sv:7115:23
									ctrl_fsm_ns = (id_ready_i ? 5'd8 : 5'd5);
								end
								data_load_event_i: begin
									// Trace: design.sv:7119:23
									ctrl_fsm_ns = (id_ready_i ? 5'd7 : 5'd5);
									// Trace: design.sv:7120:23
									halt_if_o = 1'b1;
								end
								default:
									// Trace: design.sv:7125:23
									if (is_hwlp_body) begin
										// Trace: design.sv:7132:25
										ctrl_fsm_ns = (hwlp_end0_eq_pc_plus4 || hwlp_end1_eq_pc_plus4 ? 5'd5 : 5'd15);
										// Trace: design.sv:7135:25
										if (hwlp_end0_eq_pc && hwlp_counter0_gt_1) begin
											// Trace: design.sv:7136:29
											pc_mux_o = cv32e40p_pkg_PC_HWLOOP;
											// Trace: design.sv:7137:29
											if (~jump_done_q) begin
												// Trace: design.sv:7138:31
												pc_set_o = 1'b1;
												// Trace: design.sv:7141:31
												jump_done = 1'b1;
												// Trace: design.sv:7142:31
												hwlp_dec_cnt_o[0] = 1'b1;
											end
										end
										if (hwlp_end1_eq_pc && hwlp_counter1_gt_1) begin
											// Trace: design.sv:7146:29
											pc_mux_o = cv32e40p_pkg_PC_HWLOOP;
											// Trace: design.sv:7147:29
											if (~jump_done_q) begin
												// Trace: design.sv:7148:31
												pc_set_o = 1'b1;
												// Trace: design.sv:7151:31
												jump_done = 1'b1;
												// Trace: design.sv:7152:31
												hwlp_dec_cnt_o[1] = 1'b1;
											end
										end
									end
							endcase
						if (debug_single_step_i & ~debug_mode_q) begin
							// Trace: design.sv:7163:21
							halt_if_o = 1'b1;
							// Trace: design.sv:7172:21
							if (id_ready_i)
								// Trace: design.sv:7174:25
								(* full_case, parallel_case *)
								case (1'b1)
									illegal_insn_i | ecall_insn_i:
										// Trace: design.sv:7178:29
										ctrl_fsm_ns = 5'd8;
									~ebrk_force_debug_mode & ebrk_insn_i:
										// Trace: design.sv:7183:29
										ctrl_fsm_ns = 5'd8;
									mret_insn_i | uret_insn_i:
										// Trace: design.sv:7188:29
										ctrl_fsm_ns = 5'd8;
									branch_in_id:
										// Trace: design.sv:7193:29
										ctrl_fsm_ns = 5'd14;
									default:
										// Trace: design.sv:7198:29
										ctrl_fsm_ns = 5'd13;
								endcase
						end
					end
				end
				else begin
					// Trace: design.sv:7207:13
					is_decoding_o = 1'b0;
					// Trace: design.sv:7208:13
					perf_pipeline_stall_o = data_load_event_i;
				end
			5'd15:
				// Trace: design.sv:7214:9
				if (PULP_XPULP) begin
					begin
						// Trace: design.sv:7215:11
						if (instr_valid_i) begin
							// Trace: design.sv:7218:13
							is_decoding_o = 1'b1;
							// Trace: design.sv:7220:13
							if ((debug_req_pending || trigger_match_i) & ~debug_mode_q) begin
								// Trace: design.sv:7223:17
								halt_if_o = 1'b1;
								// Trace: design.sv:7224:17
								halt_id_o = 1'b1;
								// Trace: design.sv:7225:17
								ctrl_fsm_ns = 5'd13;
								// Trace: design.sv:7226:17
								debug_req_entry_n = 1'b1;
							end
							else if (irq_req_ctrl_i && ~debug_mode_q) begin
								// Trace: design.sv:7231:17
								hwlp_mask_o = (PULP_XPULP ? 1'b1 : 1'b0);
								// Trace: design.sv:7233:17
								is_decoding_o = 1'b0;
								// Trace: design.sv:7234:17
								halt_if_o = 1'b1;
								// Trace: design.sv:7235:17
								halt_id_o = 1'b1;
								// Trace: design.sv:7237:17
								pc_set_o = 1'b1;
								// Trace: design.sv:7238:17
								pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
								// Trace: design.sv:7239:17
								exc_pc_mux_o = cv32e40p_pkg_EXC_PC_IRQ;
								// Trace: design.sv:7240:17
								exc_cause_o = irq_id_ctrl_i;
								// Trace: design.sv:7241:17
								csr_irq_sec_o = irq_sec_ctrl_i;
								// Trace: design.sv:7244:17
								irq_ack_o = 1'b1;
								// Trace: design.sv:7245:17
								irq_id_o = irq_id_ctrl_i;
								// Trace: design.sv:7247:17
								if (irq_sec_ctrl_i)
									// Trace: design.sv:7248:19
									trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
								else
									// Trace: design.sv:7250:19
									trap_addr_mux_o = (current_priv_lvl_i == 2'b00 ? cv32e40p_pkg_TRAP_USER : cv32e40p_pkg_TRAP_MACHINE);
								// Trace: design.sv:7252:17
								csr_save_cause_o = 1'b1;
								// Trace: design.sv:7253:17
								csr_cause_o = {1'b1, irq_id_ctrl_i};
								// Trace: design.sv:7254:17
								csr_save_id_o = 1'b1;
								// Trace: design.sv:7256:17
								ctrl_fsm_ns = 5'd5;
							end
							else begin
								// Trace: design.sv:7261:17
								is_hwlp_illegal = ((((((jump_in_dec || branch_in_id_dec) || mret_insn_i) || uret_insn_i) || dret_insn_i) || is_compressed_i) || fencei_insn_i) || wfi_active;
								// Trace: design.sv:7263:17
								if (illegal_insn_i || is_hwlp_illegal) begin
									// Trace: design.sv:7265:19
									halt_if_o = 1'b1;
									// Trace: design.sv:7266:19
									halt_id_o = 1'b1;
									// Trace: design.sv:7267:19
									ctrl_fsm_ns = 5'd8;
									// Trace: design.sv:7268:19
									illegal_insn_n = 1'b1;
								end
								else
									// Trace: design.sv:7273:19
									(* full_case, parallel_case *)
									case (1'b1)
										ebrk_insn_i: begin
											// Trace: design.sv:7276:23
											halt_if_o = 1'b1;
											// Trace: design.sv:7277:23
											halt_id_o = 1'b1;
											// Trace: design.sv:7279:23
											if (debug_mode_q)
												// Trace: design.sv:7281:25
												ctrl_fsm_ns = 5'd13;
											else if (ebrk_force_debug_mode)
												// Trace: design.sv:7285:25
												ctrl_fsm_ns = 5'd13;
											else
												// Trace: design.sv:7289:25
												ctrl_fsm_ns = 5'd8;
										end
										ecall_insn_i: begin
											// Trace: design.sv:7295:23
											halt_if_o = 1'b1;
											// Trace: design.sv:7296:23
											halt_id_o = 1'b1;
											// Trace: design.sv:7297:23
											ctrl_fsm_ns = 5'd8;
										end
										csr_status_i: begin
											// Trace: design.sv:7301:23
											halt_if_o = 1'b1;
											// Trace: design.sv:7302:23
											ctrl_fsm_ns = (id_ready_i ? 5'd8 : 5'd15);
										end
										data_load_event_i: begin
											// Trace: design.sv:7306:23
											ctrl_fsm_ns = (id_ready_i ? 5'd7 : 5'd15);
											// Trace: design.sv:7307:23
											halt_if_o = 1'b1;
										end
										default: begin
											// Trace: design.sv:7313:23
											if (hwlp_end1_eq_pc_plus4) begin
												begin
													// Trace: design.sv:7314:27
													if (hwlp_counter1_gt_1) begin
														// Trace: design.sv:7315:29
														hwlp_end_4_id_d = 1'b1;
														// Trace: design.sv:7316:29
														hwlp_targ_addr_o = hwlp_start_addr_i[32+:32];
														// Trace: design.sv:7317:29
														ctrl_fsm_ns = 5'd15;
													end
													else
														// Trace: design.sv:7319:29
														ctrl_fsm_ns = (is_hwlp_body ? 5'd15 : 5'd5);
												end
											end
											if (hwlp_end0_eq_pc_plus4) begin
												begin
													// Trace: design.sv:7323:27
													if (hwlp_counter0_gt_1) begin
														// Trace: design.sv:7324:29
														hwlp_end_4_id_d = 1'b1;
														// Trace: design.sv:7325:29
														hwlp_targ_addr_o = hwlp_start_addr_i[0+:32];
														// Trace: design.sv:7326:29
														ctrl_fsm_ns = 5'd15;
													end
													else
														// Trace: design.sv:7328:29
														ctrl_fsm_ns = (is_hwlp_body ? 5'd15 : 5'd5);
												end
											end
											// Trace: design.sv:7331:23
											hwlp_dec_cnt_o[0] = hwlp_end0_eq_pc;
											// Trace: design.sv:7332:23
											hwlp_dec_cnt_o[1] = hwlp_end1_eq_pc;
										end
									endcase
								if (debug_single_step_i & ~debug_mode_q) begin
									// Trace: design.sv:7340:21
									halt_if_o = 1'b1;
									// Trace: design.sv:7349:21
									if (id_ready_i)
										// Trace: design.sv:7351:25
										(* full_case, parallel_case *)
										case (1'b1)
											illegal_insn_i | ecall_insn_i:
												// Trace: design.sv:7355:29
												ctrl_fsm_ns = 5'd8;
											~ebrk_force_debug_mode & ebrk_insn_i:
												// Trace: design.sv:7360:29
												ctrl_fsm_ns = 5'd8;
											mret_insn_i | uret_insn_i:
												// Trace: design.sv:7365:29
												ctrl_fsm_ns = 5'd8;
											branch_in_id:
												// Trace: design.sv:7370:29
												ctrl_fsm_ns = 5'd14;
											default:
												// Trace: design.sv:7375:29
												ctrl_fsm_ns = 5'd13;
										endcase
								end
							end
						end
						else begin
							// Trace: design.sv:7384:13
							is_decoding_o = 1'b0;
							// Trace: design.sv:7385:13
							perf_pipeline_stall_o = data_load_event_i;
						end
					end
				end
			5'd8: begin
				// Trace: design.sv:7393:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:7395:9
				halt_if_o = 1'b1;
				// Trace: design.sv:7396:9
				halt_id_o = 1'b1;
				// Trace: design.sv:7398:9
				if (data_err_i) begin
					// Trace: design.sv:7401:13
					csr_save_ex_o = 1'b1;
					// Trace: design.sv:7402:13
					csr_save_cause_o = 1'b1;
					// Trace: design.sv:7403:13
					data_err_ack_o = 1'b1;
					// Trace: design.sv:7405:13
					csr_cause_o = {1'b0, (data_we_ex_i ? cv32e40p_pkg_EXC_CAUSE_STORE_FAULT : cv32e40p_pkg_EXC_CAUSE_LOAD_FAULT)};
					// Trace: design.sv:7406:13
					ctrl_fsm_ns = 5'd9;
					// Trace: design.sv:7409:13
					illegal_insn_n = 1'b0;
				end
				else if (ex_valid_i) begin
					// Trace: design.sv:7413:11
					ctrl_fsm_ns = 5'd9;
					// Trace: design.sv:7415:11
					if (illegal_insn_q) begin
						// Trace: design.sv:7416:13
						csr_save_id_o = 1'b1;
						// Trace: design.sv:7417:13
						csr_save_cause_o = !debug_mode_q;
						// Trace: design.sv:7418:13
						csr_cause_o = {1'b0, cv32e40p_pkg_EXC_CAUSE_ILLEGAL_INSN};
					end
					else
						// Trace: design.sv:7420:13
						(* full_case, parallel_case *)
						case (1'b1)
							ebrk_insn_i: begin
								// Trace: design.sv:7422:17
								csr_save_id_o = 1'b1;
								// Trace: design.sv:7423:17
								csr_save_cause_o = 1'b1;
								// Trace: design.sv:7424:17
								csr_cause_o = {1'b0, cv32e40p_pkg_EXC_CAUSE_BREAKPOINT};
							end
							ecall_insn_i: begin
								// Trace: design.sv:7427:17
								csr_save_id_o = 1'b1;
								// Trace: design.sv:7428:17
								csr_save_cause_o = !debug_mode_q;
								// Trace: design.sv:7429:17
								csr_cause_o = {1'b0, (current_priv_lvl_i == 2'b00 ? cv32e40p_pkg_EXC_CAUSE_ECALL_UMODE : cv32e40p_pkg_EXC_CAUSE_ECALL_MMODE)};
							end
							default:
								;
						endcase
				end
			end
			5'd6:
				// Trace: design.sv:7440:9
				if (PULP_CLUSTER == 1'b1) begin
					// Trace: design.sv:7441:11
					is_decoding_o = 1'b0;
					// Trace: design.sv:7443:11
					halt_if_o = 1'b1;
					// Trace: design.sv:7444:11
					halt_id_o = 1'b1;
					// Trace: design.sv:7446:11
					ctrl_fsm_ns = 5'd5;
					// Trace: design.sv:7448:11
					perf_pipeline_stall_o = data_load_event_i;
					// Trace: design.sv:7450:11
					if (irq_req_ctrl_i && ~(debug_req_pending || debug_mode_q)) begin
						// Trace: design.sv:7452:13
						is_decoding_o = 1'b0;
						// Trace: design.sv:7453:13
						halt_if_o = 1'b1;
						// Trace: design.sv:7454:13
						halt_id_o = 1'b1;
						// Trace: design.sv:7456:13
						pc_set_o = 1'b1;
						// Trace: design.sv:7457:13
						pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
						// Trace: design.sv:7458:13
						exc_pc_mux_o = cv32e40p_pkg_EXC_PC_IRQ;
						// Trace: design.sv:7459:13
						exc_cause_o = irq_id_ctrl_i;
						// Trace: design.sv:7460:13
						csr_irq_sec_o = irq_sec_ctrl_i;
						// Trace: design.sv:7463:13
						irq_ack_o = 1'b1;
						// Trace: design.sv:7464:13
						irq_id_o = irq_id_ctrl_i;
						// Trace: design.sv:7466:13
						if (irq_sec_ctrl_i)
							// Trace: design.sv:7467:15
							trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
						else
							// Trace: design.sv:7469:15
							trap_addr_mux_o = (current_priv_lvl_i == 2'b00 ? cv32e40p_pkg_TRAP_USER : cv32e40p_pkg_TRAP_MACHINE);
						// Trace: design.sv:7471:13
						csr_save_cause_o = 1'b1;
						// Trace: design.sv:7472:13
						csr_cause_o = {1'b1, irq_id_ctrl_i};
						// Trace: design.sv:7473:13
						csr_save_id_o = 1'b1;
					end
				end
			5'd7:
				// Trace: design.sv:7480:9
				if (PULP_CLUSTER == 1'b1) begin
					// Trace: design.sv:7481:11
					is_decoding_o = 1'b0;
					// Trace: design.sv:7483:11
					halt_if_o = 1'b1;
					// Trace: design.sv:7484:11
					halt_id_o = 1'b1;
					// Trace: design.sv:7491:11
					if (id_ready_i)
						// Trace: design.sv:7492:13
						ctrl_fsm_ns = ((debug_req_pending || trigger_match_i) & ~debug_mode_q ? 5'd13 : 5'd6);
					else
						// Trace: design.sv:7496:13
						ctrl_fsm_ns = 5'd7;
					// Trace: design.sv:7498:11
					perf_pipeline_stall_o = data_load_event_i;
				end
			5'd9: begin
				// Trace: design.sv:7505:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:7507:9
				halt_if_o = 1'b1;
				// Trace: design.sv:7508:9
				halt_id_o = 1'b1;
				// Trace: design.sv:7510:9
				ctrl_fsm_ns = 5'd5;
				// Trace: design.sv:7512:9
				if (data_err_q) begin
					// Trace: design.sv:7514:13
					pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
					// Trace: design.sv:7515:13
					pc_set_o = 1'b1;
					// Trace: design.sv:7516:13
					trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
					// Trace: design.sv:7518:13
					exc_pc_mux_o = cv32e40p_pkg_EXC_PC_EXCEPTION;
					// Trace: design.sv:7519:13
					exc_cause_o = (data_we_ex_i ? cv32e40p_pkg_EXC_CAUSE_LOAD_FAULT : cv32e40p_pkg_EXC_CAUSE_STORE_FAULT);
				end
				else if (is_fetch_failed_i) begin
					// Trace: design.sv:7524:13
					pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
					// Trace: design.sv:7525:13
					pc_set_o = 1'b1;
					// Trace: design.sv:7526:13
					trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
					// Trace: design.sv:7527:13
					exc_pc_mux_o = (debug_mode_q ? cv32e40p_pkg_EXC_PC_DBE : cv32e40p_pkg_EXC_PC_EXCEPTION);
					// Trace: design.sv:7528:13
					exc_cause_o = cv32e40p_pkg_EXC_CAUSE_INSTR_FAULT;
				end
				else
					// Trace: design.sv:7532:11
					if (illegal_insn_q) begin
						// Trace: design.sv:7534:15
						pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
						// Trace: design.sv:7535:15
						pc_set_o = 1'b1;
						// Trace: design.sv:7536:15
						trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
						// Trace: design.sv:7537:15
						exc_pc_mux_o = (debug_mode_q ? cv32e40p_pkg_EXC_PC_DBE : cv32e40p_pkg_EXC_PC_EXCEPTION);
						// Trace: design.sv:7538:15
						illegal_insn_n = 1'b0;
						// Trace: design.sv:7539:15
						if (debug_single_step_i && ~debug_mode_q)
							// Trace: design.sv:7540:19
							ctrl_fsm_ns = 5'd12;
					end
					else
						// Trace: design.sv:7542:13
						(* full_case, parallel_case *)
						case (1'b1)
							ebrk_insn_i: begin
								// Trace: design.sv:7545:19
								pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
								// Trace: design.sv:7546:19
								pc_set_o = 1'b1;
								// Trace: design.sv:7547:19
								trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
								// Trace: design.sv:7548:19
								exc_pc_mux_o = cv32e40p_pkg_EXC_PC_EXCEPTION;
								// Trace: design.sv:7550:19
								if (debug_single_step_i && ~debug_mode_q)
									// Trace: design.sv:7551:23
									ctrl_fsm_ns = 5'd12;
							end
							ecall_insn_i: begin
								// Trace: design.sv:7555:19
								pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
								// Trace: design.sv:7556:19
								pc_set_o = 1'b1;
								// Trace: design.sv:7557:19
								trap_addr_mux_o = cv32e40p_pkg_TRAP_MACHINE;
								// Trace: design.sv:7558:19
								exc_pc_mux_o = (debug_mode_q ? cv32e40p_pkg_EXC_PC_DBE : cv32e40p_pkg_EXC_PC_EXCEPTION);
								// Trace: design.sv:7560:19
								if (debug_single_step_i && ~debug_mode_q)
									// Trace: design.sv:7561:23
									ctrl_fsm_ns = 5'd12;
							end
							mret_insn_i: begin
								// Trace: design.sv:7565:18
								csr_restore_mret_id_o = !debug_mode_q;
								// Trace: design.sv:7566:18
								ctrl_fsm_ns = 5'd10;
							end
							uret_insn_i: begin
								// Trace: design.sv:7569:18
								csr_restore_uret_id_o = !debug_mode_q;
								// Trace: design.sv:7570:18
								ctrl_fsm_ns = 5'd10;
							end
							dret_insn_i: begin
								// Trace: design.sv:7573:19
								csr_restore_dret_id_o = 1'b1;
								// Trace: design.sv:7574:19
								ctrl_fsm_ns = 5'd10;
							end
							csr_status_i: begin
								// Trace: design.sv:7579:17
								if (hwlp_end0_eq_pc && hwlp_counter0_gt_1) begin
									// Trace: design.sv:7580:21
									pc_mux_o = cv32e40p_pkg_PC_HWLOOP;
									// Trace: design.sv:7581:21
									pc_set_o = 1'b1;
									// Trace: design.sv:7582:21
									hwlp_dec_cnt_o[0] = 1'b1;
								end
								if (hwlp_end1_eq_pc && hwlp_counter1_gt_1) begin
									// Trace: design.sv:7585:21
									pc_mux_o = cv32e40p_pkg_PC_HWLOOP;
									// Trace: design.sv:7586:21
									pc_set_o = 1'b1;
									// Trace: design.sv:7587:21
									hwlp_dec_cnt_o[1] = 1'b1;
								end
							end
							wfi_i:
								// Trace: design.sv:7592:19
								if (debug_req_pending) begin
									// Trace: design.sv:7593:23
									ctrl_fsm_ns = 5'd12;
									// Trace: design.sv:7594:23
									debug_force_wakeup_n = 1'b1;
								end
								else
									// Trace: design.sv:7596:21
									ctrl_fsm_ns = 5'd3;
							fencei_insn_i: begin
								// Trace: design.sv:7602:19
								pc_mux_o = cv32e40p_pkg_PC_FENCEI;
								// Trace: design.sv:7603:19
								pc_set_o = 1'b1;
							end
							default:
								;
						endcase
			end
			5'd10: begin
				// Trace: design.sv:7614:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:7615:9
				ctrl_fsm_ns = 5'd5;
				// Trace: design.sv:7616:9
				(* full_case, parallel_case *)
				case (1'b1)
					mret_dec_i: begin
						// Trace: design.sv:7619:15
						pc_mux_o = (debug_mode_q ? cv32e40p_pkg_PC_EXCEPTION : cv32e40p_pkg_PC_MRET);
						// Trace: design.sv:7620:15
						pc_set_o = 1'b1;
						// Trace: design.sv:7621:15
						exc_pc_mux_o = cv32e40p_pkg_EXC_PC_DBE;
					end
					uret_dec_i: begin
						// Trace: design.sv:7625:15
						pc_mux_o = (debug_mode_q ? cv32e40p_pkg_PC_EXCEPTION : cv32e40p_pkg_PC_URET);
						// Trace: design.sv:7626:15
						pc_set_o = 1'b1;
						// Trace: design.sv:7627:15
						exc_pc_mux_o = cv32e40p_pkg_EXC_PC_DBE;
					end
					dret_dec_i: begin
						// Trace: design.sv:7632:15
						pc_mux_o = cv32e40p_pkg_PC_DRET;
						// Trace: design.sv:7633:15
						pc_set_o = 1'b1;
						// Trace: design.sv:7634:15
						debug_mode_n = 1'b0;
					end
					default:
						;
				endcase
				if (debug_single_step_i && ~debug_mode_q)
					// Trace: design.sv:7640:11
					ctrl_fsm_ns = 5'd12;
			end
			5'd14: begin
				// Trace: design.sv:7648:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:7649:9
				halt_if_o = 1'b1;
				// Trace: design.sv:7651:9
				if (branch_taken_ex_i) begin
					// Trace: design.sv:7653:11
					pc_mux_o = cv32e40p_pkg_PC_BRANCH;
					// Trace: design.sv:7654:11
					pc_set_o = 1'b1;
				end
				// Trace: design.sv:7657:9
				ctrl_fsm_ns = 5'd13;
			end
			5'd11: begin
				// Trace: design.sv:7671:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:7672:9
				pc_set_o = 1'b1;
				// Trace: design.sv:7673:9
				pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
				// Trace: design.sv:7674:9
				exc_pc_mux_o = cv32e40p_pkg_EXC_PC_DBD;
				// Trace: design.sv:7677:9
				if (~debug_mode_q) begin
					// Trace: design.sv:7678:13
					csr_save_cause_o = 1'b1;
					// Trace: design.sv:7679:13
					csr_save_id_o = 1'b1;
					// Trace: design.sv:7680:13
					debug_csr_save_o = 1'b1;
					// Trace: design.sv:7681:13
					if (trigger_match_i)
						// Trace: design.sv:7682:17
						debug_cause_o = cv32e40p_pkg_DBG_CAUSE_TRIGGER;
					else if (ebrk_force_debug_mode & ebrk_insn_i)
						// Trace: design.sv:7684:17
						debug_cause_o = cv32e40p_pkg_DBG_CAUSE_EBREAK;
					else if (debug_req_entry_q)
						// Trace: design.sv:7686:17
						debug_cause_o = cv32e40p_pkg_DBG_CAUSE_HALTREQ;
				end
				// Trace: design.sv:7689:9
				debug_req_entry_n = 1'b0;
				// Trace: design.sv:7690:9
				ctrl_fsm_ns = 5'd5;
				// Trace: design.sv:7691:9
				debug_mode_n = 1'b1;
			end
			5'd12: begin
				// Trace: design.sv:7698:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:7699:9
				pc_set_o = 1'b1;
				// Trace: design.sv:7700:9
				pc_mux_o = cv32e40p_pkg_PC_EXCEPTION;
				// Trace: design.sv:7701:9
				exc_pc_mux_o = cv32e40p_pkg_EXC_PC_DBD;
				// Trace: design.sv:7702:9
				csr_save_cause_o = 1'b1;
				// Trace: design.sv:7703:9
				debug_csr_save_o = 1'b1;
				// Trace: design.sv:7704:9
				if (debug_force_wakeup_q)
					// Trace: design.sv:7705:13
					debug_cause_o = cv32e40p_pkg_DBG_CAUSE_HALTREQ;
				else if (debug_single_step_i)
					// Trace: design.sv:7707:13
					debug_cause_o = cv32e40p_pkg_DBG_CAUSE_STEP;
				// Trace: design.sv:7708:9
				csr_save_if_o = 1'b1;
				// Trace: design.sv:7709:9
				ctrl_fsm_ns = 5'd5;
				// Trace: design.sv:7710:9
				debug_mode_n = 1'b1;
				// Trace: design.sv:7711:9
				debug_force_wakeup_n = 1'b0;
			end
			5'd13: begin
				// Trace: design.sv:7717:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:7719:9
				halt_if_o = 1'b1;
				// Trace: design.sv:7720:9
				halt_id_o = 1'b1;
				// Trace: design.sv:7722:9
				perf_pipeline_stall_o = data_load_event_i;
				// Trace: design.sv:7724:9
				if (data_err_i) begin
					// Trace: design.sv:7727:13
					csr_save_ex_o = 1'b1;
					// Trace: design.sv:7728:13
					csr_save_cause_o = 1'b1;
					// Trace: design.sv:7729:13
					data_err_ack_o = 1'b1;
					// Trace: design.sv:7731:13
					csr_cause_o = {1'b0, (data_we_ex_i ? cv32e40p_pkg_EXC_CAUSE_STORE_FAULT : cv32e40p_pkg_EXC_CAUSE_LOAD_FAULT)};
					// Trace: design.sv:7732:13
					ctrl_fsm_ns = 5'd9;
				end
				else
					// Trace: design.sv:7735:11
					if ((((debug_mode_q | trigger_match_i) | (ebrk_force_debug_mode & ebrk_insn_i)) | data_load_event_i) | debug_req_entry_q)
						// Trace: design.sv:7741:15
						ctrl_fsm_ns = 5'd11;
					else
						// Trace: design.sv:7745:15
						ctrl_fsm_ns = 5'd12;
			end
			default: begin
				// Trace: design.sv:7752:9
				is_decoding_o = 1'b0;
				// Trace: design.sv:7753:9
				instr_req_o = 1'b0;
				// Trace: design.sv:7754:9
				ctrl_fsm_ns = 5'd0;
			end
		endcase
	end
	// Trace: design.sv:7761:1
	generate
		if (PULP_XPULP) begin : gen_hwlp
			// Trace: design.sv:7774:5
			assign hwlp_jump_o = (hwlp_end_4_id_d && !hwlp_end_4_id_q ? 1'b1 : 1'b0);
			// Trace: design.sv:7776:5
			always @(posedge clk or negedge rst_n)
				// Trace: design.sv:7777:7
				if (!rst_n)
					// Trace: design.sv:7778:9
					hwlp_end_4_id_q <= 1'b0;
				else
					// Trace: design.sv:7780:9
					hwlp_end_4_id_q <= hwlp_end_4_id_d;
			// Trace: design.sv:7784:5
			assign hwlp_end0_eq_pc = hwlp_end_addr_i[0+:32] == pc_id_i;
			// Trace: design.sv:7785:5
			assign hwlp_end1_eq_pc = hwlp_end_addr_i[32+:32] == pc_id_i;
			// Trace: design.sv:7786:5
			assign hwlp_counter0_gt_1 = hwlp_counter_i[0+:32] > 1;
			// Trace: design.sv:7787:5
			assign hwlp_counter1_gt_1 = hwlp_counter_i[32+:32] > 1;
			// Trace: design.sv:7788:5
			assign hwlp_end0_eq_pc_plus4 = hwlp_end_addr_i[0+:32] == (pc_id_i + 4);
			// Trace: design.sv:7789:5
			assign hwlp_end1_eq_pc_plus4 = hwlp_end_addr_i[32+:32] == (pc_id_i + 4);
			// Trace: design.sv:7790:5
			assign hwlp_start0_leq_pc = hwlp_start_addr_i[0+:32] <= pc_id_i;
			// Trace: design.sv:7791:5
			assign hwlp_start1_leq_pc = hwlp_start_addr_i[32+:32] <= pc_id_i;
			// Trace: design.sv:7792:5
			assign hwlp_end0_geq_pc = hwlp_end_addr_i[0+:32] >= pc_id_i;
			// Trace: design.sv:7793:5
			assign hwlp_end1_geq_pc = hwlp_end_addr_i[32+:32] >= pc_id_i;
			// Trace: design.sv:7794:5
			assign is_hwlp_body = ((hwlp_start0_leq_pc && hwlp_end0_geq_pc) && hwlp_counter0_gt_1) || ((hwlp_start1_leq_pc && hwlp_end1_geq_pc) && hwlp_counter1_gt_1);
		end
		else begin : gen_no_hwlp
			// Trace: design.sv:7798:5
			assign hwlp_jump_o = 1'b0;
			// Trace: design.sv:7799:5
			wire [1:1] sv2v_tmp_6074E;
			assign sv2v_tmp_6074E = 1'b0;
			always @(*) hwlp_end_4_id_q = sv2v_tmp_6074E;
			// Trace: design.sv:7800:5
			assign hwlp_end0_eq_pc = 1'b0;
			// Trace: design.sv:7801:5
			assign hwlp_end1_eq_pc = 1'b0;
			// Trace: design.sv:7802:5
			assign hwlp_counter0_gt_1 = 1'b0;
			// Trace: design.sv:7803:5
			assign hwlp_counter1_gt_1 = 1'b0;
			// Trace: design.sv:7804:5
			assign hwlp_end0_eq_pc_plus4 = 1'b0;
			// Trace: design.sv:7805:5
			assign hwlp_end1_eq_pc_plus4 = 1'b0;
			// Trace: design.sv:7806:5
			assign hwlp_start0_leq_pc = 1'b0;
			// Trace: design.sv:7807:5
			assign hwlp_start1_leq_pc = 1'b0;
			// Trace: design.sv:7808:5
			assign hwlp_end0_geq_pc = 1'b0;
			// Trace: design.sv:7809:5
			assign hwlp_end1_geq_pc = 1'b0;
			// Trace: design.sv:7810:5
			assign is_hwlp_body = 1'b0;
		end
	endgenerate
	// Trace: design.sv:7824:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:7826:5
		load_stall_o = 1'b0;
		// Trace: design.sv:7827:5
		deassert_we_o = 1'b0;
		// Trace: design.sv:7830:5
		if (~is_decoding_o)
			// Trace: design.sv:7831:7
			deassert_we_o = 1'b1;
		if (illegal_insn_i)
			// Trace: design.sv:7835:7
			deassert_we_o = 1'b1;
		if ((((data_req_ex_i == 1'b1) && (regfile_we_ex_i == 1'b1)) || ((wb_ready_i == 1'b0) && (regfile_we_wb_i == 1'b1))) && ((((reg_d_ex_is_reg_a_i == 1'b1) || (reg_d_ex_is_reg_b_i == 1'b1)) || (reg_d_ex_is_reg_c_i == 1'b1)) || ((is_decoding_o && (regfile_we_id_i && !data_misaligned_i)) && (regfile_waddr_ex_i == regfile_alu_waddr_id_i)))) begin
			// Trace: design.sv:7846:7
			deassert_we_o = 1'b1;
			// Trace: design.sv:7847:7
			load_stall_o = 1'b1;
		end
		if ((ctrl_transfer_insn_in_dec_i == cv32e40p_pkg_BRANCH_JALR) && ((((regfile_we_wb_i == 1'b1) && (reg_d_wb_is_reg_a_i == 1'b1)) || ((regfile_we_ex_i == 1'b1) && (reg_d_ex_is_reg_a_i == 1'b1))) || ((regfile_alu_we_fw_i == 1'b1) && (reg_d_alu_is_reg_a_i == 1'b1)))) begin
			// Trace: design.sv:7859:7
			jr_stall_o = 1'b1;
			// Trace: design.sv:7860:7
			deassert_we_o = 1'b1;
		end
		else
			// Trace: design.sv:7864:7
			jr_stall_o = 1'b0;
	end
	// Trace: design.sv:7870:3
	assign misaligned_stall_o = data_misaligned_i;
	// Trace: design.sv:7873:3
	assign apu_stall_o = apu_read_dep_i | (apu_write_dep_i & ~apu_en_i);
	// Trace: design.sv:7876:3
	localparam cv32e40p_pkg_SEL_FW_EX = 2'b01;
	localparam cv32e40p_pkg_SEL_FW_WB = 2'b10;
	localparam cv32e40p_pkg_SEL_REGFILE = 2'b00;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:7879:5
		operand_a_fw_mux_sel_o = cv32e40p_pkg_SEL_REGFILE;
		// Trace: design.sv:7880:5
		operand_b_fw_mux_sel_o = cv32e40p_pkg_SEL_REGFILE;
		// Trace: design.sv:7881:5
		operand_c_fw_mux_sel_o = cv32e40p_pkg_SEL_REGFILE;
		// Trace: design.sv:7884:5
		if (regfile_we_wb_i == 1'b1) begin
			// Trace: design.sv:7886:7
			if (reg_d_wb_is_reg_a_i == 1'b1)
				// Trace: design.sv:7887:9
				operand_a_fw_mux_sel_o = cv32e40p_pkg_SEL_FW_WB;
			if (reg_d_wb_is_reg_b_i == 1'b1)
				// Trace: design.sv:7889:9
				operand_b_fw_mux_sel_o = cv32e40p_pkg_SEL_FW_WB;
			if (reg_d_wb_is_reg_c_i == 1'b1)
				// Trace: design.sv:7891:9
				operand_c_fw_mux_sel_o = cv32e40p_pkg_SEL_FW_WB;
		end
		if (regfile_alu_we_fw_i == 1'b1) begin
			// Trace: design.sv:7897:6
			if (reg_d_alu_is_reg_a_i == 1'b1)
				// Trace: design.sv:7898:8
				operand_a_fw_mux_sel_o = cv32e40p_pkg_SEL_FW_EX;
			if (reg_d_alu_is_reg_b_i == 1'b1)
				// Trace: design.sv:7900:8
				operand_b_fw_mux_sel_o = cv32e40p_pkg_SEL_FW_EX;
			if (reg_d_alu_is_reg_c_i == 1'b1)
				// Trace: design.sv:7902:8
				operand_c_fw_mux_sel_o = cv32e40p_pkg_SEL_FW_EX;
		end
		if (data_misaligned_i) begin
			// Trace: design.sv:7908:7
			operand_a_fw_mux_sel_o = cv32e40p_pkg_SEL_FW_EX;
			// Trace: design.sv:7909:7
			operand_b_fw_mux_sel_o = cv32e40p_pkg_SEL_REGFILE;
		end
		else if (mult_multicycle_i)
			// Trace: design.sv:7911:7
			operand_c_fw_mux_sel_o = cv32e40p_pkg_SEL_FW_EX;
	end
	// Trace: design.sv:7916:3
	always @(posedge clk or negedge rst_n) begin : UPDATE_REGS
		// Trace: design.sv:7918:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:7920:7
			ctrl_fsm_cs <= 5'd0;
			// Trace: design.sv:7921:7
			jump_done_q <= 1'b0;
			// Trace: design.sv:7922:7
			data_err_q <= 1'b0;
			// Trace: design.sv:7924:7
			debug_mode_q <= 1'b0;
			// Trace: design.sv:7925:7
			illegal_insn_q <= 1'b0;
			// Trace: design.sv:7927:7
			debug_req_entry_q <= 1'b0;
			// Trace: design.sv:7928:7
			debug_force_wakeup_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:7932:7
			ctrl_fsm_cs <= ctrl_fsm_ns;
			// Trace: design.sv:7935:7
			jump_done_q <= jump_done & ~id_ready_i;
			// Trace: design.sv:7937:7
			data_err_q <= data_err_i;
			// Trace: design.sv:7939:7
			debug_mode_q <= debug_mode_n;
			// Trace: design.sv:7941:7
			illegal_insn_q <= illegal_insn_n;
			// Trace: design.sv:7943:7
			debug_req_entry_q <= debug_req_entry_n;
			// Trace: design.sv:7944:7
			debug_force_wakeup_q <= debug_force_wakeup_n;
		end
	end
	// Trace: design.sv:7949:3
	assign wake_from_sleep_o = (irq_wu_ctrl_i || debug_req_pending) || debug_mode_q;
	// Trace: design.sv:7952:3
	assign debug_mode_o = debug_mode_q;
	// Trace: design.sv:7953:3
	assign debug_req_pending = debug_req_i || debug_req_q;
	// Trace: design.sv:7956:3
	assign debug_p_elw_no_sleep_o = ((debug_mode_q || debug_req_q) || debug_single_step_i) || trigger_match_i;
	// Trace: design.sv:7963:3
	assign debug_wfi_no_sleep_o = (((debug_mode_q || debug_req_pending) || debug_single_step_i) || trigger_match_i) || PULP_CLUSTER;
	// Trace: design.sv:7966:3
	assign wfi_active = wfi_i & ~debug_wfi_no_sleep_o;
	// Trace: design.sv:7969:3
	always @(posedge clk_ungated_i or negedge rst_n)
		if (!rst_n)
			// Trace: design.sv:7971:7
			debug_req_q <= 1'b0;
		else if (debug_req_i)
			// Trace: design.sv:7974:9
			debug_req_q <= 1'b1;
		else if (debug_mode_q)
			// Trace: design.sv:7976:9
			debug_req_q <= 1'b0;
	// Trace: design.sv:7979:3
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:7981:5
		if (rst_n == 1'b0)
			// Trace: design.sv:7983:7
			debug_fsm_cs <= 3'b001;
		else
			// Trace: design.sv:7987:7
			debug_fsm_cs <= debug_fsm_ns;
	// Trace: design.sv:7991:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:7993:5
		debug_fsm_ns = debug_fsm_cs;
		// Trace: design.sv:7995:5
		case (debug_fsm_cs)
			3'b001:
				// Trace: design.sv:7998:9
				if (debug_mode_n || (ctrl_fsm_ns == 5'd4)) begin
					begin
						// Trace: design.sv:7999:11
						if (debug_mode_n)
							// Trace: design.sv:8000:13
							debug_fsm_ns = 3'b100;
						else
							// Trace: design.sv:8002:13
							debug_fsm_ns = 3'b010;
					end
				end
			3'b010:
				// Trace: design.sv:8009:9
				if (debug_mode_n)
					// Trace: design.sv:8010:11
					debug_fsm_ns = 3'b100;
			3'b100:
				// Trace: design.sv:8016:9
				if (!debug_mode_n)
					// Trace: design.sv:8017:11
					debug_fsm_ns = 3'b010;
			default:
				// Trace: design.sv:8022:9
				debug_fsm_ns = 3'b001;
		endcase
	end
	// Trace: design.sv:8027:3
	localparam cv32e40p_pkg_HAVERESET_INDEX = 0;
	assign debug_havereset_o = debug_fsm_cs[cv32e40p_pkg_HAVERESET_INDEX];
	// Trace: design.sv:8028:3
	localparam cv32e40p_pkg_RUNNING_INDEX = 1;
	assign debug_running_o = debug_fsm_cs[cv32e40p_pkg_RUNNING_INDEX];
	// Trace: design.sv:8029:3
	localparam cv32e40p_pkg_HALTED_INDEX = 2;
	assign debug_halted_o = debug_fsm_cs[cv32e40p_pkg_HALTED_INDEX];
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_cs_registers (
	clk,
	rst_n,
	hart_id_i,
	mtvec_o,
	utvec_o,
	mtvec_mode_o,
	utvec_mode_o,
	mtvec_addr_i,
	csr_mtvec_init_i,
	csr_addr_i,
	csr_wdata_i,
	csr_op_i,
	csr_rdata_o,
	frm_o,
	fflags_i,
	fflags_we_i,
	mie_bypass_o,
	mip_i,
	m_irq_enable_o,
	u_irq_enable_o,
	csr_irq_sec_i,
	sec_lvl_o,
	mepc_o,
	uepc_o,
	mcounteren_o,
	debug_mode_i,
	debug_cause_i,
	debug_csr_save_i,
	depc_o,
	debug_single_step_o,
	debug_ebreakm_o,
	debug_ebreaku_o,
	trigger_match_o,
	pmp_addr_o,
	pmp_cfg_o,
	priv_lvl_o,
	pc_if_i,
	pc_id_i,
	pc_ex_i,
	csr_save_if_i,
	csr_save_id_i,
	csr_save_ex_i,
	csr_restore_mret_i,
	csr_restore_uret_i,
	csr_restore_dret_i,
	csr_cause_i,
	csr_save_cause_i,
	hwlp_start_i,
	hwlp_end_i,
	hwlp_cnt_i,
	hwlp_data_o,
	hwlp_regid_o,
	hwlp_we_o,
	mhpmevent_minstret_i,
	mhpmevent_load_i,
	mhpmevent_store_i,
	mhpmevent_jump_i,
	mhpmevent_branch_i,
	mhpmevent_branch_taken_i,
	mhpmevent_compressed_i,
	mhpmevent_jr_stall_i,
	mhpmevent_imiss_i,
	mhpmevent_ld_stall_i,
	mhpmevent_pipe_stall_i,
	apu_typeconflict_i,
	apu_contention_i,
	apu_dep_i,
	apu_wb_i
);
	reg _sv2v_0;
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:8138:15
	parameter N_HWLP = 2;
	// Trace: design.sv:8139:15
	parameter N_HWLP_BITS = $clog2(N_HWLP);
	// Trace: design.sv:8140:15
	parameter APU = 0;
	// Trace: design.sv:8141:15
	parameter A_EXTENSION = 0;
	// Trace: design.sv:8142:15
	parameter FPU = 0;
	// Trace: design.sv:8143:15
	parameter PULP_SECURE = 0;
	// Trace: design.sv:8144:15
	parameter USE_PMP = 0;
	// Trace: design.sv:8145:15
	parameter N_PMP_ENTRIES = 16;
	// Trace: design.sv:8146:15
	parameter NUM_MHPMCOUNTERS = 1;
	// Trace: design.sv:8147:15
	parameter PULP_XPULP = 0;
	// Trace: design.sv:8148:15
	parameter PULP_CLUSTER = 0;
	// Trace: design.sv:8149:15
	parameter DEBUG_TRIGGER_EN = 1;
	// Trace: design.sv:8152:5
	input wire clk;
	// Trace: design.sv:8153:5
	input wire rst_n;
	// Trace: design.sv:8156:5
	input wire [31:0] hart_id_i;
	// Trace: design.sv:8157:5
	output wire [23:0] mtvec_o;
	// Trace: design.sv:8158:5
	output wire [23:0] utvec_o;
	// Trace: design.sv:8159:5
	output wire [1:0] mtvec_mode_o;
	// Trace: design.sv:8160:5
	output wire [1:0] utvec_mode_o;
	// Trace: design.sv:8163:5
	input wire [31:0] mtvec_addr_i;
	// Trace: design.sv:8164:5
	input wire csr_mtvec_init_i;
	// Trace: design.sv:8167:5
	// removed localparam type cv32e40p_pkg_csr_num_e
	input wire [11:0] csr_addr_i;
	// Trace: design.sv:8168:5
	input wire [31:0] csr_wdata_i;
	// Trace: design.sv:8169:5
	localparam cv32e40p_pkg_CSR_OP_WIDTH = 2;
	// removed localparam type cv32e40p_pkg_csr_opcode_e
	input wire [1:0] csr_op_i;
	// Trace: design.sv:8170:5
	output wire [31:0] csr_rdata_o;
	// Trace: design.sv:8172:5
	output wire [2:0] frm_o;
	// Trace: design.sv:8173:5
	localparam cv32e40p_pkg_C_FFLAG = 5;
	input wire [4:0] fflags_i;
	// Trace: design.sv:8174:5
	input wire fflags_we_i;
	// Trace: design.sv:8177:5
	output wire [31:0] mie_bypass_o;
	// Trace: design.sv:8178:5
	input wire [31:0] mip_i;
	// Trace: design.sv:8179:5
	output wire m_irq_enable_o;
	// Trace: design.sv:8180:5
	output wire u_irq_enable_o;
	// Trace: design.sv:8183:5
	input wire csr_irq_sec_i;
	// Trace: design.sv:8184:5
	output wire sec_lvl_o;
	// Trace: design.sv:8185:5
	output wire [31:0] mepc_o;
	// Trace: design.sv:8186:5
	output wire [31:0] uepc_o;
	// Trace: design.sv:8188:5
	output wire [31:0] mcounteren_o;
	// Trace: design.sv:8191:5
	input wire debug_mode_i;
	// Trace: design.sv:8192:5
	input wire [2:0] debug_cause_i;
	// Trace: design.sv:8193:5
	input wire debug_csr_save_i;
	// Trace: design.sv:8194:5
	output wire [31:0] depc_o;
	// Trace: design.sv:8195:5
	output wire debug_single_step_o;
	// Trace: design.sv:8196:5
	output wire debug_ebreakm_o;
	// Trace: design.sv:8197:5
	output wire debug_ebreaku_o;
	// Trace: design.sv:8198:5
	output wire trigger_match_o;
	// Trace: design.sv:8201:5
	output wire [(N_PMP_ENTRIES * 32) - 1:0] pmp_addr_o;
	// Trace: design.sv:8202:5
	output wire [(N_PMP_ENTRIES * 8) - 1:0] pmp_cfg_o;
	// Trace: design.sv:8204:5
	// removed localparam type cv32e40p_pkg_PrivLvl_t
	output wire [1:0] priv_lvl_o;
	// Trace: design.sv:8206:5
	input wire [31:0] pc_if_i;
	// Trace: design.sv:8207:5
	input wire [31:0] pc_id_i;
	// Trace: design.sv:8208:5
	input wire [31:0] pc_ex_i;
	// Trace: design.sv:8210:5
	input wire csr_save_if_i;
	// Trace: design.sv:8211:5
	input wire csr_save_id_i;
	// Trace: design.sv:8212:5
	input wire csr_save_ex_i;
	// Trace: design.sv:8214:5
	input wire csr_restore_mret_i;
	// Trace: design.sv:8215:5
	input wire csr_restore_uret_i;
	// Trace: design.sv:8217:5
	input wire csr_restore_dret_i;
	// Trace: design.sv:8219:5
	input wire [5:0] csr_cause_i;
	// Trace: design.sv:8221:5
	input wire csr_save_cause_i;
	// Trace: design.sv:8223:5
	input wire [(N_HWLP * 32) - 1:0] hwlp_start_i;
	// Trace: design.sv:8224:5
	input wire [(N_HWLP * 32) - 1:0] hwlp_end_i;
	// Trace: design.sv:8225:5
	input wire [(N_HWLP * 32) - 1:0] hwlp_cnt_i;
	// Trace: design.sv:8227:5
	output wire [31:0] hwlp_data_o;
	// Trace: design.sv:8228:5
	output reg [N_HWLP_BITS - 1:0] hwlp_regid_o;
	// Trace: design.sv:8229:5
	output reg [2:0] hwlp_we_o;
	// Trace: design.sv:8232:5
	input wire mhpmevent_minstret_i;
	// Trace: design.sv:8233:5
	input wire mhpmevent_load_i;
	// Trace: design.sv:8234:5
	input wire mhpmevent_store_i;
	// Trace: design.sv:8235:5
	input wire mhpmevent_jump_i;
	// Trace: design.sv:8236:5
	input wire mhpmevent_branch_i;
	// Trace: design.sv:8237:5
	input wire mhpmevent_branch_taken_i;
	// Trace: design.sv:8238:5
	input wire mhpmevent_compressed_i;
	// Trace: design.sv:8239:5
	input wire mhpmevent_jr_stall_i;
	// Trace: design.sv:8240:5
	input wire mhpmevent_imiss_i;
	// Trace: design.sv:8241:5
	input wire mhpmevent_ld_stall_i;
	// Trace: design.sv:8242:5
	input wire mhpmevent_pipe_stall_i;
	// Trace: design.sv:8243:5
	input wire apu_typeconflict_i;
	// Trace: design.sv:8244:5
	input wire apu_contention_i;
	// Trace: design.sv:8245:5
	input wire apu_dep_i;
	// Trace: design.sv:8246:5
	input wire apu_wb_i;
	// Trace: design.sv:8249:3
	localparam NUM_HPM_EVENTS = 16;
	// Trace: design.sv:8251:3
	localparam MTVEC_MODE = 2'b01;
	// Trace: design.sv:8253:3
	localparam MAX_N_PMP_ENTRIES = 16;
	// Trace: design.sv:8254:3
	localparam MAX_N_PMP_CFG = 4;
	// Trace: design.sv:8255:3
	localparam N_PMP_CFG = ((N_PMP_ENTRIES % 4) == 0 ? N_PMP_ENTRIES / 4 : (N_PMP_ENTRIES / 4) + 1);
	// Trace: design.sv:8257:3
	localparam MSTATUS_UIE_BIT = 0;
	// Trace: design.sv:8258:3
	localparam MSTATUS_SIE_BIT = 1;
	// Trace: design.sv:8259:3
	localparam MSTATUS_MIE_BIT = 3;
	// Trace: design.sv:8260:3
	localparam MSTATUS_UPIE_BIT = 4;
	// Trace: design.sv:8261:3
	localparam MSTATUS_SPIE_BIT = 5;
	// Trace: design.sv:8262:3
	localparam MSTATUS_MPIE_BIT = 7;
	// Trace: design.sv:8263:3
	localparam MSTATUS_SPP_BIT = 8;
	// Trace: design.sv:8264:3
	localparam MSTATUS_MPP_BIT_HIGH = 12;
	// Trace: design.sv:8265:3
	localparam MSTATUS_MPP_BIT_LOW = 11;
	// Trace: design.sv:8266:3
	localparam MSTATUS_MPRV_BIT = 17;
	// Trace: design.sv:8269:3
	localparam [1:0] MXL = 2'd1;
	// Trace: design.sv:8270:3
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	localparam [31:0] MISA_VALUE = (((((((((((A_EXTENSION << 0) | 4) | 0) | 0) | (FPU << 5)) | 256) | 4096) | 0) | 0) | (PULP_SECURE << 20)) | (sv2v_cast_32(PULP_XPULP || PULP_CLUSTER) << 23)) | (sv2v_cast_32(MXL) << 30);
	// Trace: design.sv:8283:3
	localparam MHPMCOUNTER_WIDTH = 64;
	// Trace: design.sv:8288:3
	localparam PULP_PERF_COUNTERS = 0;
	// Trace: design.sv:8290:3
	// removed localparam type Status_t
	// Trace: design.sv:8305:3
	// removed localparam type Dcsr_t
	// Trace: design.sv:8323:3
	// removed localparam type Pmp_t
	// Trace: design.sv:8330:3
	reg [31:0] csr_wdata_int;
	// Trace: design.sv:8331:3
	reg [31:0] csr_rdata_int;
	// Trace: design.sv:8332:3
	reg csr_we_int;
	// Trace: design.sv:8333:3
	localparam cv32e40p_pkg_C_RM = 3;
	reg [2:0] frm_q;
	reg [2:0] frm_n;
	// Trace: design.sv:8334:3
	reg [4:0] fflags_q;
	reg [4:0] fflags_n;
	// Trace: design.sv:8337:3
	reg [31:0] mepc_q;
	reg [31:0] mepc_n;
	// Trace: design.sv:8338:3
	reg [31:0] uepc_q;
	reg [31:0] uepc_n;
	// Trace: design.sv:8340:3
	wire [31:0] tmatch_control_rdata;
	// Trace: design.sv:8341:3
	wire [31:0] tmatch_value_rdata;
	// Trace: design.sv:8342:3
	wire [15:0] tinfo_types;
	// Trace: design.sv:8344:3
	reg [31:0] dcsr_q;
	reg [31:0] dcsr_n;
	// Trace: design.sv:8345:3
	reg [31:0] depc_q;
	reg [31:0] depc_n;
	// Trace: design.sv:8346:3
	reg [31:0] dscratch0_q;
	reg [31:0] dscratch0_n;
	// Trace: design.sv:8347:3
	reg [31:0] dscratch1_q;
	reg [31:0] dscratch1_n;
	// Trace: design.sv:8348:3
	reg [31:0] mscratch_q;
	reg [31:0] mscratch_n;
	// Trace: design.sv:8350:3
	reg [31:0] exception_pc;
	// Trace: design.sv:8351:3
	reg [6:0] mstatus_q;
	reg [6:0] mstatus_n;
	// Trace: design.sv:8352:3
	reg [5:0] mcause_q;
	reg [5:0] mcause_n;
	// Trace: design.sv:8353:3
	reg [5:0] ucause_q;
	reg [5:0] ucause_n;
	// Trace: design.sv:8355:3
	reg [23:0] mtvec_n;
	reg [23:0] mtvec_q;
	// Trace: design.sv:8356:3
	reg [23:0] utvec_n;
	reg [23:0] utvec_q;
	// Trace: design.sv:8357:3
	reg [1:0] mtvec_mode_n;
	reg [1:0] mtvec_mode_q;
	// Trace: design.sv:8358:3
	reg [1:0] utvec_mode_n;
	reg [1:0] utvec_mode_q;
	// Trace: design.sv:8360:3
	wire [31:0] mip;
	// Trace: design.sv:8361:3
	reg [31:0] mie_q;
	reg [31:0] mie_n;
	// Trace: design.sv:8363:3
	reg [31:0] csr_mie_wdata;
	// Trace: design.sv:8364:3
	reg csr_mie_we;
	// Trace: design.sv:8366:3
	wire is_irq;
	// Trace: design.sv:8367:3
	reg [1:0] priv_lvl_n;
	reg [1:0] priv_lvl_q;
	// Trace: design.sv:8368:3
	reg [767:0] pmp_reg_q;
	reg [767:0] pmp_reg_n;
	// Trace: design.sv:8370:3
	reg [15:0] pmpaddr_we;
	// Trace: design.sv:8371:3
	reg [15:0] pmpcfg_we;
	// Trace: design.sv:8374:3
	reg [2047:0] mhpmcounter_q;
	// Trace: design.sv:8375:3
	reg [1023:0] mhpmevent_q;
	reg [1023:0] mhpmevent_n;
	// Trace: design.sv:8376:3
	reg [31:0] mcounteren_q;
	reg [31:0] mcounteren_n;
	// Trace: design.sv:8377:3
	reg [31:0] mcountinhibit_q;
	reg [31:0] mcountinhibit_n;
	// Trace: design.sv:8378:3
	wire [15:0] hpm_events;
	// Trace: design.sv:8379:3
	wire [2047:0] mhpmcounter_increment;
	// Trace: design.sv:8380:3
	wire [31:0] mhpmcounter_write_lower;
	// Trace: design.sv:8381:3
	wire [31:0] mhpmcounter_write_upper;
	// Trace: design.sv:8382:3
	wire [31:0] mhpmcounter_write_increment;
	// Trace: design.sv:8384:3
	assign is_irq = csr_cause_i[5];
	// Trace: design.sv:8387:3
	assign mip = mip_i;
	// Trace: design.sv:8393:3
	function automatic [1:0] sv2v_cast_EB06E;
		input reg [1:0] inp;
		sv2v_cast_EB06E = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:8394:5
		csr_mie_wdata = csr_wdata_i;
		// Trace: design.sv:8395:5
		csr_mie_we = 1'b1;
		// Trace: design.sv:8397:5
		case (csr_op_i)
			sv2v_cast_EB06E(2'b01):
				// Trace: design.sv:8398:21
				csr_mie_wdata = csr_wdata_i;
			sv2v_cast_EB06E(2'b10):
				// Trace: design.sv:8399:21
				csr_mie_wdata = csr_wdata_i | mie_q;
			sv2v_cast_EB06E(2'b11):
				// Trace: design.sv:8400:21
				csr_mie_wdata = ~csr_wdata_i & mie_q;
			sv2v_cast_EB06E(2'b00): begin
				// Trace: design.sv:8402:9
				csr_mie_wdata = csr_wdata_i;
				// Trace: design.sv:8403:9
				csr_mie_we = 1'b0;
			end
		endcase
	end
	// Trace: design.sv:8408:3
	localparam cv32e40p_pkg_IRQ_MASK = 32'hffff0888;
	assign mie_bypass_o = ((csr_addr_i == 12'h304) && csr_mie_we ? csr_mie_wdata & cv32e40p_pkg_IRQ_MASK : mie_q);
	// Trace: design.sv:8422:3
	genvar _gv_j_3;
	// Trace: design.sv:8425:3
	localparam cv32e40p_pkg_MARCHID = 32'h00000004;
	localparam cv32e40p_pkg_MVENDORID_BANK = 25'h000000c;
	localparam cv32e40p_pkg_MVENDORID_OFFSET = 7'h02;
	generate
		if (PULP_SECURE == 1) begin : gen_pulp_secure_read_logic
			// Trace: design.sv:8427:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:8428:7
				case (csr_addr_i)
					12'h001:
						// Trace: design.sv:8430:21
						csr_rdata_int = (FPU == 1 ? {27'b000000000000000000000000000, fflags_q} : {32 {1'sb0}});
					12'h002:
						// Trace: design.sv:8431:21
						csr_rdata_int = (FPU == 1 ? {29'b00000000000000000000000000000, frm_q} : {32 {1'sb0}});
					12'h003:
						// Trace: design.sv:8432:21
						csr_rdata_int = (FPU == 1 ? {24'b000000000000000000000000, frm_q, fflags_q} : {32 {1'sb0}});
					12'h300:
						// Trace: design.sv:8436:9
						csr_rdata_int = {14'b00000000000000, mstatus_q[0], 4'b0000, mstatus_q[2-:2], 3'b000, mstatus_q[3], 2'h0, mstatus_q[4], mstatus_q[5], 2'h0, mstatus_q[6]};
					12'h301:
						// Trace: design.sv:8451:19
						csr_rdata_int = MISA_VALUE;
					12'h304:
						// Trace: design.sv:8455:11
						csr_rdata_int = mie_q;
					12'h305:
						// Trace: design.sv:8459:20
						csr_rdata_int = {mtvec_q, 6'h00, mtvec_mode_q};
					12'h340:
						// Trace: design.sv:8461:23
						csr_rdata_int = mscratch_q;
					12'h341:
						// Trace: design.sv:8463:19
						csr_rdata_int = mepc_q;
					12'h342:
						// Trace: design.sv:8465:21
						csr_rdata_int = {mcause_q[5], 26'b00000000000000000000000000, mcause_q[4:0]};
					12'h344:
						// Trace: design.sv:8468:11
						csr_rdata_int = mip;
					12'hf14:
						// Trace: design.sv:8472:22
						csr_rdata_int = hart_id_i;
					12'hf11:
						// Trace: design.sv:8475:24
						csr_rdata_int = {cv32e40p_pkg_MVENDORID_BANK, cv32e40p_pkg_MVENDORID_OFFSET};
					12'hf12:
						// Trace: design.sv:8478:22
						csr_rdata_int = cv32e40p_pkg_MARCHID;
					12'hf13, 12'h343:
						// Trace: design.sv:8481:32
						csr_rdata_int = 'b0;
					12'h306:
						// Trace: design.sv:8484:25
						csr_rdata_int = mcounteren_q;
					12'h7a0, 12'h7a3, 12'h7a8, 12'h7aa:
						// Trace: design.sv:8486:62
						csr_rdata_int = 'b0;
					12'h7a1:
						// Trace: design.sv:8487:21
						csr_rdata_int = tmatch_control_rdata;
					12'h7a2:
						// Trace: design.sv:8488:21
						csr_rdata_int = tmatch_value_rdata;
					12'h7a4:
						// Trace: design.sv:8489:20
						csr_rdata_int = tinfo_types;
					12'h7b0:
						// Trace: design.sv:8491:19
						csr_rdata_int = dcsr_q;
					12'h7b1:
						// Trace: design.sv:8492:18
						csr_rdata_int = depc_q;
					12'h7b2:
						// Trace: design.sv:8493:24
						csr_rdata_int = dscratch0_q;
					12'h7b3:
						// Trace: design.sv:8494:24
						csr_rdata_int = dscratch1_q;
					12'hb00, 12'hb02, 12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f, 12'hc00, 12'hc02, 12'hc03, 12'hc04, 12'hc05, 12'hc06, 12'hc07, 12'hc08, 12'hc09, 12'hc0a, 12'hc0b, 12'hc0c, 12'hc0d, 12'hc0e, 12'hc0f, 12'hc10, 12'hc11, 12'hc12, 12'hc13, 12'hc14, 12'hc15, 12'hc16, 12'hc17, 12'hc18, 12'hc19, 12'hc1a, 12'hc1b, 12'hc1c, 12'hc1d, 12'hc1e, 12'hc1f:
						// Trace: design.sv:8517:9
						csr_rdata_int = mhpmcounter_q[(csr_addr_i[4:0] * 64) + 31-:32];
					12'hb80, 12'hb82, 12'hb83, 12'hb84, 12'hb85, 12'hb86, 12'hb87, 12'hb88, 12'hb89, 12'hb8a, 12'hb8b, 12'hb8c, 12'hb8d, 12'hb8e, 12'hb8f, 12'hb90, 12'hb91, 12'hb92, 12'hb93, 12'hb94, 12'hb95, 12'hb96, 12'hb97, 12'hb98, 12'hb99, 12'hb9a, 12'hb9b, 12'hb9c, 12'hb9d, 12'hb9e, 12'hb9f, 12'hc80, 12'hc82, 12'hc83, 12'hc84, 12'hc85, 12'hc86, 12'hc87, 12'hc88, 12'hc89, 12'hc8a, 12'hc8b, 12'hc8c, 12'hc8d, 12'hc8e, 12'hc8f, 12'hc90, 12'hc91, 12'hc92, 12'hc93, 12'hc94, 12'hc95, 12'hc96, 12'hc97, 12'hc98, 12'hc99, 12'hc9a, 12'hc9b, 12'hc9c, 12'hc9d, 12'hc9e, 12'hc9f:
						// Trace: design.sv:8539:9
						csr_rdata_int = mhpmcounter_q[(csr_addr_i[4:0] * 64) + 63-:32];
					12'h320:
						// Trace: design.sv:8541:28
						csr_rdata_int = mcountinhibit_q;
					12'h323, 12'h324, 12'h325, 12'h326, 12'h327, 12'h328, 12'h329, 12'h32a, 12'h32b, 12'h32c, 12'h32d, 12'h32e, 12'h32f, 12'h330, 12'h331, 12'h332, 12'h333, 12'h334, 12'h335, 12'h336, 12'h337, 12'h338, 12'h339, 12'h33a, 12'h33b, 12'h33c, 12'h33d, 12'h33e, 12'h33f:
						// Trace: design.sv:8551:9
						csr_rdata_int = mhpmevent_q[csr_addr_i[4:0] * 32+:32];
					12'h800:
						// Trace: design.sv:8554:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_start_i[0+:32]);
					12'h801:
						// Trace: design.sv:8555:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_end_i[0+:32]);
					12'h802:
						// Trace: design.sv:8556:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_cnt_i[0+:32]);
					12'h804:
						// Trace: design.sv:8557:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_start_i[32+:32]);
					12'h805:
						// Trace: design.sv:8558:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_end_i[32+:32]);
					12'h806:
						// Trace: design.sv:8559:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_cnt_i[32+:32]);
					12'h3a0:
						// Trace: design.sv:8562:22
						csr_rdata_int = (USE_PMP ? pmp_reg_q[128+:32] : {32 {1'sb0}});
					12'h3a1:
						// Trace: design.sv:8563:22
						csr_rdata_int = (USE_PMP ? pmp_reg_q[160+:32] : {32 {1'sb0}});
					12'h3a2:
						// Trace: design.sv:8564:22
						csr_rdata_int = (USE_PMP ? pmp_reg_q[192+:32] : {32 {1'sb0}});
					12'h3a3:
						// Trace: design.sv:8565:22
						csr_rdata_int = (USE_PMP ? pmp_reg_q[224+:32] : {32 {1'sb0}});
					12'h3b0, 12'h3b1, 12'h3b2, 12'h3b3, 12'h3b4, 12'h3b5, 12'h3b6, 12'h3b7, 12'h3b8, 12'h3b9, 12'h3ba, 12'h3bb, 12'h3bc, 12'h3bd, 12'h3be, 12'h3bf:
						// Trace: design.sv:8571:9
						csr_rdata_int = (USE_PMP ? pmp_reg_q[256 + (csr_addr_i[3:0] * 32)+:32] : {32 {1'sb0}});
					12'h000:
						// Trace: design.sv:8575:22
						csr_rdata_int = {27'b000000000000000000000000000, mstatus_q[4], 3'h0, mstatus_q[6]};
					12'h005:
						// Trace: design.sv:8577:20
						csr_rdata_int = {utvec_q, 6'h00, utvec_mode_q};
					12'hcc0:
						// Trace: design.sv:8579:22
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hart_id_i);
					12'h041:
						// Trace: design.sv:8581:19
						csr_rdata_int = uepc_q;
					12'h042:
						// Trace: design.sv:8583:21
						csr_rdata_int = {ucause_q[5], 26'h0000000, ucause_q[4:0]};
					12'hcc1:
						// Trace: design.sv:8586:21
						csr_rdata_int = (!PULP_XPULP ? 'b0 : {30'h00000000, priv_lvl_q});
					default:
						// Trace: design.sv:8588:18
						csr_rdata_int = 1'sb0;
				endcase
			end
		end
		else begin : gen_no_pulp_secure_read_logic
			// Trace: design.sv:8593:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:8595:7
				case (csr_addr_i)
					12'h001:
						// Trace: design.sv:8597:21
						csr_rdata_int = (FPU == 1 ? {27'b000000000000000000000000000, fflags_q} : {32 {1'sb0}});
					12'h002:
						// Trace: design.sv:8598:18
						csr_rdata_int = (FPU == 1 ? {29'b00000000000000000000000000000, frm_q} : {32 {1'sb0}});
					12'h003:
						// Trace: design.sv:8599:19
						csr_rdata_int = (FPU == 1 ? {24'b000000000000000000000000, frm_q, fflags_q} : {32 {1'sb0}});
					12'h300:
						// Trace: design.sv:8602:9
						csr_rdata_int = {14'b00000000000000, mstatus_q[0], 4'b0000, mstatus_q[2-:2], 3'b000, mstatus_q[3], 2'h0, mstatus_q[4], mstatus_q[5], 2'h0, mstatus_q[6]};
					12'h301:
						// Trace: design.sv:8616:19
						csr_rdata_int = MISA_VALUE;
					12'h304:
						// Trace: design.sv:8619:11
						csr_rdata_int = mie_q;
					12'h305:
						// Trace: design.sv:8623:20
						csr_rdata_int = {mtvec_q, 6'h00, mtvec_mode_q};
					12'h340:
						// Trace: design.sv:8625:23
						csr_rdata_int = mscratch_q;
					12'h341:
						// Trace: design.sv:8627:19
						csr_rdata_int = mepc_q;
					12'h342:
						// Trace: design.sv:8629:21
						csr_rdata_int = {mcause_q[5], 26'b00000000000000000000000000, mcause_q[4:0]};
					12'h344:
						// Trace: design.sv:8632:11
						csr_rdata_int = mip;
					12'hf14:
						// Trace: design.sv:8635:22
						csr_rdata_int = hart_id_i;
					12'hf11:
						// Trace: design.sv:8638:24
						csr_rdata_int = {cv32e40p_pkg_MVENDORID_BANK, cv32e40p_pkg_MVENDORID_OFFSET};
					12'hf12:
						// Trace: design.sv:8641:22
						csr_rdata_int = cv32e40p_pkg_MARCHID;
					12'hf13, 12'h343:
						// Trace: design.sv:8644:32
						csr_rdata_int = 'b0;
					12'h7a0, 12'h7a3, 12'h7a8, 12'h7aa:
						// Trace: design.sv:8646:62
						csr_rdata_int = 'b0;
					12'h7a1:
						// Trace: design.sv:8647:21
						csr_rdata_int = tmatch_control_rdata;
					12'h7a2:
						// Trace: design.sv:8648:21
						csr_rdata_int = tmatch_value_rdata;
					12'h7a4:
						// Trace: design.sv:8649:20
						csr_rdata_int = tinfo_types;
					12'h7b0:
						// Trace: design.sv:8651:19
						csr_rdata_int = dcsr_q;
					12'h7b1:
						// Trace: design.sv:8652:18
						csr_rdata_int = depc_q;
					12'h7b2:
						// Trace: design.sv:8653:24
						csr_rdata_int = dscratch0_q;
					12'h7b3:
						// Trace: design.sv:8654:24
						csr_rdata_int = dscratch1_q;
					12'hb00, 12'hb02, 12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f, 12'hc00, 12'hc02, 12'hc03, 12'hc04, 12'hc05, 12'hc06, 12'hc07, 12'hc08, 12'hc09, 12'hc0a, 12'hc0b, 12'hc0c, 12'hc0d, 12'hc0e, 12'hc0f, 12'hc10, 12'hc11, 12'hc12, 12'hc13, 12'hc14, 12'hc15, 12'hc16, 12'hc17, 12'hc18, 12'hc19, 12'hc1a, 12'hc1b, 12'hc1c, 12'hc1d, 12'hc1e, 12'hc1f:
						// Trace: design.sv:8677:9
						csr_rdata_int = mhpmcounter_q[(csr_addr_i[4:0] * 64) + 31-:32];
					12'hb80, 12'hb82, 12'hb83, 12'hb84, 12'hb85, 12'hb86, 12'hb87, 12'hb88, 12'hb89, 12'hb8a, 12'hb8b, 12'hb8c, 12'hb8d, 12'hb8e, 12'hb8f, 12'hb90, 12'hb91, 12'hb92, 12'hb93, 12'hb94, 12'hb95, 12'hb96, 12'hb97, 12'hb98, 12'hb99, 12'hb9a, 12'hb9b, 12'hb9c, 12'hb9d, 12'hb9e, 12'hb9f, 12'hc80, 12'hc82, 12'hc83, 12'hc84, 12'hc85, 12'hc86, 12'hc87, 12'hc88, 12'hc89, 12'hc8a, 12'hc8b, 12'hc8c, 12'hc8d, 12'hc8e, 12'hc8f, 12'hc90, 12'hc91, 12'hc92, 12'hc93, 12'hc94, 12'hc95, 12'hc96, 12'hc97, 12'hc98, 12'hc99, 12'hc9a, 12'hc9b, 12'hc9c, 12'hc9d, 12'hc9e, 12'hc9f:
						// Trace: design.sv:8699:9
						csr_rdata_int = mhpmcounter_q[(csr_addr_i[4:0] * 64) + 63-:32];
					12'h320:
						// Trace: design.sv:8701:28
						csr_rdata_int = mcountinhibit_q;
					12'h323, 12'h324, 12'h325, 12'h326, 12'h327, 12'h328, 12'h329, 12'h32a, 12'h32b, 12'h32c, 12'h32d, 12'h32e, 12'h32f, 12'h330, 12'h331, 12'h332, 12'h333, 12'h334, 12'h335, 12'h336, 12'h337, 12'h338, 12'h339, 12'h33a, 12'h33b, 12'h33c, 12'h33d, 12'h33e, 12'h33f:
						// Trace: design.sv:8711:9
						csr_rdata_int = mhpmevent_q[csr_addr_i[4:0] * 32+:32];
					12'h800:
						// Trace: design.sv:8714:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_start_i[0+:32]);
					12'h801:
						// Trace: design.sv:8715:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_end_i[0+:32]);
					12'h802:
						// Trace: design.sv:8716:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_cnt_i[0+:32]);
					12'h804:
						// Trace: design.sv:8717:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_start_i[32+:32]);
					12'h805:
						// Trace: design.sv:8718:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_end_i[32+:32]);
					12'h806:
						// Trace: design.sv:8719:23
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hwlp_cnt_i[32+:32]);
					12'hcc0:
						// Trace: design.sv:8723:22
						csr_rdata_int = (!PULP_XPULP ? 'b0 : hart_id_i);
					12'hcc1:
						// Trace: design.sv:8725:21
						csr_rdata_int = (!PULP_XPULP ? 'b0 : {30'h00000000, priv_lvl_q});
					default:
						// Trace: design.sv:8726:18
						csr_rdata_int = 1'sb0;
				endcase
			end
		end
	endgenerate
	// Trace: design.sv:8731:3
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		if (PULP_SECURE == 1) begin : gen_pulp_secure_write_logic
			// Trace: design.sv:8733:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:8734:7
				fflags_n = fflags_q;
				// Trace: design.sv:8735:7
				frm_n = frm_q;
				// Trace: design.sv:8736:7
				mscratch_n = mscratch_q;
				// Trace: design.sv:8737:7
				mepc_n = mepc_q;
				// Trace: design.sv:8738:7
				uepc_n = uepc_q;
				// Trace: design.sv:8739:7
				depc_n = depc_q;
				// Trace: design.sv:8740:7
				dcsr_n = dcsr_q;
				// Trace: design.sv:8741:7
				dscratch0_n = dscratch0_q;
				// Trace: design.sv:8742:7
				dscratch1_n = dscratch1_q;
				// Trace: design.sv:8744:7
				mstatus_n = mstatus_q;
				// Trace: design.sv:8745:7
				mcause_n = mcause_q;
				// Trace: design.sv:8746:7
				ucause_n = ucause_q;
				// Trace: design.sv:8747:7
				hwlp_we_o = 1'sb0;
				// Trace: design.sv:8748:7
				hwlp_regid_o = 1'sb0;
				// Trace: design.sv:8749:7
				exception_pc = pc_id_i;
				// Trace: design.sv:8750:7
				priv_lvl_n = priv_lvl_q;
				// Trace: design.sv:8751:7
				mtvec_n = (csr_mtvec_init_i ? mtvec_addr_i[31:8] : mtvec_q);
				// Trace: design.sv:8752:7
				utvec_n = utvec_q;
				// Trace: design.sv:8753:7
				mtvec_mode_n = mtvec_mode_q;
				// Trace: design.sv:8754:7
				utvec_mode_n = utvec_mode_q;
				// Trace: design.sv:8755:7
				pmp_reg_n[767-:512] = pmp_reg_q[767-:512];
				// Trace: design.sv:8756:7
				pmp_reg_n[255-:128] = pmp_reg_q[255-:128];
				// Trace: design.sv:8757:7
				pmpaddr_we = 1'sb0;
				// Trace: design.sv:8758:7
				pmpcfg_we = 1'sb0;
				// Trace: design.sv:8760:7
				mie_n = mie_q;
				// Trace: design.sv:8762:7
				if (FPU == 1) begin
					if (fflags_we_i)
						// Trace: design.sv:8762:38
						fflags_n = fflags_i | fflags_q;
				end
				case (csr_addr_i)
					12'h001:
						if (csr_we_int)
							// Trace: design.sv:8766:37
							fflags_n = (FPU == 1 ? csr_wdata_int[4:0] : {5 {1'sb0}});
					12'h002:
						if (csr_we_int)
							// Trace: design.sv:8767:37
							frm_n = (FPU == 1 ? csr_wdata_int[2:0] : {3 {1'sb0}});
					12'h003:
						if (csr_we_int) begin
							// Trace: design.sv:8770:11
							fflags_n = (FPU == 1 ? csr_wdata_int[4:0] : {5 {1'sb0}});
							// Trace: design.sv:8771:11
							frm_n = (FPU == 1 ? csr_wdata_int[7:cv32e40p_pkg_C_FFLAG] : {3 {1'sb0}});
						end
					12'h300:
						if (csr_we_int)
							// Trace: design.sv:8777:11
							mstatus_n = {csr_wdata_int[MSTATUS_UIE_BIT], csr_wdata_int[MSTATUS_MIE_BIT], csr_wdata_int[MSTATUS_UPIE_BIT], csr_wdata_int[MSTATUS_MPIE_BIT], sv2v_cast_2(csr_wdata_int[MSTATUS_MPP_BIT_HIGH:MSTATUS_MPP_BIT_LOW]), csr_wdata_int[MSTATUS_MPRV_BIT]};
					12'h304:
						if (csr_we_int)
							// Trace: design.sv:8789:11
							mie_n = csr_wdata_int & cv32e40p_pkg_IRQ_MASK;
					12'h305:
						if (csr_we_int) begin
							// Trace: design.sv:8794:11
							mtvec_n = csr_wdata_int[31:8];
							// Trace: design.sv:8795:11
							mtvec_mode_n = {1'b0, csr_wdata_int[0]};
						end
					12'h340:
						if (csr_we_int)
							// Trace: design.sv:8800:11
							mscratch_n = csr_wdata_int;
					12'h341:
						if (csr_we_int)
							// Trace: design.sv:8805:11
							mepc_n = csr_wdata_int & ~32'b00000000000000000000000000000001;
					12'h342:
						if (csr_we_int)
							// Trace: design.sv:8808:37
							mcause_n = {csr_wdata_int[31], csr_wdata_int[4:0]};
					12'h7b0:
						if (csr_we_int) begin
							// Trace: design.sv:8819:11
							dcsr_n[15] = csr_wdata_int[15];
							// Trace: design.sv:8820:11
							dcsr_n[13] = 1'b0;
							// Trace: design.sv:8821:11
							dcsr_n[12] = csr_wdata_int[12];
							// Trace: design.sv:8822:11
							dcsr_n[11] = csr_wdata_int[11];
							// Trace: design.sv:8823:11
							dcsr_n[10] = 1'b0;
							// Trace: design.sv:8824:11
							dcsr_n[9] = 1'b0;
							// Trace: design.sv:8825:11
							dcsr_n[4] = 1'b0;
							// Trace: design.sv:8826:11
							dcsr_n[2] = csr_wdata_int[2];
							// Trace: design.sv:8827:11
							dcsr_n[1-:2] = (csr_wdata_int[1:0] == 2'b11 ? 2'b11 : 2'b00);
						end
					12'h7b1:
						if (csr_we_int)
							// Trace: design.sv:8832:11
							depc_n = csr_wdata_int & ~32'b00000000000000000000000000000001;
					12'h7b2:
						if (csr_we_int)
							// Trace: design.sv:8837:11
							dscratch0_n = csr_wdata_int;
					12'h7b3:
						if (csr_we_int)
							// Trace: design.sv:8842:11
							dscratch1_n = csr_wdata_int;
					12'h800:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:8848:11
							hwlp_we_o = 3'b001;
							// Trace: design.sv:8849:11
							hwlp_regid_o = 1'b0;
						end
					12'h801:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:8853:11
							hwlp_we_o = 3'b010;
							// Trace: design.sv:8854:11
							hwlp_regid_o = 1'b0;
						end
					12'h802:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:8858:11
							hwlp_we_o = 3'b100;
							// Trace: design.sv:8859:11
							hwlp_regid_o = 1'b0;
						end
					12'h804:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:8863:11
							hwlp_we_o = 3'b001;
							// Trace: design.sv:8864:11
							hwlp_regid_o = 1'b1;
						end
					12'h805:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:8868:11
							hwlp_we_o = 3'b010;
							// Trace: design.sv:8869:11
							hwlp_regid_o = 1'b1;
						end
					12'h806:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:8873:11
							hwlp_we_o = 3'b100;
							// Trace: design.sv:8874:11
							hwlp_regid_o = 1'b1;
						end
					12'h3a0:
						if (csr_we_int) begin
							// Trace: design.sv:8880:11
							pmp_reg_n[128+:32] = csr_wdata_int;
							// Trace: design.sv:8881:11
							pmpcfg_we[3:0] = 4'b1111;
						end
					12'h3a1:
						if (csr_we_int) begin
							// Trace: design.sv:8885:11
							pmp_reg_n[160+:32] = csr_wdata_int;
							// Trace: design.sv:8886:11
							pmpcfg_we[7:4] = 4'b1111;
						end
					12'h3a2:
						if (csr_we_int) begin
							// Trace: design.sv:8890:11
							pmp_reg_n[192+:32] = csr_wdata_int;
							// Trace: design.sv:8891:11
							pmpcfg_we[11:8] = 4'b1111;
						end
					12'h3a3:
						if (csr_we_int) begin
							// Trace: design.sv:8895:11
							pmp_reg_n[224+:32] = csr_wdata_int;
							// Trace: design.sv:8896:11
							pmpcfg_we[15:12] = 4'b1111;
						end
					12'h3b0, 12'h3b1, 12'h3b2, 12'h3b3, 12'h3b4, 12'h3b5, 12'h3b6, 12'h3b7, 12'h3b8, 12'h3b9, 12'h3ba, 12'h3bb, 12'h3bc, 12'h3bd, 12'h3be, 12'h3bf:
						if (csr_we_int) begin
							// Trace: design.sv:8904:11
							pmp_reg_n[256 + (csr_addr_i[3:0] * 32)+:32] = csr_wdata_int;
							// Trace: design.sv:8905:11
							pmpaddr_we[csr_addr_i[3:0]] = 1'b1;
						end
					12'h000:
						if (csr_we_int)
							// Trace: design.sv:8913:11
							mstatus_n = {csr_wdata_int[MSTATUS_UIE_BIT], mstatus_q[5], csr_wdata_int[MSTATUS_UPIE_BIT], mstatus_q[3], sv2v_cast_2(mstatus_q[2-:2]), mstatus_q[0]};
					12'h005:
						if (csr_we_int) begin
							// Trace: design.sv:8925:11
							utvec_n = csr_wdata_int[31:8];
							// Trace: design.sv:8926:11
							utvec_mode_n = {1'b0, csr_wdata_int[0]};
						end
					12'h041:
						if (csr_we_int)
							// Trace: design.sv:8931:11
							uepc_n = csr_wdata_int;
					12'h042:
						if (csr_we_int)
							// Trace: design.sv:8934:37
							ucause_n = {csr_wdata_int[31], csr_wdata_int[4:0]};
				endcase
				(* full_case, parallel_case *)
				case (1'b1)
					csr_save_cause_i: begin
						// Trace: design.sv:8942:11
						(* full_case, parallel_case *)
						case (1'b1)
							csr_save_if_i:
								// Trace: design.sv:8943:28
								exception_pc = pc_if_i;
							csr_save_id_i:
								// Trace: design.sv:8944:28
								exception_pc = pc_id_i;
							csr_save_ex_i:
								// Trace: design.sv:8945:28
								exception_pc = pc_ex_i;
							default:
								;
						endcase
						(* full_case, parallel_case *)
						case (priv_lvl_q)
							2'b00:
								// Trace: design.sv:8952:15
								if (~is_irq) begin
									// Trace: design.sv:8954:17
									priv_lvl_n = 2'b11;
									// Trace: design.sv:8955:17
									mstatus_n[3] = mstatus_q[6];
									// Trace: design.sv:8956:17
									mstatus_n[5] = 1'b0;
									// Trace: design.sv:8957:17
									mstatus_n[2-:2] = 2'b00;
									// Trace: design.sv:8958:17
									if (debug_csr_save_i)
										// Trace: design.sv:8958:39
										depc_n = exception_pc;
									else
										// Trace: design.sv:8959:22
										mepc_n = exception_pc;
									// Trace: design.sv:8960:17
									mcause_n = csr_cause_i;
								end
								else
									// Trace: design.sv:8963:17
									if (~csr_irq_sec_i) begin
										// Trace: design.sv:8965:19
										priv_lvl_n = 2'b00;
										// Trace: design.sv:8966:19
										mstatus_n[4] = mstatus_q[6];
										// Trace: design.sv:8967:19
										mstatus_n[6] = 1'b0;
										// Trace: design.sv:8968:19
										if (debug_csr_save_i)
											// Trace: design.sv:8968:41
											depc_n = exception_pc;
										else
											// Trace: design.sv:8969:24
											uepc_n = exception_pc;
										// Trace: design.sv:8970:19
										ucause_n = csr_cause_i;
									end
									else begin
										// Trace: design.sv:8974:19
										priv_lvl_n = 2'b11;
										// Trace: design.sv:8975:19
										mstatus_n[3] = mstatus_q[6];
										// Trace: design.sv:8976:19
										mstatus_n[5] = 1'b0;
										// Trace: design.sv:8977:19
										mstatus_n[2-:2] = 2'b00;
										// Trace: design.sv:8978:19
										if (debug_csr_save_i)
											// Trace: design.sv:8978:41
											depc_n = exception_pc;
										else
											// Trace: design.sv:8979:24
											mepc_n = exception_pc;
										// Trace: design.sv:8980:19
										mcause_n = csr_cause_i;
									end
							2'b11:
								// Trace: design.sv:8986:15
								if (debug_csr_save_i) begin
									// Trace: design.sv:8989:17
									dcsr_n[1-:2] = 2'b11;
									// Trace: design.sv:8990:17
									dcsr_n[8-:3] = debug_cause_i;
									// Trace: design.sv:8991:17
									depc_n = exception_pc;
								end
								else begin
									// Trace: design.sv:8994:17
									priv_lvl_n = 2'b11;
									// Trace: design.sv:8995:17
									mstatus_n[3] = mstatus_q[5];
									// Trace: design.sv:8996:17
									mstatus_n[5] = 1'b0;
									// Trace: design.sv:8997:17
									mstatus_n[2-:2] = 2'b11;
									// Trace: design.sv:8998:17
									mepc_n = exception_pc;
									// Trace: design.sv:8999:17
									mcause_n = csr_cause_i;
								end
							default:
								;
						endcase
					end
					csr_restore_uret_i: begin
						// Trace: design.sv:9010:11
						mstatus_n[6] = mstatus_q[4];
						// Trace: design.sv:9011:11
						priv_lvl_n = 2'b00;
						// Trace: design.sv:9012:11
						mstatus_n[4] = 1'b1;
					end
					csr_restore_mret_i:
						// Trace: design.sv:9016:11
						(* full_case, parallel_case *)
						case (mstatus_q[2-:2])
							2'b00: begin
								// Trace: design.sv:9018:15
								mstatus_n[6] = mstatus_q[3];
								// Trace: design.sv:9019:15
								priv_lvl_n = 2'b00;
								// Trace: design.sv:9020:15
								mstatus_n[3] = 1'b1;
								// Trace: design.sv:9021:15
								mstatus_n[2-:2] = 2'b00;
							end
							2'b11: begin
								// Trace: design.sv:9024:15
								mstatus_n[5] = mstatus_q[3];
								// Trace: design.sv:9025:15
								priv_lvl_n = 2'b11;
								// Trace: design.sv:9026:15
								mstatus_n[3] = 1'b1;
								// Trace: design.sv:9027:15
								mstatus_n[2-:2] = 2'b00;
							end
							default:
								;
						endcase
					csr_restore_dret_i:
						// Trace: design.sv:9036:11
						priv_lvl_n = dcsr_q[1-:2];
					default:
						;
				endcase
			end
		end
		else begin : gen_no_pulp_secure_write_logic
			// Trace: design.sv:9045:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:9046:7
				fflags_n = fflags_q;
				// Trace: design.sv:9047:7
				frm_n = frm_q;
				// Trace: design.sv:9048:7
				mscratch_n = mscratch_q;
				// Trace: design.sv:9049:7
				mepc_n = mepc_q;
				// Trace: design.sv:9050:7
				uepc_n = 'b0;
				// Trace: design.sv:9051:7
				depc_n = depc_q;
				// Trace: design.sv:9052:7
				dcsr_n = dcsr_q;
				// Trace: design.sv:9053:7
				dscratch0_n = dscratch0_q;
				// Trace: design.sv:9054:7
				dscratch1_n = dscratch1_q;
				// Trace: design.sv:9056:7
				mstatus_n = mstatus_q;
				// Trace: design.sv:9057:7
				mcause_n = mcause_q;
				// Trace: design.sv:9058:7
				ucause_n = 1'sb0;
				// Trace: design.sv:9059:7
				hwlp_we_o = 1'sb0;
				// Trace: design.sv:9060:7
				hwlp_regid_o = 1'sb0;
				// Trace: design.sv:9061:7
				exception_pc = pc_id_i;
				// Trace: design.sv:9062:7
				priv_lvl_n = priv_lvl_q;
				// Trace: design.sv:9063:7
				mtvec_n = (csr_mtvec_init_i ? mtvec_addr_i[31:8] : mtvec_q);
				// Trace: design.sv:9064:7
				utvec_n = 1'sb0;
				// Trace: design.sv:9065:7
				pmp_reg_n[767-:512] = 1'sb0;
				// Trace: design.sv:9066:7
				pmp_reg_n[255-:128] = 1'sb0;
				// Trace: design.sv:9067:7
				pmp_reg_n[127-:128] = 1'sb0;
				// Trace: design.sv:9068:7
				pmpaddr_we = 1'sb0;
				// Trace: design.sv:9069:7
				pmpcfg_we = 1'sb0;
				// Trace: design.sv:9071:7
				mie_n = mie_q;
				// Trace: design.sv:9072:7
				mtvec_mode_n = mtvec_mode_q;
				// Trace: design.sv:9073:7
				utvec_mode_n = 1'sb0;
				// Trace: design.sv:9075:7
				if (FPU == 1) begin
					if (fflags_we_i)
						// Trace: design.sv:9075:38
						fflags_n = fflags_i | fflags_q;
				end
				case (csr_addr_i)
					12'h001:
						if (csr_we_int)
							// Trace: design.sv:9079:37
							fflags_n = (FPU == 1 ? csr_wdata_int[4:0] : {5 {1'sb0}});
					12'h002:
						if (csr_we_int)
							// Trace: design.sv:9080:37
							frm_n = (FPU == 1 ? csr_wdata_int[2:0] : {3 {1'sb0}});
					12'h003:
						if (csr_we_int) begin
							// Trace: design.sv:9083:11
							fflags_n = (FPU == 1 ? csr_wdata_int[4:0] : {5 {1'sb0}});
							// Trace: design.sv:9084:11
							frm_n = (FPU == 1 ? csr_wdata_int[7:cv32e40p_pkg_C_FFLAG] : {3 {1'sb0}});
						end
					12'h300:
						if (csr_we_int)
							// Trace: design.sv:9090:11
							mstatus_n = {csr_wdata_int[MSTATUS_UIE_BIT], csr_wdata_int[MSTATUS_MIE_BIT], csr_wdata_int[MSTATUS_UPIE_BIT], csr_wdata_int[MSTATUS_MPIE_BIT], sv2v_cast_2(csr_wdata_int[MSTATUS_MPP_BIT_HIGH:MSTATUS_MPP_BIT_LOW]), csr_wdata_int[MSTATUS_MPRV_BIT]};
					12'h304:
						if (csr_we_int)
							// Trace: design.sv:9102:11
							mie_n = csr_wdata_int & cv32e40p_pkg_IRQ_MASK;
					12'h305:
						if (csr_we_int) begin
							// Trace: design.sv:9107:11
							mtvec_n = csr_wdata_int[31:8];
							// Trace: design.sv:9108:11
							mtvec_mode_n = {1'b0, csr_wdata_int[0]};
						end
					12'h340:
						if (csr_we_int)
							// Trace: design.sv:9113:11
							mscratch_n = csr_wdata_int;
					12'h341:
						if (csr_we_int)
							// Trace: design.sv:9118:11
							mepc_n = csr_wdata_int & ~32'b00000000000000000000000000000001;
					12'h342:
						if (csr_we_int)
							// Trace: design.sv:9121:37
							mcause_n = {csr_wdata_int[31], csr_wdata_int[4:0]};
					12'h7b0:
						if (csr_we_int) begin
							// Trace: design.sv:9131:11
							dcsr_n[15] = csr_wdata_int[15];
							// Trace: design.sv:9132:11
							dcsr_n[13] = 1'b0;
							// Trace: design.sv:9133:11
							dcsr_n[12] = 1'b0;
							// Trace: design.sv:9134:11
							dcsr_n[11] = csr_wdata_int[11];
							// Trace: design.sv:9135:11
							dcsr_n[10] = 1'b0;
							// Trace: design.sv:9136:11
							dcsr_n[9] = 1'b0;
							// Trace: design.sv:9137:11
							dcsr_n[4] = 1'b0;
							// Trace: design.sv:9138:11
							dcsr_n[2] = csr_wdata_int[2];
							// Trace: design.sv:9139:11
							dcsr_n[1-:2] = 2'b11;
						end
					12'h7b1:
						if (csr_we_int)
							// Trace: design.sv:9144:11
							depc_n = csr_wdata_int & ~32'b00000000000000000000000000000001;
					12'h7b2:
						if (csr_we_int)
							// Trace: design.sv:9149:11
							dscratch0_n = csr_wdata_int;
					12'h7b3:
						if (csr_we_int)
							// Trace: design.sv:9154:11
							dscratch1_n = csr_wdata_int;
					12'h800:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:9160:11
							hwlp_we_o = 3'b001;
							// Trace: design.sv:9161:11
							hwlp_regid_o = 1'b0;
						end
					12'h801:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:9165:11
							hwlp_we_o = 3'b010;
							// Trace: design.sv:9166:11
							hwlp_regid_o = 1'b0;
						end
					12'h802:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:9170:11
							hwlp_we_o = 3'b100;
							// Trace: design.sv:9171:11
							hwlp_regid_o = 1'b0;
						end
					12'h804:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:9175:11
							hwlp_we_o = 3'b001;
							// Trace: design.sv:9176:11
							hwlp_regid_o = 1'b1;
						end
					12'h805:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:9180:11
							hwlp_we_o = 3'b010;
							// Trace: design.sv:9181:11
							hwlp_regid_o = 1'b1;
						end
					12'h806:
						if (PULP_XPULP && csr_we_int) begin
							// Trace: design.sv:9185:11
							hwlp_we_o = 3'b100;
							// Trace: design.sv:9186:11
							hwlp_regid_o = 1'b1;
						end
				endcase
				(* full_case, parallel_case *)
				case (1'b1)
					csr_save_cause_i: begin
						// Trace: design.sv:9194:11
						(* full_case, parallel_case *)
						case (1'b1)
							csr_save_if_i:
								// Trace: design.sv:9195:28
								exception_pc = pc_if_i;
							csr_save_id_i:
								// Trace: design.sv:9196:28
								exception_pc = pc_id_i;
							csr_save_ex_i:
								// Trace: design.sv:9197:28
								exception_pc = pc_ex_i;
							default:
								;
						endcase
						if (debug_csr_save_i) begin
							// Trace: design.sv:9204:13
							dcsr_n[1-:2] = 2'b11;
							// Trace: design.sv:9205:13
							dcsr_n[8-:3] = debug_cause_i;
							// Trace: design.sv:9206:13
							depc_n = exception_pc;
						end
						else begin
							// Trace: design.sv:9208:13
							priv_lvl_n = 2'b11;
							// Trace: design.sv:9209:13
							mstatus_n[3] = mstatus_q[5];
							// Trace: design.sv:9210:13
							mstatus_n[5] = 1'b0;
							// Trace: design.sv:9211:13
							mstatus_n[2-:2] = 2'b11;
							// Trace: design.sv:9212:13
							mepc_n = exception_pc;
							// Trace: design.sv:9213:13
							mcause_n = csr_cause_i;
						end
					end
					csr_restore_mret_i: begin
						// Trace: design.sv:9218:11
						mstatus_n[5] = mstatus_q[3];
						// Trace: design.sv:9219:11
						priv_lvl_n = 2'b11;
						// Trace: design.sv:9220:11
						mstatus_n[3] = 1'b1;
						// Trace: design.sv:9221:11
						mstatus_n[2-:2] = 2'b11;
					end
					csr_restore_dret_i:
						// Trace: design.sv:9226:11
						priv_lvl_n = dcsr_q[1-:2];
					default:
						;
				endcase
			end
		end
	endgenerate
	// Trace: design.sv:9234:3
	assign hwlp_data_o = (PULP_XPULP ? csr_wdata_int : {32 {1'sb0}});
	// Trace: design.sv:9237:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:9238:5
		csr_wdata_int = csr_wdata_i;
		// Trace: design.sv:9239:5
		csr_we_int = 1'b1;
		// Trace: design.sv:9241:5
		case (csr_op_i)
			sv2v_cast_EB06E(2'b01):
				// Trace: design.sv:9242:21
				csr_wdata_int = csr_wdata_i;
			sv2v_cast_EB06E(2'b10):
				// Trace: design.sv:9243:21
				csr_wdata_int = csr_wdata_i | csr_rdata_o;
			sv2v_cast_EB06E(2'b11):
				// Trace: design.sv:9244:21
				csr_wdata_int = ~csr_wdata_i & csr_rdata_o;
			sv2v_cast_EB06E(2'b00): begin
				// Trace: design.sv:9247:9
				csr_wdata_int = csr_wdata_i;
				// Trace: design.sv:9248:9
				csr_we_int = 1'b0;
			end
		endcase
	end
	// Trace: design.sv:9253:3
	assign csr_rdata_o = csr_rdata_int;
	// Trace: design.sv:9256:3
	assign m_irq_enable_o = mstatus_q[5] && !(dcsr_q[2] && !dcsr_q[11]);
	// Trace: design.sv:9257:3
	assign u_irq_enable_o = mstatus_q[6] && !(dcsr_q[2] && !dcsr_q[11]);
	// Trace: design.sv:9258:3
	assign priv_lvl_o = priv_lvl_q;
	// Trace: design.sv:9259:3
	assign sec_lvl_o = priv_lvl_q[0];
	// Trace: design.sv:9260:3
	assign frm_o = (FPU == 1 ? frm_q : {3 {1'sb0}});
	// Trace: design.sv:9262:3
	assign mtvec_o = mtvec_q;
	// Trace: design.sv:9263:3
	assign utvec_o = utvec_q;
	// Trace: design.sv:9264:3
	assign mtvec_mode_o = mtvec_mode_q;
	// Trace: design.sv:9265:3
	assign utvec_mode_o = utvec_mode_q;
	// Trace: design.sv:9267:3
	assign mepc_o = mepc_q;
	// Trace: design.sv:9268:3
	assign uepc_o = uepc_q;
	// Trace: design.sv:9270:3
	assign mcounteren_o = (PULP_SECURE ? mcounteren_q : {32 {1'sb0}});
	// Trace: design.sv:9272:3
	assign depc_o = depc_q;
	// Trace: design.sv:9274:3
	assign pmp_addr_o = pmp_reg_q[767-:512];
	// Trace: design.sv:9275:3
	assign pmp_cfg_o = pmp_reg_q[127-:128];
	// Trace: design.sv:9277:3
	assign debug_single_step_o = dcsr_q[2];
	// Trace: design.sv:9278:3
	assign debug_ebreakm_o = dcsr_q[15];
	// Trace: design.sv:9279:3
	assign debug_ebreaku_o = dcsr_q[12];
	// Trace: design.sv:9281:3
	generate
		if (PULP_SECURE == 1) begin : gen_pmp_user
			for (_gv_j_3 = 0; _gv_j_3 < N_PMP_ENTRIES; _gv_j_3 = _gv_j_3 + 1) begin : CS_PMP_CFG
				localparam j = _gv_j_3;
				// Trace: design.sv:9285:9
				wire [8:1] sv2v_tmp_9A7A7;
				assign sv2v_tmp_9A7A7 = pmp_reg_n[128 + (((j / 4) * 32) + (((8 * ((j % 4) + 1)) - 1) >= (8 * (j % 4)) ? (8 * ((j % 4) + 1)) - 1 : (((8 * ((j % 4) + 1)) - 1) + (((8 * ((j % 4) + 1)) - 1) >= (8 * (j % 4)) ? (((8 * ((j % 4) + 1)) - 1) - (8 * (j % 4))) + 1 : ((8 * (j % 4)) - ((8 * ((j % 4) + 1)) - 1)) + 1)) - 1))-:(((8 * ((j % 4) + 1)) - 1) >= (8 * (j % 4)) ? (((8 * ((j % 4) + 1)) - 1) - (8 * (j % 4))) + 1 : ((8 * (j % 4)) - ((8 * ((j % 4) + 1)) - 1)) + 1)];
				always @(*) pmp_reg_n[0 + (j * 8)+:8] = sv2v_tmp_9A7A7;
				// Trace: design.sv:9286:9
				wire [(((8 * ((j % 4) + 1)) - 1) >= (8 * (j % 4)) ? (((8 * ((j % 4) + 1)) - 1) - (8 * (j % 4))) + 1 : ((8 * (j % 4)) - ((8 * ((j % 4) + 1)) - 1)) + 1) * 1:1] sv2v_tmp_D6B27;
				assign sv2v_tmp_D6B27 = pmp_reg_q[0 + (j * 8)+:8];
				always @(*) pmp_reg_q[128 + (((j / 4) * 32) + (((8 * ((j % 4) + 1)) - 1) >= (8 * (j % 4)) ? (8 * ((j % 4) + 1)) - 1 : (((8 * ((j % 4) + 1)) - 1) + (((8 * ((j % 4) + 1)) - 1) >= (8 * (j % 4)) ? (((8 * ((j % 4) + 1)) - 1) - (8 * (j % 4))) + 1 : ((8 * (j % 4)) - ((8 * ((j % 4) + 1)) - 1)) + 1)) - 1))-:(((8 * ((j % 4) + 1)) - 1) >= (8 * (j % 4)) ? (((8 * ((j % 4) + 1)) - 1) - (8 * (j % 4))) + 1 : ((8 * (j % 4)) - ((8 * ((j % 4) + 1)) - 1)) + 1)] = sv2v_tmp_D6B27;
			end
			for (_gv_j_3 = 0; _gv_j_3 < N_PMP_ENTRIES; _gv_j_3 = _gv_j_3 + 1) begin : CS_PMP_REGS_FF
				localparam j = _gv_j_3;
				// Trace: design.sv:9290:9
				always @(posedge clk or negedge rst_n)
					// Trace: design.sv:9291:11
					if (rst_n == 1'b0) begin
						// Trace: design.sv:9292:13
						pmp_reg_q[0 + (j * 8)+:8] <= 1'sb0;
						// Trace: design.sv:9293:13
						pmp_reg_q[256 + (j * 32)+:32] <= 1'sb0;
					end
					else begin
						// Trace: design.sv:9295:13
						if (pmpcfg_we[j])
							// Trace: design.sv:9295:31
							pmp_reg_q[0 + (j * 8)+:8] <= (USE_PMP ? pmp_reg_n[0 + (j * 8)+:8] : {8 {1'sb0}});
						if (pmpaddr_we[j])
							// Trace: design.sv:9296:32
							pmp_reg_q[256 + (j * 32)+:32] <= (USE_PMP ? pmp_reg_n[256 + (j * 32)+:32] : {32 {1'sb0}});
					end
			end
			// Trace: design.sv:9301:7
			always @(posedge clk or negedge rst_n)
				// Trace: design.sv:9302:9
				if (rst_n == 1'b0) begin
					// Trace: design.sv:9303:11
					uepc_q <= 1'sb0;
					// Trace: design.sv:9304:11
					ucause_q <= 1'sb0;
					// Trace: design.sv:9305:11
					utvec_q <= 1'sb0;
					// Trace: design.sv:9306:11
					utvec_mode_q <= MTVEC_MODE;
					// Trace: design.sv:9307:11
					priv_lvl_q <= 2'b11;
				end
				else begin
					// Trace: design.sv:9309:11
					uepc_q <= uepc_n;
					// Trace: design.sv:9310:11
					ucause_q <= ucause_n;
					// Trace: design.sv:9311:11
					utvec_q <= utvec_n;
					// Trace: design.sv:9312:11
					utvec_mode_q <= utvec_mode_n;
					// Trace: design.sv:9313:11
					priv_lvl_q <= priv_lvl_n;
				end
		end
		else begin : gen_no_pmp_user
			// Trace: design.sv:9317:7
			wire [768:1] sv2v_tmp_E1062;
			assign sv2v_tmp_E1062 = 1'sb0;
			always @(*) pmp_reg_q = sv2v_tmp_E1062;
			// Trace: design.sv:9318:7
			wire [32:1] sv2v_tmp_1316C;
			assign sv2v_tmp_1316C = 1'sb0;
			always @(*) uepc_q = sv2v_tmp_1316C;
			// Trace: design.sv:9319:7
			wire [6:1] sv2v_tmp_55E05;
			assign sv2v_tmp_55E05 = 1'sb0;
			always @(*) ucause_q = sv2v_tmp_55E05;
			// Trace: design.sv:9320:7
			wire [24:1] sv2v_tmp_382EF;
			assign sv2v_tmp_382EF = 1'sb0;
			always @(*) utvec_q = sv2v_tmp_382EF;
			// Trace: design.sv:9321:7
			wire [2:1] sv2v_tmp_828F8;
			assign sv2v_tmp_828F8 = 1'sb0;
			always @(*) utvec_mode_q = sv2v_tmp_828F8;
			// Trace: design.sv:9322:7
			wire [2:1] sv2v_tmp_86FE7;
			assign sv2v_tmp_86FE7 = 2'b11;
			always @(*) priv_lvl_q = sv2v_tmp_86FE7;
		end
	endgenerate
	// Trace: design.sv:9327:3
	localparam cv32e40p_pkg_DBG_CAUSE_NONE = 3'h0;
	// removed localparam type cv32e40p_pkg_x_debug_ver_e
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:9328:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:9329:7
			frm_q <= 1'sb0;
			// Trace: design.sv:9330:7
			fflags_q <= 1'sb0;
			// Trace: design.sv:9331:7
			mstatus_q <= 7'b0000110;
			// Trace: design.sv:9339:7
			mepc_q <= 1'sb0;
			// Trace: design.sv:9340:7
			mcause_q <= 1'sb0;
			// Trace: design.sv:9342:7
			depc_q <= 1'sb0;
			// Trace: design.sv:9343:7
			dcsr_q <= {23'h200000, cv32e40p_pkg_DBG_CAUSE_NONE, 6'b000011};
			// Trace: design.sv:9349:7
			dscratch0_q <= 1'sb0;
			// Trace: design.sv:9350:7
			dscratch1_q <= 1'sb0;
			// Trace: design.sv:9351:7
			mscratch_q <= 1'sb0;
			// Trace: design.sv:9352:7
			mie_q <= 1'sb0;
			// Trace: design.sv:9353:7
			mtvec_q <= 1'sb0;
			// Trace: design.sv:9354:7
			mtvec_mode_q <= MTVEC_MODE;
		end
		else begin
			// Trace: design.sv:9357:7
			if (FPU == 1) begin
				// Trace: design.sv:9358:9
				frm_q <= frm_n;
				// Trace: design.sv:9359:9
				fflags_q <= fflags_n;
			end
			else begin
				// Trace: design.sv:9361:9
				frm_q <= 'b0;
				// Trace: design.sv:9362:9
				fflags_q <= 'b0;
			end
			if (PULP_SECURE == 1)
				// Trace: design.sv:9365:9
				mstatus_q <= mstatus_n;
			else
				// Trace: design.sv:9367:9
				mstatus_q <= {1'b0, mstatus_n[5], 1'b0, mstatus_n[3], 3'b110};
			// Trace: design.sv:9376:7
			mepc_q <= mepc_n;
			// Trace: design.sv:9377:7
			mcause_q <= mcause_n;
			// Trace: design.sv:9378:7
			depc_q <= depc_n;
			// Trace: design.sv:9379:7
			dcsr_q <= dcsr_n;
			// Trace: design.sv:9380:7
			dscratch0_q <= dscratch0_n;
			// Trace: design.sv:9381:7
			dscratch1_q <= dscratch1_n;
			// Trace: design.sv:9382:7
			mscratch_q <= mscratch_n;
			// Trace: design.sv:9383:7
			mie_q <= mie_n;
			// Trace: design.sv:9384:7
			mtvec_q <= mtvec_n;
			// Trace: design.sv:9385:7
			mtvec_mode_q <= mtvec_mode_n;
		end
	// Trace: design.sv:9397:3
	// removed localparam type cv32e40p_pkg_trigger_type_e
	generate
		if (DEBUG_TRIGGER_EN) begin : gen_trigger_regs
			// Trace: design.sv:9399:5
			reg tmatch_control_exec_q;
			// Trace: design.sv:9400:5
			reg [31:0] tmatch_value_q;
			// Trace: design.sv:9402:5
			wire tmatch_control_we;
			// Trace: design.sv:9403:5
			wire tmatch_value_we;
			// Trace: design.sv:9406:5
			assign tmatch_control_we = (csr_we_int & debug_mode_i) & (csr_addr_i == 12'h7a1);
			// Trace: design.sv:9407:5
			assign tmatch_value_we = (csr_we_int & debug_mode_i) & (csr_addr_i == 12'h7a2);
			// Trace: design.sv:9411:5
			always @(posedge clk or negedge rst_n)
				// Trace: design.sv:9412:7
				if (!rst_n) begin
					// Trace: design.sv:9413:9
					tmatch_control_exec_q <= 'b0;
					// Trace: design.sv:9414:9
					tmatch_value_q <= 'b0;
				end
				else begin
					// Trace: design.sv:9416:9
					if (tmatch_control_we)
						// Trace: design.sv:9416:32
						tmatch_control_exec_q <= csr_wdata_int[2];
					if (tmatch_value_we)
						// Trace: design.sv:9417:30
						tmatch_value_q <= csr_wdata_int[31:0];
				end
			// Trace: design.sv:9422:5
			assign tinfo_types = 4;
			// Trace: design.sv:9426:5
			assign tmatch_control_rdata = {28'h2800104, PULP_SECURE == 1, tmatch_control_exec_q, 2'b00};
			// Trace: design.sv:9447:5
			assign tmatch_value_rdata = tmatch_value_q;
			// Trace: design.sv:9451:5
			assign trigger_match_o = tmatch_control_exec_q & (pc_id_i[31:0] == tmatch_value_q[31:0]);
		end
		else begin : gen_no_trigger_regs
			// Trace: design.sv:9454:5
			assign tinfo_types = 'b0;
			// Trace: design.sv:9455:5
			assign tmatch_control_rdata = 'b0;
			// Trace: design.sv:9456:5
			assign tmatch_value_rdata = 'b0;
			// Trace: design.sv:9457:5
			assign trigger_match_o = 'b0;
		end
	endgenerate
	// Trace: design.sv:9471:3
	assign hpm_events[0] = 1'b1;
	// Trace: design.sv:9472:3
	assign hpm_events[1] = mhpmevent_minstret_i;
	// Trace: design.sv:9473:3
	assign hpm_events[2] = mhpmevent_ld_stall_i;
	// Trace: design.sv:9474:3
	assign hpm_events[3] = mhpmevent_jr_stall_i;
	// Trace: design.sv:9475:3
	assign hpm_events[4] = mhpmevent_imiss_i;
	// Trace: design.sv:9476:3
	assign hpm_events[5] = mhpmevent_load_i;
	// Trace: design.sv:9477:3
	assign hpm_events[6] = mhpmevent_store_i;
	// Trace: design.sv:9478:3
	assign hpm_events[7] = mhpmevent_jump_i;
	// Trace: design.sv:9479:3
	assign hpm_events[8] = mhpmevent_branch_i;
	// Trace: design.sv:9480:3
	assign hpm_events[9] = mhpmevent_branch_taken_i;
	// Trace: design.sv:9481:3
	assign hpm_events[10] = mhpmevent_compressed_i;
	// Trace: design.sv:9482:3
	assign hpm_events[11] = (PULP_CLUSTER ? mhpmevent_pipe_stall_i : 1'b0);
	// Trace: design.sv:9483:3
	assign hpm_events[12] = (!APU ? 1'b0 : apu_typeconflict_i && !apu_dep_i);
	// Trace: design.sv:9484:3
	assign hpm_events[13] = (!APU ? 1'b0 : apu_contention_i);
	// Trace: design.sv:9485:3
	assign hpm_events[14] = (!APU ? 1'b0 : apu_dep_i && !apu_contention_i);
	// Trace: design.sv:9486:3
	assign hpm_events[15] = (!APU ? 1'b0 : apu_wb_i);
	// Trace: design.sv:9490:3
	wire mcounteren_we;
	// Trace: design.sv:9491:3
	wire mcountinhibit_we;
	// Trace: design.sv:9492:3
	wire mhpmevent_we;
	// Trace: design.sv:9494:3
	assign mcounteren_we = csr_we_int & (csr_addr_i == 12'h306);
	// Trace: design.sv:9495:3
	assign mcountinhibit_we = csr_we_int & (csr_addr_i == 12'h320);
	// Trace: design.sv:9496:3
	assign mhpmevent_we = csr_we_int & (((((((((((((((((((((((((((((csr_addr_i == 12'h323) || (csr_addr_i == 12'h324)) || (csr_addr_i == 12'h325)) || (csr_addr_i == 12'h326)) || (csr_addr_i == 12'h327)) || (csr_addr_i == 12'h328)) || (csr_addr_i == 12'h329)) || (csr_addr_i == 12'h32a)) || (csr_addr_i == 12'h32b)) || (csr_addr_i == 12'h32c)) || (csr_addr_i == 12'h32d)) || (csr_addr_i == 12'h32e)) || (csr_addr_i == 12'h32f)) || (csr_addr_i == 12'h330)) || (csr_addr_i == 12'h331)) || (csr_addr_i == 12'h332)) || (csr_addr_i == 12'h333)) || (csr_addr_i == 12'h334)) || (csr_addr_i == 12'h335)) || (csr_addr_i == 12'h336)) || (csr_addr_i == 12'h337)) || (csr_addr_i == 12'h338)) || (csr_addr_i == 12'h339)) || (csr_addr_i == 12'h33a)) || (csr_addr_i == 12'h33b)) || (csr_addr_i == 12'h33c)) || (csr_addr_i == 12'h33d)) || (csr_addr_i == 12'h33e)) || (csr_addr_i == 12'h33f));
	// Trace: design.sv:9528:3
	genvar _gv_incr_gidx_1;
	// Trace: design.sv:9529:3
	generate
		for (_gv_incr_gidx_1 = 0; _gv_incr_gidx_1 < 32; _gv_incr_gidx_1 = _gv_incr_gidx_1 + 1) begin : gen_mhpmcounter_increment
			localparam incr_gidx = _gv_incr_gidx_1;
			// Trace: design.sv:9531:7
			assign mhpmcounter_increment[incr_gidx * 64+:64] = mhpmcounter_q[incr_gidx * 64+:64] + 1;
		end
	endgenerate
	// Trace: design.sv:9537:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:9538:5
		mcounteren_n = mcounteren_q;
		// Trace: design.sv:9539:5
		mcountinhibit_n = mcountinhibit_q;
		// Trace: design.sv:9540:5
		mhpmevent_n = mhpmevent_q;
		// Trace: design.sv:9543:5
		if (PULP_SECURE && mcounteren_we)
			// Trace: design.sv:9543:39
			mcounteren_n = csr_wdata_int;
		if (mcountinhibit_we)
			// Trace: design.sv:9546:27
			mcountinhibit_n = csr_wdata_int;
		if (mhpmevent_we)
			// Trace: design.sv:9549:23
			mhpmevent_n[csr_addr_i[4:0] * 32+:32] = csr_wdata_int;
	end
	// Trace: design.sv:9552:3
	genvar _gv_wcnt_gidx_1;
	// Trace: design.sv:9553:3
	generate
		for (_gv_wcnt_gidx_1 = 0; _gv_wcnt_gidx_1 < 32; _gv_wcnt_gidx_1 = _gv_wcnt_gidx_1 + 1) begin : gen_mhpmcounter_write
			localparam wcnt_gidx = _gv_wcnt_gidx_1;
			// Trace: design.sv:9557:7
			assign mhpmcounter_write_lower[wcnt_gidx] = csr_we_int && (csr_addr_i == (12'hb00 + wcnt_gidx));
			// Trace: design.sv:9560:7
			assign mhpmcounter_write_upper[wcnt_gidx] = ((!mhpmcounter_write_lower[wcnt_gidx] && csr_we_int) && (csr_addr_i == (12'hb80 + wcnt_gidx))) && 1'd1;
			if (!PULP_PERF_COUNTERS) begin : gen_no_pulp_perf_counters
				if (wcnt_gidx == 0) begin : gen_mhpmcounter_mcycle
					// Trace: design.sv:9567:11
					assign mhpmcounter_write_increment[wcnt_gidx] = (!mhpmcounter_write_lower[wcnt_gidx] && !mhpmcounter_write_upper[wcnt_gidx]) && !mcountinhibit_q[wcnt_gidx];
				end
				else if (wcnt_gidx == 2) begin : gen_mhpmcounter_minstret
					// Trace: design.sv:9572:11
					assign mhpmcounter_write_increment[wcnt_gidx] = ((!mhpmcounter_write_lower[wcnt_gidx] && !mhpmcounter_write_upper[wcnt_gidx]) && !mcountinhibit_q[wcnt_gidx]) && hpm_events[1];
				end
				else if ((wcnt_gidx > 2) && (wcnt_gidx < (NUM_MHPMCOUNTERS + 3))) begin : gen_mhpmcounter
					// Trace: design.sv:9578:11
					assign mhpmcounter_write_increment[wcnt_gidx] = ((!mhpmcounter_write_lower[wcnt_gidx] && !mhpmcounter_write_upper[wcnt_gidx]) && !mcountinhibit_q[wcnt_gidx]) && |(hpm_events & mhpmevent_q[(wcnt_gidx * 32) + 15-:16]);
				end
				else begin : gen_mhpmcounter_not_implemented
					// Trace: design.sv:9583:11
					assign mhpmcounter_write_increment[wcnt_gidx] = 1'b0;
				end
			end
			else begin : gen_pulp_perf_counters
				// Trace: design.sv:9587:9
				assign mhpmcounter_write_increment[wcnt_gidx] = ((!mhpmcounter_write_lower[wcnt_gidx] && !mhpmcounter_write_upper[wcnt_gidx]) && !mcountinhibit_q[wcnt_gidx]) && |(hpm_events & mhpmevent_q[(wcnt_gidx * 32) + 15-:16]);
			end
		end
	endgenerate
	// Trace: design.sv:9598:3
	genvar _gv_cnt_gidx_1;
	// Trace: design.sv:9599:3
	generate
		for (_gv_cnt_gidx_1 = 0; _gv_cnt_gidx_1 < 32; _gv_cnt_gidx_1 = _gv_cnt_gidx_1 + 1) begin : gen_mhpmcounter
			localparam cnt_gidx = _gv_cnt_gidx_1;
			if ((cnt_gidx == 1) || (cnt_gidx >= (NUM_MHPMCOUNTERS + 3))) begin : gen_non_implemented
				// Trace: design.sv:9606:9
				always @(posedge clk)
					// Trace: design.sv:9606:34
					mhpmcounter_q[cnt_gidx * 64+:64] <= 'b0;
			end
			else begin : gen_implemented
				// Trace: design.sv:9608:9
				always @(posedge clk or negedge rst_n)
					if (!rst_n)
						// Trace: design.sv:9610:13
						mhpmcounter_q[cnt_gidx * 64+:64] <= 'b0;
					else begin
						// Trace: design.sv:9612:13
						// Trace: design.sv:9615:15
						if (mhpmcounter_write_lower[cnt_gidx])
							// Trace: design.sv:9616:17
							mhpmcounter_q[(cnt_gidx * 64) + 31-:32] <= csr_wdata_int;
						else if (mhpmcounter_write_upper[cnt_gidx])
							// Trace: design.sv:9618:17
							mhpmcounter_q[(cnt_gidx * 64) + 63-:32] <= csr_wdata_int;
						else if (mhpmcounter_write_increment[cnt_gidx])
							// Trace: design.sv:9620:17
							mhpmcounter_q[cnt_gidx * 64+:64] <= mhpmcounter_increment[cnt_gidx * 64+:64];
					end
			end
		end
	endgenerate
	// Trace: design.sv:9629:3
	genvar _gv_evt_gidx_1;
	// Trace: design.sv:9630:3
	generate
		for (_gv_evt_gidx_1 = 0; _gv_evt_gidx_1 < 32; _gv_evt_gidx_1 = _gv_evt_gidx_1 + 1) begin : gen_mhpmevent
			localparam evt_gidx = _gv_evt_gidx_1;
			if ((evt_gidx < 3) || (evt_gidx >= (NUM_MHPMCOUNTERS + 3))) begin : gen_non_implemented
				// Trace: design.sv:9634:9
				always @(posedge clk)
					// Trace: design.sv:9634:34
					mhpmevent_q[evt_gidx * 32+:32] <= 'b0;
			end
			else begin : gen_implemented
				if (1) begin : gen_tie_off
					// Trace: design.sv:9637:11
					always @(posedge clk)
						// Trace: design.sv:9637:36
						mhpmevent_q[(evt_gidx * 32) + 31-:16] <= 'b0;
				end
				// Trace: design.sv:9639:9
				always @(posedge clk or negedge rst_n)
					if (!rst_n)
						// Trace: design.sv:9640:23
						mhpmevent_q[(evt_gidx * 32) + 15-:16] <= 'b0;
					else
						// Trace: design.sv:9642:13
						mhpmevent_q[(evt_gidx * 32) + 15-:16] <= mhpmevent_n[(evt_gidx * 32) + 15-:16];
			end
		end
	endgenerate
	// Trace: design.sv:9648:3
	genvar _gv_en_gidx_1;
	// Trace: design.sv:9649:3
	generate
		for (_gv_en_gidx_1 = 0; _gv_en_gidx_1 < 32; _gv_en_gidx_1 = _gv_en_gidx_1 + 1) begin : gen_mcounteren
			localparam en_gidx = _gv_en_gidx_1;
			if (((PULP_SECURE == 0) || (en_gidx == 1)) || (en_gidx >= (NUM_MHPMCOUNTERS + 3))) begin : gen_non_implemented
				// Trace: design.sv:9655:9
				always @(posedge clk)
					// Trace: design.sv:9655:34
					mcounteren_q[en_gidx] <= 'b0;
			end
			else begin : gen_implemented
				// Trace: design.sv:9657:9
				always @(posedge clk or negedge rst_n)
					if (!rst_n)
						// Trace: design.sv:9658:23
						mcounteren_q[en_gidx] <= 'b0;
					else
						// Trace: design.sv:9659:16
						mcounteren_q[en_gidx] <= mcounteren_n[en_gidx];
			end
		end
	endgenerate
	// Trace: design.sv:9666:3
	genvar _gv_inh_gidx_1;
	// Trace: design.sv:9667:3
	generate
		for (_gv_inh_gidx_1 = 0; _gv_inh_gidx_1 < 32; _gv_inh_gidx_1 = _gv_inh_gidx_1 + 1) begin : gen_mcountinhibit
			localparam inh_gidx = _gv_inh_gidx_1;
			if ((inh_gidx == 1) || (inh_gidx >= (NUM_MHPMCOUNTERS + 3))) begin : gen_non_implemented
				// Trace: design.sv:9670:9
				always @(posedge clk)
					// Trace: design.sv:9670:34
					mcountinhibit_q[inh_gidx] <= 'b0;
			end
			else begin : gen_implemented
				// Trace: design.sv:9672:9
				always @(posedge clk or negedge rst_n)
					if (!rst_n)
						// Trace: design.sv:9673:23
						mcountinhibit_q[inh_gidx] <= 'b1;
					else
						// Trace: design.sv:9674:16
						mcountinhibit_q[inh_gidx] <= mcountinhibit_n[inh_gidx];
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_decoder (
	deassert_we_i,
	illegal_insn_o,
	ebrk_insn_o,
	mret_insn_o,
	uret_insn_o,
	dret_insn_o,
	mret_dec_o,
	uret_dec_o,
	dret_dec_o,
	ecall_insn_o,
	wfi_o,
	fencei_insn_o,
	rega_used_o,
	regb_used_o,
	regc_used_o,
	reg_fp_a_o,
	reg_fp_b_o,
	reg_fp_c_o,
	reg_fp_d_o,
	bmask_a_mux_o,
	bmask_b_mux_o,
	alu_bmask_a_mux_sel_o,
	alu_bmask_b_mux_sel_o,
	instr_rdata_i,
	illegal_c_insn_i,
	alu_en_o,
	alu_operator_o,
	alu_op_a_mux_sel_o,
	alu_op_b_mux_sel_o,
	alu_op_c_mux_sel_o,
	alu_vec_mode_o,
	scalar_replication_o,
	scalar_replication_c_o,
	imm_a_mux_sel_o,
	imm_b_mux_sel_o,
	regc_mux_o,
	is_clpx_o,
	is_subrot_o,
	mult_operator_o,
	mult_int_en_o,
	mult_dot_en_o,
	mult_imm_mux_o,
	mult_sel_subword_o,
	mult_signed_mode_o,
	mult_dot_signed_o,
	frm_i,
	fpu_dst_fmt_o,
	fpu_src_fmt_o,
	fpu_int_fmt_o,
	apu_en_o,
	apu_op_o,
	apu_lat_o,
	fp_rnd_mode_o,
	regfile_mem_we_o,
	regfile_alu_we_o,
	regfile_alu_we_dec_o,
	regfile_alu_waddr_sel_o,
	csr_access_o,
	csr_status_o,
	csr_op_o,
	current_priv_lvl_i,
	data_req_o,
	data_we_o,
	prepost_useincr_o,
	data_type_o,
	data_sign_extension_o,
	data_reg_offset_o,
	data_load_event_o,
	atop_o,
	hwlp_we_o,
	hwlp_target_mux_sel_o,
	hwlp_start_mux_sel_o,
	hwlp_cnt_mux_sel_o,
	debug_mode_i,
	debug_wfi_no_sleep_i,
	ctrl_transfer_insn_in_dec_o,
	ctrl_transfer_insn_in_id_o,
	ctrl_transfer_target_mux_sel_o,
	mcounteren_i
);
	reg _sv2v_0;
	// removed import cv32e40p_pkg::*;
	// removed import cv32e40p_apu_core_pkg::*;
	// removed import cv32e40p_fpu_pkg::*;
	// Trace: design.sv:9722:13
	parameter PULP_XPULP = 1;
	// Trace: design.sv:9723:13
	parameter PULP_CLUSTER = 0;
	// Trace: design.sv:9724:13
	parameter A_EXTENSION = 0;
	// Trace: design.sv:9725:13
	parameter FPU = 0;
	// Trace: design.sv:9726:13
	parameter PULP_ZFINX = 0;
	// Trace: design.sv:9727:13
	parameter PULP_SECURE = 0;
	// Trace: design.sv:9728:13
	parameter USE_PMP = 0;
	// Trace: design.sv:9729:13
	parameter APU_WOP_CPU = 6;
	// Trace: design.sv:9730:13
	parameter DEBUG_TRIGGER_EN = 1;
	// Trace: design.sv:9734:3
	input wire deassert_we_i;
	// Trace: design.sv:9736:3
	output reg illegal_insn_o;
	// Trace: design.sv:9737:3
	output reg ebrk_insn_o;
	// Trace: design.sv:9739:3
	output reg mret_insn_o;
	// Trace: design.sv:9740:3
	output reg uret_insn_o;
	// Trace: design.sv:9741:3
	output reg dret_insn_o;
	// Trace: design.sv:9743:3
	output reg mret_dec_o;
	// Trace: design.sv:9744:3
	output reg uret_dec_o;
	// Trace: design.sv:9745:3
	output reg dret_dec_o;
	// Trace: design.sv:9747:3
	output reg ecall_insn_o;
	// Trace: design.sv:9748:3
	output reg wfi_o;
	// Trace: design.sv:9750:3
	output reg fencei_insn_o;
	// Trace: design.sv:9752:3
	output reg rega_used_o;
	// Trace: design.sv:9753:3
	output reg regb_used_o;
	// Trace: design.sv:9754:3
	output reg regc_used_o;
	// Trace: design.sv:9756:3
	output reg reg_fp_a_o;
	// Trace: design.sv:9757:3
	output reg reg_fp_b_o;
	// Trace: design.sv:9758:3
	output reg reg_fp_c_o;
	// Trace: design.sv:9759:3
	output reg reg_fp_d_o;
	// Trace: design.sv:9761:3
	output reg [0:0] bmask_a_mux_o;
	// Trace: design.sv:9762:3
	output reg [1:0] bmask_b_mux_o;
	// Trace: design.sv:9763:3
	output reg alu_bmask_a_mux_sel_o;
	// Trace: design.sv:9764:3
	output reg alu_bmask_b_mux_sel_o;
	// Trace: design.sv:9767:3
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:9768:3
	input wire illegal_c_insn_i;
	// Trace: design.sv:9771:3
	output wire alu_en_o;
	// Trace: design.sv:9772:3
	localparam cv32e40p_pkg_ALU_OP_WIDTH = 7;
	// removed localparam type cv32e40p_pkg_alu_opcode_e
	output reg [6:0] alu_operator_o;
	// Trace: design.sv:9773:3
	output reg [2:0] alu_op_a_mux_sel_o;
	// Trace: design.sv:9774:3
	output reg [2:0] alu_op_b_mux_sel_o;
	// Trace: design.sv:9775:3
	output reg [1:0] alu_op_c_mux_sel_o;
	// Trace: design.sv:9776:3
	output reg [1:0] alu_vec_mode_o;
	// Trace: design.sv:9777:3
	output reg scalar_replication_o;
	// Trace: design.sv:9778:3
	output reg scalar_replication_c_o;
	// Trace: design.sv:9779:3
	output reg [0:0] imm_a_mux_sel_o;
	// Trace: design.sv:9780:3
	output reg [3:0] imm_b_mux_sel_o;
	// Trace: design.sv:9781:3
	output reg [1:0] regc_mux_o;
	// Trace: design.sv:9782:3
	output reg is_clpx_o;
	// Trace: design.sv:9783:3
	output reg is_subrot_o;
	// Trace: design.sv:9786:3
	localparam cv32e40p_pkg_MUL_OP_WIDTH = 3;
	// removed localparam type cv32e40p_pkg_mul_opcode_e
	output reg [2:0] mult_operator_o;
	// Trace: design.sv:9787:3
	output wire mult_int_en_o;
	// Trace: design.sv:9788:3
	output wire mult_dot_en_o;
	// Trace: design.sv:9789:3
	output reg [0:0] mult_imm_mux_o;
	// Trace: design.sv:9790:3
	output reg mult_sel_subword_o;
	// Trace: design.sv:9791:3
	output reg [1:0] mult_signed_mode_o;
	// Trace: design.sv:9792:3
	output reg [1:0] mult_dot_signed_o;
	// Trace: design.sv:9795:3
	localparam cv32e40p_pkg_C_RM = 3;
	input wire [2:0] frm_i;
	// Trace: design.sv:9797:3
	localparam [31:0] cv32e40p_fpu_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] cv32e40p_fpu_pkg_FP_FORMAT_BITS = 3;
	output reg [2:0] fpu_dst_fmt_o;
	// Trace: design.sv:9798:3
	output reg [2:0] fpu_src_fmt_o;
	// Trace: design.sv:9799:3
	localparam [31:0] cv32e40p_fpu_pkg_NUM_INT_FORMATS = 4;
	localparam [31:0] cv32e40p_fpu_pkg_INT_FORMAT_BITS = 2;
	output reg [1:0] fpu_int_fmt_o;
	// Trace: design.sv:9802:3
	output wire apu_en_o;
	// Trace: design.sv:9803:3
	output reg [APU_WOP_CPU - 1:0] apu_op_o;
	// Trace: design.sv:9804:3
	output reg [1:0] apu_lat_o;
	// Trace: design.sv:9805:3
	output reg [2:0] fp_rnd_mode_o;
	// Trace: design.sv:9808:3
	output wire regfile_mem_we_o;
	// Trace: design.sv:9809:3
	output wire regfile_alu_we_o;
	// Trace: design.sv:9810:3
	output wire regfile_alu_we_dec_o;
	// Trace: design.sv:9811:3
	output reg regfile_alu_waddr_sel_o;
	// Trace: design.sv:9814:3
	output reg csr_access_o;
	// Trace: design.sv:9815:3
	output reg csr_status_o;
	// Trace: design.sv:9816:3
	localparam cv32e40p_pkg_CSR_OP_WIDTH = 2;
	// removed localparam type cv32e40p_pkg_csr_opcode_e
	output wire [1:0] csr_op_o;
	// Trace: design.sv:9817:3
	// removed localparam type cv32e40p_pkg_PrivLvl_t
	input wire [1:0] current_priv_lvl_i;
	// Trace: design.sv:9820:3
	output wire data_req_o;
	// Trace: design.sv:9821:3
	output reg data_we_o;
	// Trace: design.sv:9822:3
	output reg prepost_useincr_o;
	// Trace: design.sv:9823:3
	output reg [1:0] data_type_o;
	// Trace: design.sv:9824:3
	output reg [1:0] data_sign_extension_o;
	// Trace: design.sv:9825:3
	output reg [1:0] data_reg_offset_o;
	// Trace: design.sv:9826:3
	output reg data_load_event_o;
	// Trace: design.sv:9829:3
	output reg [5:0] atop_o;
	// Trace: design.sv:9832:3
	output wire [2:0] hwlp_we_o;
	// Trace: design.sv:9833:3
	output reg hwlp_target_mux_sel_o;
	// Trace: design.sv:9834:3
	output reg hwlp_start_mux_sel_o;
	// Trace: design.sv:9835:3
	output reg hwlp_cnt_mux_sel_o;
	// Trace: design.sv:9837:3
	input wire debug_mode_i;
	// Trace: design.sv:9838:3
	input wire debug_wfi_no_sleep_i;
	// Trace: design.sv:9841:3
	output wire [1:0] ctrl_transfer_insn_in_dec_o;
	// Trace: design.sv:9842:3
	output wire [1:0] ctrl_transfer_insn_in_id_o;
	// Trace: design.sv:9843:3
	output reg [1:0] ctrl_transfer_target_mux_sel_o;
	// Trace: design.sv:9846:3
	input wire [31:0] mcounteren_i;
	// Trace: design.sv:9850:3
	reg regfile_mem_we;
	// Trace: design.sv:9851:3
	reg regfile_alu_we;
	// Trace: design.sv:9852:3
	reg data_req;
	// Trace: design.sv:9853:3
	reg [2:0] hwlp_we;
	// Trace: design.sv:9854:3
	reg csr_illegal;
	// Trace: design.sv:9855:3
	reg [1:0] ctrl_transfer_insn;
	// Trace: design.sv:9857:3
	reg [1:0] csr_op;
	// Trace: design.sv:9859:3
	reg alu_en;
	// Trace: design.sv:9860:3
	reg mult_int_en;
	// Trace: design.sv:9861:3
	reg mult_dot_en;
	// Trace: design.sv:9862:3
	reg apu_en;
	// Trace: design.sv:9865:3
	reg check_fprm;
	// Trace: design.sv:9867:3
	localparam [31:0] cv32e40p_fpu_pkg_OP_BITS = 4;
	reg [3:0] fpu_op;
	// Trace: design.sv:9868:3
	reg fpu_op_mod;
	// Trace: design.sv:9869:3
	reg fpu_vec_op;
	// Trace: design.sv:9871:3
	reg [1:0] fp_op_group;
	// Trace: design.sv:9883:3
	localparam cv32e40p_apu_core_pkg_PIPE_REG_ADDSUB = 1;
	localparam cv32e40p_apu_core_pkg_PIPE_REG_CAST = 1;
	localparam cv32e40p_apu_core_pkg_PIPE_REG_MAC = 2;
	localparam cv32e40p_apu_core_pkg_PIPE_REG_MULT = 1;
	// removed localparam type cv32e40p_fpu_pkg_operation_e
	// removed localparam type cv32e40p_fpu_pkg_fp_format_e
	// removed localparam type cv32e40p_fpu_pkg_int_format_e
	localparam cv32e40p_pkg_AMO_ADD = 5'b00000;
	localparam cv32e40p_pkg_AMO_AND = 5'b01100;
	localparam cv32e40p_pkg_AMO_LR = 5'b00010;
	localparam cv32e40p_pkg_AMO_MAX = 5'b10100;
	localparam cv32e40p_pkg_AMO_MAXU = 5'b11100;
	localparam cv32e40p_pkg_AMO_MIN = 5'b10000;
	localparam cv32e40p_pkg_AMO_MINU = 5'b11000;
	localparam cv32e40p_pkg_AMO_OR = 5'b01000;
	localparam cv32e40p_pkg_AMO_SC = 5'b00011;
	localparam cv32e40p_pkg_AMO_SWAP = 5'b00001;
	localparam cv32e40p_pkg_AMO_XOR = 5'b00100;
	localparam cv32e40p_pkg_BMASK_A_IMM = 1'b1;
	localparam cv32e40p_pkg_BMASK_A_REG = 1'b0;
	localparam cv32e40p_pkg_BMASK_A_S3 = 1'b1;
	localparam cv32e40p_pkg_BMASK_A_ZERO = 1'b0;
	localparam cv32e40p_pkg_BMASK_B_IMM = 1'b1;
	localparam cv32e40p_pkg_BMASK_B_ONE = 2'b11;
	localparam cv32e40p_pkg_BMASK_B_REG = 1'b0;
	localparam cv32e40p_pkg_BMASK_B_S2 = 2'b00;
	localparam cv32e40p_pkg_BMASK_B_S3 = 2'b01;
	localparam cv32e40p_pkg_BMASK_B_ZERO = 2'b10;
	localparam cv32e40p_pkg_BRANCH_COND = 2'b11;
	localparam cv32e40p_pkg_BRANCH_JAL = 2'b01;
	localparam cv32e40p_pkg_BRANCH_JALR = 2'b10;
	localparam cv32e40p_pkg_BRANCH_NONE = 2'b00;
	// removed localparam type cv32e40p_pkg_csr_num_e
	localparam [31:0] cv32e40p_pkg_C_LAT_CONV = 'd0;
	localparam [31:0] cv32e40p_pkg_C_LAT_FP16 = 'd0;
	localparam [31:0] cv32e40p_pkg_C_LAT_FP16ALT = 'd0;
	localparam [31:0] cv32e40p_pkg_C_LAT_FP32 = 'd0;
	localparam [31:0] cv32e40p_pkg_C_LAT_FP64 = 'd0;
	localparam [31:0] cv32e40p_pkg_C_LAT_FP8 = 'd0;
	localparam [31:0] cv32e40p_pkg_C_LAT_NONCOMP = 'd0;
	localparam [0:0] cv32e40p_pkg_C_RVD = 1'b0;
	localparam [0:0] cv32e40p_pkg_C_RVF = 1'b1;
	localparam [0:0] cv32e40p_pkg_C_XF16 = 1'b0;
	localparam [0:0] cv32e40p_pkg_C_XF16ALT = 1'b0;
	localparam [0:0] cv32e40p_pkg_C_XF8 = 1'b0;
	localparam [0:0] cv32e40p_pkg_C_XFVEC = 1'b0;
	localparam cv32e40p_pkg_IMMA_Z = 1'b0;
	localparam cv32e40p_pkg_IMMA_ZERO = 1'b1;
	localparam cv32e40p_pkg_IMMB_BI = 4'b1011;
	localparam cv32e40p_pkg_IMMB_CLIP = 4'b1001;
	localparam cv32e40p_pkg_IMMB_I = 4'b0000;
	localparam cv32e40p_pkg_IMMB_PCINCR = 4'b0011;
	localparam cv32e40p_pkg_IMMB_S = 4'b0001;
	localparam cv32e40p_pkg_IMMB_S2 = 4'b0100;
	localparam cv32e40p_pkg_IMMB_SHUF = 4'b1000;
	localparam cv32e40p_pkg_IMMB_U = 4'b0010;
	localparam cv32e40p_pkg_IMMB_VS = 4'b0110;
	localparam cv32e40p_pkg_IMMB_VU = 4'b0111;
	localparam cv32e40p_pkg_JT_COND = 2'b11;
	localparam cv32e40p_pkg_JT_JAL = 2'b01;
	localparam cv32e40p_pkg_JT_JALR = 2'b10;
	localparam cv32e40p_pkg_MIMM_S3 = 1'b1;
	localparam cv32e40p_pkg_MIMM_ZERO = 1'b0;
	localparam cv32e40p_pkg_OPCODE_AMO = 7'h2f;
	localparam cv32e40p_pkg_OPCODE_AUIPC = 7'h17;
	localparam cv32e40p_pkg_OPCODE_BRANCH = 7'h63;
	localparam cv32e40p_pkg_OPCODE_FENCE = 7'h0f;
	localparam cv32e40p_pkg_OPCODE_HWLOOP = 7'h7b;
	localparam cv32e40p_pkg_OPCODE_JAL = 7'h6f;
	localparam cv32e40p_pkg_OPCODE_JALR = 7'h67;
	localparam cv32e40p_pkg_OPCODE_LOAD = 7'h03;
	localparam cv32e40p_pkg_OPCODE_LOAD_FP = 7'h07;
	localparam cv32e40p_pkg_OPCODE_LOAD_POST = 7'h0b;
	localparam cv32e40p_pkg_OPCODE_LUI = 7'h37;
	localparam cv32e40p_pkg_OPCODE_OP = 7'h33;
	localparam cv32e40p_pkg_OPCODE_OPIMM = 7'h13;
	localparam cv32e40p_pkg_OPCODE_OP_FMADD = 7'h43;
	localparam cv32e40p_pkg_OPCODE_OP_FMSUB = 7'h47;
	localparam cv32e40p_pkg_OPCODE_OP_FNMADD = 7'h4f;
	localparam cv32e40p_pkg_OPCODE_OP_FNMSUB = 7'h4b;
	localparam cv32e40p_pkg_OPCODE_OP_FP = 7'h53;
	localparam cv32e40p_pkg_OPCODE_PULP_OP = 7'h5b;
	localparam cv32e40p_pkg_OPCODE_STORE = 7'h23;
	localparam cv32e40p_pkg_OPCODE_STORE_FP = 7'h27;
	localparam cv32e40p_pkg_OPCODE_STORE_POST = 7'h2b;
	localparam cv32e40p_pkg_OPCODE_SYSTEM = 7'h73;
	localparam cv32e40p_pkg_OPCODE_VECOP = 7'h57;
	localparam cv32e40p_pkg_OP_A_CURRPC = 3'b001;
	localparam cv32e40p_pkg_OP_A_IMM = 3'b010;
	localparam cv32e40p_pkg_OP_A_REGA_OR_FWD = 3'b000;
	localparam cv32e40p_pkg_OP_A_REGB_OR_FWD = 3'b011;
	localparam cv32e40p_pkg_OP_A_REGC_OR_FWD = 3'b100;
	localparam cv32e40p_pkg_OP_B_BMASK = 3'b100;
	localparam cv32e40p_pkg_OP_B_IMM = 3'b010;
	localparam cv32e40p_pkg_OP_B_REGA_OR_FWD = 3'b011;
	localparam cv32e40p_pkg_OP_B_REGB_OR_FWD = 3'b000;
	localparam cv32e40p_pkg_OP_B_REGC_OR_FWD = 3'b001;
	localparam cv32e40p_pkg_OP_C_JT = 2'b10;
	localparam cv32e40p_pkg_OP_C_REGB_OR_FWD = 2'b01;
	localparam cv32e40p_pkg_OP_C_REGC_OR_FWD = 2'b00;
	localparam cv32e40p_pkg_REGC_RD = 2'b01;
	localparam cv32e40p_pkg_REGC_S4 = 2'b00;
	localparam cv32e40p_pkg_REGC_ZERO = 2'b11;
	localparam cv32e40p_pkg_VEC_MODE16 = 2'b10;
	localparam cv32e40p_pkg_VEC_MODE32 = 2'b00;
	localparam cv32e40p_pkg_VEC_MODE8 = 2'b11;
	function automatic [6:0] sv2v_cast_C07C4;
		input reg [6:0] inp;
		sv2v_cast_C07C4 = inp;
	endfunction
	function automatic [2:0] sv2v_cast_9F558;
		input reg [2:0] inp;
		sv2v_cast_9F558 = inp;
	endfunction
	function automatic [3:0] sv2v_cast_A1364;
		input reg [3:0] inp;
		sv2v_cast_A1364 = inp;
	endfunction
	function automatic [2:0] sv2v_cast_9D6B6;
		input reg [2:0] inp;
		sv2v_cast_9D6B6 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_1BCDC;
		input reg [1:0] inp;
		sv2v_cast_1BCDC = inp;
	endfunction
	function automatic [1:0] sv2v_cast_EB06E;
		input reg [1:0] inp;
		sv2v_cast_EB06E = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:9885:5
		ctrl_transfer_insn = cv32e40p_pkg_BRANCH_NONE;
		// Trace: design.sv:9886:5
		ctrl_transfer_target_mux_sel_o = cv32e40p_pkg_JT_JAL;
		// Trace: design.sv:9888:5
		alu_en = 1'b1;
		// Trace: design.sv:9889:5
		alu_operator_o = sv2v_cast_C07C4(7'b0000011);
		// Trace: design.sv:9890:5
		alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGA_OR_FWD;
		// Trace: design.sv:9891:5
		alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGB_OR_FWD;
		// Trace: design.sv:9892:5
		alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_REGC_OR_FWD;
		// Trace: design.sv:9893:5
		alu_vec_mode_o = cv32e40p_pkg_VEC_MODE32;
		// Trace: design.sv:9894:5
		scalar_replication_o = 1'b0;
		// Trace: design.sv:9895:5
		scalar_replication_c_o = 1'b0;
		// Trace: design.sv:9896:5
		regc_mux_o = cv32e40p_pkg_REGC_ZERO;
		// Trace: design.sv:9897:5
		imm_a_mux_sel_o = cv32e40p_pkg_IMMA_ZERO;
		// Trace: design.sv:9898:5
		imm_b_mux_sel_o = cv32e40p_pkg_IMMB_I;
		// Trace: design.sv:9900:5
		mult_operator_o = sv2v_cast_9F558(3'b010);
		// Trace: design.sv:9901:5
		mult_int_en = 1'b0;
		// Trace: design.sv:9902:5
		mult_dot_en = 1'b0;
		// Trace: design.sv:9903:5
		mult_imm_mux_o = cv32e40p_pkg_MIMM_ZERO;
		// Trace: design.sv:9904:5
		mult_signed_mode_o = 2'b00;
		// Trace: design.sv:9905:5
		mult_sel_subword_o = 1'b0;
		// Trace: design.sv:9906:5
		mult_dot_signed_o = 2'b00;
		// Trace: design.sv:9908:5
		apu_en = 1'b0;
		// Trace: design.sv:9909:5
		apu_op_o = 1'sb0;
		// Trace: design.sv:9910:5
		apu_lat_o = 1'sb0;
		// Trace: design.sv:9911:5
		fp_rnd_mode_o = 1'sb0;
		// Trace: design.sv:9912:5
		fpu_op = sv2v_cast_A1364(6);
		// Trace: design.sv:9913:5
		fpu_op_mod = 1'b0;
		// Trace: design.sv:9914:5
		fpu_vec_op = 1'b0;
		// Trace: design.sv:9915:5
		fpu_dst_fmt_o = sv2v_cast_9D6B6('d0);
		// Trace: design.sv:9916:5
		fpu_src_fmt_o = sv2v_cast_9D6B6('d0);
		// Trace: design.sv:9917:5
		fpu_int_fmt_o = sv2v_cast_1BCDC(2);
		// Trace: design.sv:9918:5
		check_fprm = 1'b0;
		// Trace: design.sv:9919:5
		fp_op_group = 2'd0;
		// Trace: design.sv:9921:5
		regfile_mem_we = 1'b0;
		// Trace: design.sv:9922:5
		regfile_alu_we = 1'b0;
		// Trace: design.sv:9923:5
		regfile_alu_waddr_sel_o = 1'b1;
		// Trace: design.sv:9925:5
		prepost_useincr_o = 1'b1;
		// Trace: design.sv:9927:5
		hwlp_we = 3'b000;
		// Trace: design.sv:9928:5
		hwlp_target_mux_sel_o = 1'b0;
		// Trace: design.sv:9929:5
		hwlp_start_mux_sel_o = 1'b0;
		// Trace: design.sv:9930:5
		hwlp_cnt_mux_sel_o = 1'b0;
		// Trace: design.sv:9932:5
		csr_access_o = 1'b0;
		// Trace: design.sv:9933:5
		csr_status_o = 1'b0;
		// Trace: design.sv:9934:5
		csr_illegal = 1'b0;
		// Trace: design.sv:9935:5
		csr_op = sv2v_cast_EB06E(2'b00);
		// Trace: design.sv:9936:5
		mret_insn_o = 1'b0;
		// Trace: design.sv:9937:5
		uret_insn_o = 1'b0;
		// Trace: design.sv:9939:5
		dret_insn_o = 1'b0;
		// Trace: design.sv:9941:5
		data_we_o = 1'b0;
		// Trace: design.sv:9942:5
		data_type_o = 2'b00;
		// Trace: design.sv:9943:5
		data_sign_extension_o = 2'b00;
		// Trace: design.sv:9944:5
		data_reg_offset_o = 2'b00;
		// Trace: design.sv:9945:5
		data_req = 1'b0;
		// Trace: design.sv:9946:5
		data_load_event_o = 1'b0;
		// Trace: design.sv:9948:5
		atop_o = 6'b000000;
		// Trace: design.sv:9950:5
		illegal_insn_o = 1'b0;
		// Trace: design.sv:9951:5
		ebrk_insn_o = 1'b0;
		// Trace: design.sv:9952:5
		ecall_insn_o = 1'b0;
		// Trace: design.sv:9953:5
		wfi_o = 1'b0;
		// Trace: design.sv:9955:5
		fencei_insn_o = 1'b0;
		// Trace: design.sv:9957:5
		rega_used_o = 1'b0;
		// Trace: design.sv:9958:5
		regb_used_o = 1'b0;
		// Trace: design.sv:9959:5
		regc_used_o = 1'b0;
		// Trace: design.sv:9960:5
		reg_fp_a_o = 1'b0;
		// Trace: design.sv:9961:5
		reg_fp_b_o = 1'b0;
		// Trace: design.sv:9962:5
		reg_fp_c_o = 1'b0;
		// Trace: design.sv:9963:5
		reg_fp_d_o = 1'b0;
		// Trace: design.sv:9965:5
		bmask_a_mux_o = cv32e40p_pkg_BMASK_A_ZERO;
		// Trace: design.sv:9966:5
		bmask_b_mux_o = cv32e40p_pkg_BMASK_B_ZERO;
		// Trace: design.sv:9967:5
		alu_bmask_a_mux_sel_o = cv32e40p_pkg_BMASK_A_IMM;
		// Trace: design.sv:9968:5
		alu_bmask_b_mux_sel_o = cv32e40p_pkg_BMASK_B_IMM;
		// Trace: design.sv:9970:5
		is_clpx_o = 1'b0;
		// Trace: design.sv:9971:5
		is_subrot_o = 1'b0;
		// Trace: design.sv:9973:5
		mret_dec_o = 1'b0;
		// Trace: design.sv:9974:5
		uret_dec_o = 1'b0;
		// Trace: design.sv:9975:5
		dret_dec_o = 1'b0;
		// Trace: design.sv:9977:5
		(* full_case, parallel_case *)
		case (instr_rdata_i[6:0])
			cv32e40p_pkg_OPCODE_JAL: begin
				// Trace: design.sv:9989:9
				ctrl_transfer_target_mux_sel_o = cv32e40p_pkg_JT_JAL;
				// Trace: design.sv:9990:9
				ctrl_transfer_insn = cv32e40p_pkg_BRANCH_JAL;
				// Trace: design.sv:9992:9
				alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_CURRPC;
				// Trace: design.sv:9993:9
				alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
				// Trace: design.sv:9994:9
				imm_b_mux_sel_o = cv32e40p_pkg_IMMB_PCINCR;
				// Trace: design.sv:9995:9
				alu_operator_o = sv2v_cast_C07C4(7'b0011000);
				// Trace: design.sv:9996:9
				regfile_alu_we = 1'b1;
			end
			cv32e40p_pkg_OPCODE_JALR: begin
				// Trace: design.sv:10001:9
				ctrl_transfer_target_mux_sel_o = cv32e40p_pkg_JT_JALR;
				// Trace: design.sv:10002:9
				ctrl_transfer_insn = cv32e40p_pkg_BRANCH_JALR;
				// Trace: design.sv:10004:9
				alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_CURRPC;
				// Trace: design.sv:10005:9
				alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
				// Trace: design.sv:10006:9
				imm_b_mux_sel_o = cv32e40p_pkg_IMMB_PCINCR;
				// Trace: design.sv:10007:9
				alu_operator_o = sv2v_cast_C07C4(7'b0011000);
				// Trace: design.sv:10008:9
				regfile_alu_we = 1'b1;
				// Trace: design.sv:10010:9
				rega_used_o = 1'b1;
				// Trace: design.sv:10012:9
				if (instr_rdata_i[14:12] != 3'b000) begin
					// Trace: design.sv:10013:11
					ctrl_transfer_insn = cv32e40p_pkg_BRANCH_NONE;
					// Trace: design.sv:10014:11
					regfile_alu_we = 1'b0;
					// Trace: design.sv:10015:11
					illegal_insn_o = 1'b1;
				end
			end
			cv32e40p_pkg_OPCODE_BRANCH: begin
				// Trace: design.sv:10020:9
				ctrl_transfer_target_mux_sel_o = cv32e40p_pkg_JT_COND;
				// Trace: design.sv:10021:9
				ctrl_transfer_insn = cv32e40p_pkg_BRANCH_COND;
				// Trace: design.sv:10022:9
				alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_JT;
				// Trace: design.sv:10023:9
				rega_used_o = 1'b1;
				// Trace: design.sv:10024:9
				regb_used_o = 1'b1;
				// Trace: design.sv:10026:9
				(* full_case, parallel_case *)
				case (instr_rdata_i[14:12])
					3'b000:
						// Trace: design.sv:10027:19
						alu_operator_o = sv2v_cast_C07C4(7'b0001100);
					3'b001:
						// Trace: design.sv:10028:19
						alu_operator_o = sv2v_cast_C07C4(7'b0001101);
					3'b100:
						// Trace: design.sv:10029:19
						alu_operator_o = sv2v_cast_C07C4(7'b0000000);
					3'b101:
						// Trace: design.sv:10030:19
						alu_operator_o = sv2v_cast_C07C4(7'b0001010);
					3'b110:
						// Trace: design.sv:10031:19
						alu_operator_o = sv2v_cast_C07C4(7'b0000001);
					3'b111:
						// Trace: design.sv:10032:19
						alu_operator_o = sv2v_cast_C07C4(7'b0001011);
					3'b010:
						// Trace: design.sv:10034:13
						if (PULP_XPULP) begin
							// Trace: design.sv:10035:15
							alu_operator_o = sv2v_cast_C07C4(7'b0001100);
							// Trace: design.sv:10036:15
							regb_used_o = 1'b0;
							// Trace: design.sv:10037:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
							// Trace: design.sv:10038:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_BI;
						end
						else
							// Trace: design.sv:10040:15
							illegal_insn_o = 1'b1;
					3'b011:
						// Trace: design.sv:10044:13
						if (PULP_XPULP) begin
							// Trace: design.sv:10045:15
							alu_operator_o = sv2v_cast_C07C4(7'b0001101);
							// Trace: design.sv:10046:15
							regb_used_o = 1'b0;
							// Trace: design.sv:10047:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
							// Trace: design.sv:10048:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_BI;
						end
						else
							// Trace: design.sv:10050:15
							illegal_insn_o = 1'b1;
				endcase
			end
			cv32e40p_pkg_OPCODE_STORE, cv32e40p_pkg_OPCODE_STORE_POST:
				// Trace: design.sv:10068:9
				if (PULP_XPULP || (instr_rdata_i[6:0] == cv32e40p_pkg_OPCODE_STORE)) begin
					// Trace: design.sv:10069:11
					data_req = 1'b1;
					// Trace: design.sv:10070:11
					data_we_o = 1'b1;
					// Trace: design.sv:10071:11
					rega_used_o = 1'b1;
					// Trace: design.sv:10072:11
					regb_used_o = 1'b1;
					// Trace: design.sv:10073:11
					alu_operator_o = sv2v_cast_C07C4(7'b0011000);
					// Trace: design.sv:10075:11
					alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_REGB_OR_FWD;
					// Trace: design.sv:10078:11
					if (instr_rdata_i[6:0] == cv32e40p_pkg_OPCODE_STORE_POST) begin
						// Trace: design.sv:10079:13
						prepost_useincr_o = 1'b0;
						// Trace: design.sv:10080:13
						regfile_alu_waddr_sel_o = 1'b0;
						// Trace: design.sv:10081:13
						regfile_alu_we = 1'b1;
					end
					if (instr_rdata_i[14] == 1'b0) begin
						// Trace: design.sv:10086:13
						imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S;
						// Trace: design.sv:10087:13
						alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
					end
					else
						// Trace: design.sv:10089:13
						if (PULP_XPULP) begin
							// Trace: design.sv:10091:15
							regc_used_o = 1'b1;
							// Trace: design.sv:10092:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGC_OR_FWD;
							// Trace: design.sv:10093:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
						end
						else
							// Trace: design.sv:10095:15
							illegal_insn_o = 1'b1;
					(* full_case, parallel_case *)
					case (instr_rdata_i[13:12])
						2'b00:
							// Trace: design.sv:10101:20
							data_type_o = 2'b10;
						2'b01:
							// Trace: design.sv:10102:20
							data_type_o = 2'b01;
						2'b10:
							// Trace: design.sv:10103:20
							data_type_o = 2'b00;
						default: begin
							// Trace: design.sv:10105:15
							data_req = 1'b0;
							// Trace: design.sv:10106:15
							data_we_o = 1'b0;
							// Trace: design.sv:10107:15
							illegal_insn_o = 1'b1;
						end
					endcase
				end
				else
					// Trace: design.sv:10111:11
					illegal_insn_o = 1'b1;
			cv32e40p_pkg_OPCODE_LOAD, cv32e40p_pkg_OPCODE_LOAD_POST:
				// Trace: design.sv:10117:9
				if (PULP_XPULP || (instr_rdata_i[6:0] == cv32e40p_pkg_OPCODE_LOAD)) begin
					// Trace: design.sv:10118:11
					data_req = 1'b1;
					// Trace: design.sv:10119:11
					regfile_mem_we = 1'b1;
					// Trace: design.sv:10120:11
					rega_used_o = 1'b1;
					// Trace: design.sv:10121:11
					data_type_o = 2'b00;
					// Trace: design.sv:10123:11
					alu_operator_o = sv2v_cast_C07C4(7'b0011000);
					// Trace: design.sv:10124:11
					alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
					// Trace: design.sv:10125:11
					imm_b_mux_sel_o = cv32e40p_pkg_IMMB_I;
					// Trace: design.sv:10128:11
					if (instr_rdata_i[6:0] == cv32e40p_pkg_OPCODE_LOAD_POST) begin
						// Trace: design.sv:10129:13
						prepost_useincr_o = 1'b0;
						// Trace: design.sv:10130:13
						regfile_alu_waddr_sel_o = 1'b0;
						// Trace: design.sv:10131:13
						regfile_alu_we = 1'b1;
					end
					// Trace: design.sv:10135:11
					data_sign_extension_o = {1'b0, ~instr_rdata_i[14]};
					(* full_case, parallel_case *)
					case (instr_rdata_i[13:12])
						2'b00:
							// Trace: design.sv:10139:22
							data_type_o = 2'b10;
						2'b01:
							// Trace: design.sv:10140:22
							data_type_o = 2'b01;
						2'b10:
							// Trace: design.sv:10141:22
							data_type_o = 2'b00;
						default:
							// Trace: design.sv:10142:22
							data_type_o = 2'b00;
					endcase
					if (instr_rdata_i[14:12] == 3'b111) begin
						begin
							// Trace: design.sv:10147:13
							if (PULP_XPULP) begin
								// Trace: design.sv:10149:15
								regb_used_o = 1'b1;
								// Trace: design.sv:10150:15
								alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGB_OR_FWD;
								// Trace: design.sv:10153:15
								data_sign_extension_o = {1'b0, ~instr_rdata_i[30]};
								// Trace: design.sv:10156:15
								(* full_case, parallel_case *)
								case (instr_rdata_i[31:25])
									7'b0000000, 7'b0100000:
										// Trace: design.sv:10158:30
										data_type_o = 2'b10;
									7'b0001000, 7'b0101000:
										// Trace: design.sv:10160:30
										data_type_o = 2'b01;
									7'b0010000:
										// Trace: design.sv:10161:30
										data_type_o = 2'b00;
									default:
										// Trace: design.sv:10163:19
										illegal_insn_o = 1'b1;
								endcase
							end
							else
								// Trace: design.sv:10167:15
								illegal_insn_o = 1'b1;
						end
					end
					if (instr_rdata_i[14:12] == 3'b110) begin
						begin
							// Trace: design.sv:10173:13
							if (PULP_CLUSTER && (instr_rdata_i[6:0] == cv32e40p_pkg_OPCODE_LOAD))
								// Trace: design.sv:10174:15
								data_load_event_o = 1'b1;
							else
								// Trace: design.sv:10177:15
								illegal_insn_o = 1'b1;
						end
					end
					if (instr_rdata_i[14:12] == 3'b011)
						// Trace: design.sv:10183:13
						illegal_insn_o = 1'b1;
				end
				else
					// Trace: design.sv:10186:11
					illegal_insn_o = 1'b1;
			cv32e40p_pkg_OPCODE_AMO:
				// Trace: design.sv:10191:9
				if (A_EXTENSION) begin : decode_amo
					// Trace: design.sv:10192:11
					if (instr_rdata_i[14:12] == 3'b010) begin
						// Trace: design.sv:10193:13
						data_req = 1'b1;
						// Trace: design.sv:10194:13
						data_type_o = 2'b00;
						// Trace: design.sv:10195:13
						rega_used_o = 1'b1;
						// Trace: design.sv:10196:13
						regb_used_o = 1'b1;
						// Trace: design.sv:10197:13
						regfile_mem_we = 1'b1;
						// Trace: design.sv:10198:13
						prepost_useincr_o = 1'b0;
						// Trace: design.sv:10199:13
						alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGA_OR_FWD;
						// Trace: design.sv:10201:13
						data_sign_extension_o = 1'b1;
						// Trace: design.sv:10204:13
						atop_o = {1'b1, instr_rdata_i[31:27]};
						// Trace: design.sv:10206:13
						(* full_case, parallel_case *)
						case (instr_rdata_i[31:27])
							cv32e40p_pkg_AMO_LR:
								// Trace: design.sv:10208:17
								data_we_o = 1'b0;
							cv32e40p_pkg_AMO_SC, cv32e40p_pkg_AMO_SWAP, cv32e40p_pkg_AMO_ADD, cv32e40p_pkg_AMO_XOR, cv32e40p_pkg_AMO_AND, cv32e40p_pkg_AMO_OR, cv32e40p_pkg_AMO_MIN, cv32e40p_pkg_AMO_MAX, cv32e40p_pkg_AMO_MINU, cv32e40p_pkg_AMO_MAXU: begin
								// Trace: design.sv:10220:17
								data_we_o = 1'b1;
								// Trace: design.sv:10221:17
								alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_REGB_OR_FWD;
							end
							default:
								// Trace: design.sv:10223:25
								illegal_insn_o = 1'b1;
						endcase
					end
					else
						// Trace: design.sv:10227:13
						illegal_insn_o = 1'b1;
				end
				else begin : no_decode_amo
					// Trace: design.sv:10230:11
					illegal_insn_o = 1'b1;
				end
			cv32e40p_pkg_OPCODE_LUI: begin
				// Trace: design.sv:10245:9
				alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_IMM;
				// Trace: design.sv:10246:9
				alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
				// Trace: design.sv:10247:9
				imm_a_mux_sel_o = cv32e40p_pkg_IMMA_ZERO;
				// Trace: design.sv:10248:9
				imm_b_mux_sel_o = cv32e40p_pkg_IMMB_U;
				// Trace: design.sv:10249:9
				alu_operator_o = sv2v_cast_C07C4(7'b0011000);
				// Trace: design.sv:10250:9
				regfile_alu_we = 1'b1;
			end
			cv32e40p_pkg_OPCODE_AUIPC: begin
				// Trace: design.sv:10254:9
				alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_CURRPC;
				// Trace: design.sv:10255:9
				alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
				// Trace: design.sv:10256:9
				imm_b_mux_sel_o = cv32e40p_pkg_IMMB_U;
				// Trace: design.sv:10257:9
				alu_operator_o = sv2v_cast_C07C4(7'b0011000);
				// Trace: design.sv:10258:9
				regfile_alu_we = 1'b1;
			end
			cv32e40p_pkg_OPCODE_OPIMM: begin
				// Trace: design.sv:10262:9
				alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
				// Trace: design.sv:10263:9
				imm_b_mux_sel_o = cv32e40p_pkg_IMMB_I;
				// Trace: design.sv:10264:9
				regfile_alu_we = 1'b1;
				// Trace: design.sv:10265:9
				rega_used_o = 1'b1;
				// Trace: design.sv:10267:9
				(* full_case, parallel_case *)
				case (instr_rdata_i[14:12])
					3'b000:
						// Trace: design.sv:10268:19
						alu_operator_o = sv2v_cast_C07C4(7'b0011000);
					3'b010:
						// Trace: design.sv:10269:19
						alu_operator_o = sv2v_cast_C07C4(7'b0000010);
					3'b011:
						// Trace: design.sv:10270:19
						alu_operator_o = sv2v_cast_C07C4(7'b0000011);
					3'b100:
						// Trace: design.sv:10271:19
						alu_operator_o = sv2v_cast_C07C4(7'b0101111);
					3'b110:
						// Trace: design.sv:10272:19
						alu_operator_o = sv2v_cast_C07C4(7'b0101110);
					3'b111:
						// Trace: design.sv:10273:19
						alu_operator_o = sv2v_cast_C07C4(7'b0010101);
					3'b001: begin
						// Trace: design.sv:10276:13
						alu_operator_o = sv2v_cast_C07C4(7'b0100111);
						// Trace: design.sv:10277:13
						if (instr_rdata_i[31:25] != 7'b0000000)
							// Trace: design.sv:10278:15
							illegal_insn_o = 1'b1;
					end
					3'b101:
						// Trace: design.sv:10282:13
						if (instr_rdata_i[31:25] == 7'b0000000)
							// Trace: design.sv:10283:15
							alu_operator_o = sv2v_cast_C07C4(7'b0100101);
						else if (instr_rdata_i[31:25] == 7'b0100000)
							// Trace: design.sv:10285:15
							alu_operator_o = sv2v_cast_C07C4(7'b0100100);
						else
							// Trace: design.sv:10287:15
							illegal_insn_o = 1'b1;
				endcase
			end
			cv32e40p_pkg_OPCODE_OP:
				// Trace: design.sv:10297:9
				if (instr_rdata_i[31:30] == 2'b11) begin
					begin
						// Trace: design.sv:10298:11
						if (PULP_XPULP) begin
							// Trace: design.sv:10303:13
							regfile_alu_we = 1'b1;
							// Trace: design.sv:10304:13
							rega_used_o = 1'b1;
							// Trace: design.sv:10307:13
							bmask_a_mux_o = cv32e40p_pkg_BMASK_A_S3;
							// Trace: design.sv:10308:13
							bmask_b_mux_o = cv32e40p_pkg_BMASK_B_S2;
							// Trace: design.sv:10309:13
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
							// Trace: design.sv:10311:13
							(* full_case, parallel_case *)
							case (instr_rdata_i[14:12])
								3'b000: begin
									// Trace: design.sv:10313:17
									alu_operator_o = sv2v_cast_C07C4(7'b0101000);
									// Trace: design.sv:10314:17
									imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S2;
									// Trace: design.sv:10315:17
									bmask_b_mux_o = cv32e40p_pkg_BMASK_B_ZERO;
								end
								3'b001: begin
									// Trace: design.sv:10318:17
									alu_operator_o = sv2v_cast_C07C4(7'b0101001);
									// Trace: design.sv:10319:17
									imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S2;
									// Trace: design.sv:10320:17
									bmask_b_mux_o = cv32e40p_pkg_BMASK_B_ZERO;
								end
								3'b010: begin
									// Trace: design.sv:10323:17
									alu_operator_o = sv2v_cast_C07C4(7'b0101010);
									// Trace: design.sv:10324:17
									imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S2;
									// Trace: design.sv:10325:17
									regc_used_o = 1'b1;
									// Trace: design.sv:10326:17
									regc_mux_o = cv32e40p_pkg_REGC_RD;
								end
								3'b011:
									// Trace: design.sv:10329:17
									alu_operator_o = sv2v_cast_C07C4(7'b0101011);
								3'b100:
									// Trace: design.sv:10332:17
									alu_operator_o = sv2v_cast_C07C4(7'b0101100);
								3'b101: begin
									// Trace: design.sv:10335:17
									alu_operator_o = sv2v_cast_C07C4(7'b1001001);
									// Trace: design.sv:10337:17
									regc_used_o = 1'b1;
									// Trace: design.sv:10338:17
									regc_mux_o = cv32e40p_pkg_REGC_RD;
									// Trace: design.sv:10340:17
									imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S2;
									// Trace: design.sv:10342:17
									alu_bmask_a_mux_sel_o = cv32e40p_pkg_BMASK_A_IMM;
									// Trace: design.sv:10343:17
									if (instr_rdata_i[29:27] != 3'b000)
										// Trace: design.sv:10344:19
										illegal_insn_o = 1'b1;
								end
								default:
									// Trace: design.sv:10347:24
									illegal_insn_o = 1'b1;
							endcase
						end
						else
							// Trace: design.sv:10350:13
							illegal_insn_o = 1'b1;
					end
				end
				else if (instr_rdata_i[31:30] == 2'b10) begin
					begin
						// Trace: design.sv:10359:11
						if (instr_rdata_i[29:25] == 5'b00000) begin
							begin
								// Trace: design.sv:10360:13
								if (PULP_XPULP) begin
									// Trace: design.sv:10361:15
									regfile_alu_we = 1'b1;
									// Trace: design.sv:10362:15
									rega_used_o = 1'b1;
									// Trace: design.sv:10364:15
									bmask_a_mux_o = cv32e40p_pkg_BMASK_A_S3;
									// Trace: design.sv:10365:15
									bmask_b_mux_o = cv32e40p_pkg_BMASK_B_S2;
									// Trace: design.sv:10366:15
									alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
									// Trace: design.sv:10368:15
									(* full_case, parallel_case *)
									case (instr_rdata_i[14:12])
										3'b000: begin
											// Trace: design.sv:10370:19
											alu_operator_o = sv2v_cast_C07C4(7'b0101000);
											// Trace: design.sv:10371:19
											imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S2;
											// Trace: design.sv:10372:19
											bmask_b_mux_o = cv32e40p_pkg_BMASK_B_ZERO;
											// Trace: design.sv:10374:19
											alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_BMASK;
											// Trace: design.sv:10375:19
											alu_bmask_a_mux_sel_o = cv32e40p_pkg_BMASK_A_REG;
											// Trace: design.sv:10376:19
											regb_used_o = 1'b1;
										end
										3'b001: begin
											// Trace: design.sv:10379:19
											alu_operator_o = sv2v_cast_C07C4(7'b0101001);
											// Trace: design.sv:10380:19
											imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S2;
											// Trace: design.sv:10381:19
											bmask_b_mux_o = cv32e40p_pkg_BMASK_B_ZERO;
											// Trace: design.sv:10383:19
											alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_BMASK;
											// Trace: design.sv:10384:19
											alu_bmask_a_mux_sel_o = cv32e40p_pkg_BMASK_A_REG;
											// Trace: design.sv:10385:19
											regb_used_o = 1'b1;
										end
										3'b010: begin
											// Trace: design.sv:10388:19
											alu_operator_o = sv2v_cast_C07C4(7'b0101010);
											// Trace: design.sv:10389:19
											imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S2;
											// Trace: design.sv:10390:19
											regc_used_o = 1'b1;
											// Trace: design.sv:10391:19
											regc_mux_o = cv32e40p_pkg_REGC_RD;
											// Trace: design.sv:10393:19
											alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_BMASK;
											// Trace: design.sv:10394:19
											alu_bmask_a_mux_sel_o = cv32e40p_pkg_BMASK_A_REG;
											// Trace: design.sv:10395:19
											alu_bmask_b_mux_sel_o = cv32e40p_pkg_BMASK_B_REG;
											// Trace: design.sv:10396:19
											regb_used_o = 1'b1;
										end
										3'b011: begin
											// Trace: design.sv:10399:19
											alu_operator_o = sv2v_cast_C07C4(7'b0101011);
											// Trace: design.sv:10401:19
											regb_used_o = 1'b1;
											// Trace: design.sv:10402:19
											alu_bmask_a_mux_sel_o = cv32e40p_pkg_BMASK_A_REG;
											// Trace: design.sv:10403:19
											alu_bmask_b_mux_sel_o = cv32e40p_pkg_BMASK_B_REG;
										end
										3'b100: begin
											// Trace: design.sv:10406:19
											alu_operator_o = sv2v_cast_C07C4(7'b0101100);
											// Trace: design.sv:10408:19
											regb_used_o = 1'b1;
											// Trace: design.sv:10409:19
											alu_bmask_a_mux_sel_o = cv32e40p_pkg_BMASK_A_REG;
											// Trace: design.sv:10410:19
											alu_bmask_b_mux_sel_o = cv32e40p_pkg_BMASK_B_REG;
										end
										default:
											// Trace: design.sv:10412:26
											illegal_insn_o = 1'b1;
									endcase
								end
								else
									// Trace: design.sv:10415:15
									illegal_insn_o = 1'b1;
							end
						end
						else
							// Trace: design.sv:10423:13
							if ((FPU == 1) && cv32e40p_pkg_C_XFVEC) begin
								// Trace: design.sv:10426:15
								apu_en = 1'b1;
								// Trace: design.sv:10427:15
								alu_en = 1'b0;
								// Trace: design.sv:10429:15
								rega_used_o = 1'b1;
								// Trace: design.sv:10430:15
								regb_used_o = 1'b1;
								// Trace: design.sv:10431:15
								if (PULP_ZFINX == 0) begin
									// Trace: design.sv:10432:17
									reg_fp_a_o = 1'b1;
									// Trace: design.sv:10433:17
									reg_fp_b_o = 1'b1;
									// Trace: design.sv:10434:17
									reg_fp_d_o = 1'b1;
								end
								else begin
									// Trace: design.sv:10436:17
									reg_fp_a_o = 1'b0;
									// Trace: design.sv:10437:17
									reg_fp_b_o = 1'b0;
									// Trace: design.sv:10438:17
									reg_fp_d_o = 1'b0;
								end
								// Trace: design.sv:10440:15
								fpu_vec_op = 1'b1;
								// Trace: design.sv:10442:15
								scalar_replication_o = instr_rdata_i[14];
								// Trace: design.sv:10444:15
								check_fprm = 1'b1;
								// Trace: design.sv:10445:15
								fp_rnd_mode_o = frm_i;
								(* full_case, parallel_case *)
								case (instr_rdata_i[13:12])
									2'b00: begin
										// Trace: design.sv:10451:19
										fpu_dst_fmt_o = sv2v_cast_9D6B6('d0);
										// Trace: design.sv:10452:19
										alu_vec_mode_o = cv32e40p_pkg_VEC_MODE32;
									end
									2'b01: begin
										// Trace: design.sv:10456:19
										fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
										// Trace: design.sv:10457:19
										alu_vec_mode_o = cv32e40p_pkg_VEC_MODE16;
									end
									2'b10: begin
										// Trace: design.sv:10461:19
										fpu_dst_fmt_o = sv2v_cast_9D6B6('d2);
										// Trace: design.sv:10462:19
										alu_vec_mode_o = cv32e40p_pkg_VEC_MODE16;
									end
									2'b11: begin
										// Trace: design.sv:10466:19
										fpu_dst_fmt_o = sv2v_cast_9D6B6('d3);
										// Trace: design.sv:10467:19
										alu_vec_mode_o = cv32e40p_pkg_VEC_MODE8;
									end
								endcase
								// Trace: design.sv:10472:15
								fpu_src_fmt_o = fpu_dst_fmt_o;
								(* full_case, parallel_case *)
								if (instr_rdata_i[29:25] == 5'b00001) begin
									// Trace: design.sv:10478:19
									fpu_op = sv2v_cast_A1364(2);
									// Trace: design.sv:10479:19
									fp_op_group = 2'd0;
									// Trace: design.sv:10481:19
									alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
									// Trace: design.sv:10482:19
									alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_REGB_OR_FWD;
									// Trace: design.sv:10483:19
									scalar_replication_o = 1'b0;
									// Trace: design.sv:10484:19
									scalar_replication_c_o = instr_rdata_i[14];
								end
								else if (instr_rdata_i[29:25] == 5'b00010) begin
									// Trace: design.sv:10488:19
									fpu_op = sv2v_cast_A1364(2);
									// Trace: design.sv:10489:19
									fpu_op_mod = 1'b1;
									// Trace: design.sv:10490:19
									fp_op_group = 2'd0;
									// Trace: design.sv:10492:19
									alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
									// Trace: design.sv:10493:19
									alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_REGB_OR_FWD;
									// Trace: design.sv:10494:19
									scalar_replication_o = 1'b0;
									// Trace: design.sv:10495:19
									scalar_replication_c_o = instr_rdata_i[14];
								end
								else if (instr_rdata_i[29:25] == 5'b00011) begin
									// Trace: design.sv:10499:19
									fpu_op = sv2v_cast_A1364(3);
									// Trace: design.sv:10500:19
									fp_op_group = 2'd0;
								end
								else if (instr_rdata_i[29:25] == 5'b00100) begin
									// Trace: design.sv:10504:19
									fpu_op = sv2v_cast_A1364(4);
									// Trace: design.sv:10505:19
									fp_op_group = 2'd1;
								end
								else if (instr_rdata_i[29:25] == 5'b00101) begin
									// Trace: design.sv:10509:19
									fpu_op = sv2v_cast_A1364(7);
									// Trace: design.sv:10510:19
									fp_rnd_mode_o = 3'b000;
									// Trace: design.sv:10511:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10512:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b00110) begin
									// Trace: design.sv:10516:19
									fpu_op = sv2v_cast_A1364(7);
									// Trace: design.sv:10517:19
									fp_rnd_mode_o = 3'b001;
									// Trace: design.sv:10518:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10519:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b00111) begin
									// Trace: design.sv:10523:19
									regb_used_o = 1'b0;
									// Trace: design.sv:10524:19
									fpu_op = sv2v_cast_A1364(5);
									// Trace: design.sv:10525:19
									fp_op_group = 2'd1;
									// Trace: design.sv:10527:19
									if ((instr_rdata_i[24:20] != 5'b00000) || instr_rdata_i[14])
										// Trace: design.sv:10528:21
										illegal_insn_o = 1'b1;
								end
								else if (instr_rdata_i[29:25] == 5'b01000) begin
									// Trace: design.sv:10533:19
									regc_used_o = 1'b1;
									// Trace: design.sv:10534:19
									regc_mux_o = cv32e40p_pkg_REGC_RD;
									// Trace: design.sv:10535:19
									if (PULP_ZFINX == 0)
										// Trace: design.sv:10536:21
										reg_fp_c_o = 1'b1;
									else
										// Trace: design.sv:10538:21
										reg_fp_c_o = 1'b0;
									// Trace: design.sv:10540:19
									fpu_op = sv2v_cast_A1364(0);
									// Trace: design.sv:10541:19
									fp_op_group = 2'd0;
								end
								else if (instr_rdata_i[29:25] == 5'b01001) begin
									// Trace: design.sv:10545:19
									regc_used_o = 1'b1;
									// Trace: design.sv:10546:19
									regc_mux_o = cv32e40p_pkg_REGC_RD;
									// Trace: design.sv:10547:19
									if (PULP_ZFINX == 0)
										// Trace: design.sv:10548:21
										reg_fp_c_o = 1'b1;
									else
										// Trace: design.sv:10550:21
										reg_fp_c_o = 1'b0;
									// Trace: design.sv:10552:19
									fpu_op = sv2v_cast_A1364(0);
									// Trace: design.sv:10553:19
									fpu_op_mod = 1'b1;
									// Trace: design.sv:10554:19
									fp_op_group = 2'd0;
								end
								else if (instr_rdata_i[29:25] == 5'b01100) begin
									// Trace: design.sv:10558:19
									regb_used_o = 1'b0;
									// Trace: design.sv:10559:19
									scalar_replication_o = 1'b0;
									// Trace: design.sv:10561:19
									(* full_case, parallel_case *)
									if (instr_rdata_i[24:20] == 5'b00000) begin
										// Trace: design.sv:10564:23
										alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
										// Trace: design.sv:10565:23
										fpu_op = sv2v_cast_A1364(6);
										// Trace: design.sv:10566:23
										fp_rnd_mode_o = 3'b011;
										// Trace: design.sv:10567:23
										fp_op_group = 2'd2;
										// Trace: design.sv:10568:23
										check_fprm = 1'b0;
										// Trace: design.sv:10570:23
										if (instr_rdata_i[14]) begin
											// Trace: design.sv:10571:25
											reg_fp_a_o = 1'b0;
											// Trace: design.sv:10572:25
											fpu_op_mod = 1'b0;
										end
										else begin
											// Trace: design.sv:10576:25
											reg_fp_d_o = 1'b0;
											// Trace: design.sv:10577:25
											fpu_op_mod = 1'b1;
										end
									end
									else if (instr_rdata_i[24:20] == 5'b00001) begin
										// Trace: design.sv:10582:23
										reg_fp_d_o = 1'b0;
										// Trace: design.sv:10583:23
										fpu_op = sv2v_cast_A1364(9);
										// Trace: design.sv:10584:23
										fp_rnd_mode_o = 3'b000;
										// Trace: design.sv:10585:23
										fp_op_group = 2'd2;
										// Trace: design.sv:10586:23
										check_fprm = 1'b0;
										// Trace: design.sv:10588:23
										if (instr_rdata_i[14])
											// Trace: design.sv:10588:46
											illegal_insn_o = 1'b1;
									end
									else if ((instr_rdata_i[24:20] | 5'b00001) == 5'b00011) begin
										// Trace: design.sv:10592:23
										fp_op_group = 2'd3;
										// Trace: design.sv:10593:23
										fpu_op_mod = instr_rdata_i[14];
										// Trace: design.sv:10595:23
										(* full_case, parallel_case *)
										case (instr_rdata_i[13:12])
											2'b00:
												// Trace: design.sv:10597:33
												fpu_int_fmt_o = sv2v_cast_1BCDC(2);
											2'b01, 2'b10:
												// Trace: design.sv:10600:32
												fpu_int_fmt_o = sv2v_cast_1BCDC(1);
											2'b11:
												// Trace: design.sv:10602:32
												fpu_int_fmt_o = sv2v_cast_1BCDC(0);
										endcase
										if (instr_rdata_i[20]) begin
											// Trace: design.sv:10606:25
											reg_fp_a_o = 1'b0;
											// Trace: design.sv:10607:25
											fpu_op = sv2v_cast_A1364(12);
										end
										else begin
											// Trace: design.sv:10611:25
											reg_fp_d_o = 1'b0;
											// Trace: design.sv:10612:25
											fpu_op = sv2v_cast_A1364(11);
										end
									end
									else if ((instr_rdata_i[24:20] | 5'b00011) == 5'b00111) begin
										// Trace: design.sv:10617:23
										fpu_op = sv2v_cast_A1364(10);
										// Trace: design.sv:10618:23
										fp_op_group = 2'd3;
										// Trace: design.sv:10620:23
										(* full_case, parallel_case *)
										case (instr_rdata_i[21:20])
											2'b00: begin
												// Trace: design.sv:10623:27
												fpu_src_fmt_o = sv2v_cast_9D6B6('d0);
												// Trace: design.sv:10624:27
												if (~cv32e40p_pkg_C_RVF)
													// Trace: design.sv:10624:39
													illegal_insn_o = 1'b1;
											end
											2'b01: begin
												// Trace: design.sv:10627:27
												fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
												// Trace: design.sv:10628:27
												if (~cv32e40p_pkg_C_XF16ALT)
													// Trace: design.sv:10628:43
													illegal_insn_o = 1'b1;
											end
											2'b10: begin
												// Trace: design.sv:10631:27
												fpu_src_fmt_o = sv2v_cast_9D6B6('d2);
												// Trace: design.sv:10632:27
												if (~cv32e40p_pkg_C_XF16)
													// Trace: design.sv:10632:40
													illegal_insn_o = 1'b1;
											end
											2'b11: begin
												// Trace: design.sv:10635:27
												fpu_src_fmt_o = sv2v_cast_9D6B6('d3);
												// Trace: design.sv:10636:27
												if (~cv32e40p_pkg_C_XF8)
													// Trace: design.sv:10636:39
													illegal_insn_o = 1'b1;
											end
										endcase
										if (instr_rdata_i[14])
											// Trace: design.sv:10640:46
											illegal_insn_o = 1'b1;
									end
									else
										// Trace: design.sv:10643:31
										illegal_insn_o = 1'b1;
								end
								else if (instr_rdata_i[29:25] == 5'b01101) begin
									// Trace: design.sv:10648:19
									fpu_op = sv2v_cast_A1364(6);
									// Trace: design.sv:10649:19
									fp_rnd_mode_o = 3'b000;
									// Trace: design.sv:10650:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10651:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b01110) begin
									// Trace: design.sv:10655:19
									fpu_op = sv2v_cast_A1364(6);
									// Trace: design.sv:10656:19
									fp_rnd_mode_o = 3'b001;
									// Trace: design.sv:10657:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10658:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b01111) begin
									// Trace: design.sv:10662:19
									fpu_op = sv2v_cast_A1364(6);
									// Trace: design.sv:10663:19
									fp_rnd_mode_o = 3'b010;
									// Trace: design.sv:10664:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10665:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b10000) begin
									// Trace: design.sv:10669:19
									reg_fp_d_o = 1'b0;
									// Trace: design.sv:10670:19
									fpu_op = sv2v_cast_A1364(8);
									// Trace: design.sv:10671:19
									fp_rnd_mode_o = 3'b010;
									// Trace: design.sv:10672:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10673:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b10001) begin
									// Trace: design.sv:10677:19
									reg_fp_d_o = 1'b0;
									// Trace: design.sv:10678:19
									fpu_op = sv2v_cast_A1364(8);
									// Trace: design.sv:10679:19
									fpu_op_mod = 1'b1;
									// Trace: design.sv:10680:19
									fp_rnd_mode_o = 3'b010;
									// Trace: design.sv:10681:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10682:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b10010) begin
									// Trace: design.sv:10686:19
									reg_fp_d_o = 1'b0;
									// Trace: design.sv:10687:19
									fpu_op = sv2v_cast_A1364(8);
									// Trace: design.sv:10688:19
									fp_rnd_mode_o = 3'b001;
									// Trace: design.sv:10689:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10690:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b10011) begin
									// Trace: design.sv:10694:19
									reg_fp_d_o = 1'b0;
									// Trace: design.sv:10695:19
									fpu_op = sv2v_cast_A1364(8);
									// Trace: design.sv:10696:19
									fpu_op_mod = 1'b1;
									// Trace: design.sv:10697:19
									fp_rnd_mode_o = 3'b001;
									// Trace: design.sv:10698:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10699:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b10100) begin
									// Trace: design.sv:10703:19
									reg_fp_d_o = 1'b0;
									// Trace: design.sv:10704:19
									fpu_op = sv2v_cast_A1364(8);
									// Trace: design.sv:10705:19
									fp_rnd_mode_o = 3'b000;
									// Trace: design.sv:10706:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10707:19
									check_fprm = 1'b0;
								end
								else if (instr_rdata_i[29:25] == 5'b10101) begin
									// Trace: design.sv:10711:19
									reg_fp_d_o = 1'b0;
									// Trace: design.sv:10712:19
									fpu_op = sv2v_cast_A1364(8);
									// Trace: design.sv:10713:19
									fpu_op_mod = 1'b1;
									// Trace: design.sv:10714:19
									fp_rnd_mode_o = 3'b000;
									// Trace: design.sv:10715:19
									fp_op_group = 2'd2;
									// Trace: design.sv:10716:19
									check_fprm = 1'b0;
								end
								else if ((instr_rdata_i[29:25] | 5'b00011) == 5'b11011) begin
									// Trace: design.sv:10721:19
									fpu_op_mod = instr_rdata_i[14];
									// Trace: design.sv:10722:19
									fp_op_group = 2'd3;
									// Trace: design.sv:10723:19
									scalar_replication_o = 1'b0;
									// Trace: design.sv:10725:19
									if (instr_rdata_i[25])
										// Trace: design.sv:10725:42
										fpu_op = sv2v_cast_A1364(14);
									else
										// Trace: design.sv:10726:24
										fpu_op = sv2v_cast_A1364(13);
									if (instr_rdata_i[26]) begin
										// Trace: design.sv:10730:21
										fpu_src_fmt_o = sv2v_cast_9D6B6('d1);
										// Trace: design.sv:10731:21
										if (~cv32e40p_pkg_C_RVD)
											// Trace: design.sv:10731:33
											illegal_insn_o = 1'b1;
									end
									else begin
										// Trace: design.sv:10735:21
										fpu_src_fmt_o = sv2v_cast_9D6B6('d0);
										// Trace: design.sv:10736:21
										if (~cv32e40p_pkg_C_RVF)
											// Trace: design.sv:10736:33
											illegal_insn_o = 1'b1;
									end
									if (fpu_op == sv2v_cast_A1364(14)) begin
										begin
											// Trace: design.sv:10740:21
											if (~cv32e40p_pkg_C_XF8 || ~cv32e40p_pkg_C_RVD)
												// Trace: design.sv:10740:43
												illegal_insn_o = 1'b1;
										end
									end
									else
										// Trace: design.sv:10742:21
										if (instr_rdata_i[14]) begin
											// Trace: design.sv:10744:23
											if (fpu_dst_fmt_o == sv2v_cast_9D6B6('d0))
												// Trace: design.sv:10744:68
												illegal_insn_o = 1'b1;
											if (~cv32e40p_pkg_C_RVD && (fpu_dst_fmt_o != sv2v_cast_9D6B6('d3)))
												// Trace: design.sv:10746:79
												illegal_insn_o = 1'b1;
										end
								end
								else
									// Trace: design.sv:10752:19
									illegal_insn_o = 1'b1;
								if ((~cv32e40p_pkg_C_RVF || ~cv32e40p_pkg_C_RVD) && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d0)))
									// Trace: design.sv:10758:82
									illegal_insn_o = 1'b1;
								if ((~cv32e40p_pkg_C_XF16 || ~cv32e40p_pkg_C_RVF) && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d2)))
									// Trace: design.sv:10760:83
									illegal_insn_o = 1'b1;
								if ((~cv32e40p_pkg_C_XF16ALT || ~cv32e40p_pkg_C_RVF) && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d4)))
									// Trace: design.sv:10763:17
									illegal_insn_o = 1'b1;
								if ((~cv32e40p_pkg_C_XF8 || (~cv32e40p_pkg_C_XF16 && ~cv32e40p_pkg_C_XF16ALT)) && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d3)))
									// Trace: design.sv:10767:17
									illegal_insn_o = 1'b1;
								if (check_fprm) begin
									begin
										// Trace: design.sv:10772:17
										(* full_case, parallel_case *)
										if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
											;
										else
											// Trace: design.sv:10774:37
											illegal_insn_o = 1'b1;
									end
								end
								case (fp_op_group)
									2'd0:
										// Trace: design.sv:10784:19
										(* full_case, parallel_case *)
										case (fpu_dst_fmt_o)
											sv2v_cast_9D6B6('d0):
												// Trace: design.sv:10785:49
												apu_lat_o = 1;
											sv2v_cast_9D6B6('d2):
												// Trace: design.sv:10786:49
												apu_lat_o = 1;
											sv2v_cast_9D6B6('d4):
												// Trace: design.sv:10787:49
												apu_lat_o = 1;
											sv2v_cast_9D6B6('d3):
												// Trace: design.sv:10788:49
												apu_lat_o = 1;
											default:
												;
										endcase
									2'd1:
										// Trace: design.sv:10793:27
										apu_lat_o = 2'h3;
									2'd2:
										// Trace: design.sv:10795:27
										apu_lat_o = 1;
									2'd3:
										// Trace: design.sv:10797:27
										apu_lat_o = 1;
								endcase
								// Trace: design.sv:10801:15
								apu_op_o = {fpu_vec_op, fpu_op_mod, fpu_op};
							end
							else
								// Trace: design.sv:10805:15
								illegal_insn_o = 1'b1;
					end
				end
				else begin
					// Trace: design.sv:10814:11
					regfile_alu_we = 1'b1;
					// Trace: design.sv:10815:11
					rega_used_o = 1'b1;
					// Trace: design.sv:10817:11
					if (~instr_rdata_i[28])
						// Trace: design.sv:10817:35
						regb_used_o = 1'b1;
					(* full_case, parallel_case *)
					case ({instr_rdata_i[30:25], instr_rdata_i[14:12]})
						9'b000000000:
							// Trace: design.sv:10821:35
							alu_operator_o = sv2v_cast_C07C4(7'b0011000);
						9'b100000000:
							// Trace: design.sv:10822:35
							alu_operator_o = sv2v_cast_C07C4(7'b0011001);
						9'b000000010:
							// Trace: design.sv:10823:35
							alu_operator_o = sv2v_cast_C07C4(7'b0000010);
						9'b000000011:
							// Trace: design.sv:10824:35
							alu_operator_o = sv2v_cast_C07C4(7'b0000011);
						9'b000000100:
							// Trace: design.sv:10825:35
							alu_operator_o = sv2v_cast_C07C4(7'b0101111);
						9'b000000110:
							// Trace: design.sv:10826:35
							alu_operator_o = sv2v_cast_C07C4(7'b0101110);
						9'b000000111:
							// Trace: design.sv:10827:35
							alu_operator_o = sv2v_cast_C07C4(7'b0010101);
						9'b000000001:
							// Trace: design.sv:10828:35
							alu_operator_o = sv2v_cast_C07C4(7'b0100111);
						9'b000000101:
							// Trace: design.sv:10829:35
							alu_operator_o = sv2v_cast_C07C4(7'b0100101);
						9'b100000101:
							// Trace: design.sv:10830:35
							alu_operator_o = sv2v_cast_C07C4(7'b0100100);
						9'b000001000: begin
							// Trace: design.sv:10834:15
							alu_en = 1'b0;
							// Trace: design.sv:10835:15
							mult_int_en = 1'b1;
							// Trace: design.sv:10836:15
							mult_operator_o = sv2v_cast_9F558(3'b000);
							// Trace: design.sv:10837:15
							regc_mux_o = cv32e40p_pkg_REGC_ZERO;
						end
						9'b000001001: begin
							// Trace: design.sv:10840:15
							alu_en = 1'b0;
							// Trace: design.sv:10841:15
							regc_used_o = 1'b1;
							// Trace: design.sv:10842:15
							regc_mux_o = cv32e40p_pkg_REGC_ZERO;
							// Trace: design.sv:10843:15
							mult_signed_mode_o = 2'b11;
							// Trace: design.sv:10844:15
							mult_int_en = 1'b1;
							// Trace: design.sv:10845:15
							mult_operator_o = sv2v_cast_9F558(3'b110);
						end
						9'b000001010: begin
							// Trace: design.sv:10848:15
							alu_en = 1'b0;
							// Trace: design.sv:10849:15
							regc_used_o = 1'b1;
							// Trace: design.sv:10850:15
							regc_mux_o = cv32e40p_pkg_REGC_ZERO;
							// Trace: design.sv:10851:15
							mult_signed_mode_o = 2'b01;
							// Trace: design.sv:10852:15
							mult_int_en = 1'b1;
							// Trace: design.sv:10853:15
							mult_operator_o = sv2v_cast_9F558(3'b110);
						end
						9'b000001011: begin
							// Trace: design.sv:10856:15
							alu_en = 1'b0;
							// Trace: design.sv:10857:15
							regc_used_o = 1'b1;
							// Trace: design.sv:10858:15
							regc_mux_o = cv32e40p_pkg_REGC_ZERO;
							// Trace: design.sv:10859:15
							mult_signed_mode_o = 2'b00;
							// Trace: design.sv:10860:15
							mult_int_en = 1'b1;
							// Trace: design.sv:10861:15
							mult_operator_o = sv2v_cast_9F558(3'b110);
						end
						9'b000001100: begin
							// Trace: design.sv:10864:15
							alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGB_OR_FWD;
							// Trace: design.sv:10865:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
							// Trace: design.sv:10866:15
							regb_used_o = 1'b1;
							// Trace: design.sv:10867:15
							alu_operator_o = sv2v_cast_C07C4(7'b0110001);
						end
						9'b000001101: begin
							// Trace: design.sv:10870:15
							alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGB_OR_FWD;
							// Trace: design.sv:10871:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
							// Trace: design.sv:10872:15
							regb_used_o = 1'b1;
							// Trace: design.sv:10873:15
							alu_operator_o = sv2v_cast_C07C4(7'b0110000);
						end
						9'b000001110: begin
							// Trace: design.sv:10876:15
							alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGB_OR_FWD;
							// Trace: design.sv:10877:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
							// Trace: design.sv:10878:15
							regb_used_o = 1'b1;
							// Trace: design.sv:10879:15
							alu_operator_o = sv2v_cast_C07C4(7'b0110011);
						end
						9'b000001111: begin
							// Trace: design.sv:10882:15
							alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGB_OR_FWD;
							// Trace: design.sv:10883:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
							// Trace: design.sv:10884:15
							regb_used_o = 1'b1;
							// Trace: design.sv:10885:15
							alu_operator_o = sv2v_cast_C07C4(7'b0110010);
						end
						9'b100001000:
							// Trace: design.sv:10890:15
							if (PULP_XPULP) begin
								// Trace: design.sv:10891:17
								alu_en = 1'b0;
								// Trace: design.sv:10892:17
								regc_used_o = 1'b1;
								// Trace: design.sv:10893:17
								regc_mux_o = cv32e40p_pkg_REGC_RD;
								// Trace: design.sv:10894:17
								mult_int_en = 1'b1;
								// Trace: design.sv:10895:17
								mult_operator_o = sv2v_cast_9F558(3'b000);
							end
							else
								// Trace: design.sv:10897:17
								illegal_insn_o = 1'b1;
						9'b100001001:
							// Trace: design.sv:10901:15
							if (PULP_XPULP) begin
								// Trace: design.sv:10902:17
								alu_en = 1'b0;
								// Trace: design.sv:10903:17
								regc_used_o = 1'b1;
								// Trace: design.sv:10904:17
								regc_mux_o = cv32e40p_pkg_REGC_RD;
								// Trace: design.sv:10905:17
								mult_int_en = 1'b1;
								// Trace: design.sv:10906:17
								mult_operator_o = sv2v_cast_9F558(3'b001);
							end
							else
								// Trace: design.sv:10908:17
								illegal_insn_o = 1'b1;
						9'b000010010:
							// Trace: design.sv:10912:15
							if (PULP_XPULP)
								// Trace: design.sv:10913:17
								alu_operator_o = sv2v_cast_C07C4(7'b0000110);
							else
								// Trace: design.sv:10915:17
								illegal_insn_o = 1'b1;
						9'b000010011:
							// Trace: design.sv:10919:15
							if (PULP_XPULP)
								// Trace: design.sv:10920:17
								alu_operator_o = sv2v_cast_C07C4(7'b0000111);
							else
								// Trace: design.sv:10922:17
								illegal_insn_o = 1'b1;
						9'b000010100:
							// Trace: design.sv:10926:15
							if (PULP_XPULP)
								// Trace: design.sv:10927:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010000);
							else
								// Trace: design.sv:10929:17
								illegal_insn_o = 1'b1;
						9'b000010101:
							// Trace: design.sv:10933:15
							if (PULP_XPULP)
								// Trace: design.sv:10934:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010001);
							else
								// Trace: design.sv:10936:17
								illegal_insn_o = 1'b1;
						9'b000010110:
							// Trace: design.sv:10940:15
							if (PULP_XPULP)
								// Trace: design.sv:10941:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010010);
							else
								// Trace: design.sv:10943:17
								illegal_insn_o = 1'b1;
						9'b000010111:
							// Trace: design.sv:10947:15
							if (PULP_XPULP)
								// Trace: design.sv:10948:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010011);
							else
								// Trace: design.sv:10950:17
								illegal_insn_o = 1'b1;
						9'b000100101:
							// Trace: design.sv:10954:15
							if (PULP_XPULP)
								// Trace: design.sv:10955:17
								alu_operator_o = sv2v_cast_C07C4(7'b0100110);
							else
								// Trace: design.sv:10957:17
								illegal_insn_o = 1'b1;
						9'b001000000:
							// Trace: design.sv:10964:15
							if (PULP_XPULP) begin
								// Trace: design.sv:10965:17
								alu_operator_o = sv2v_cast_C07C4(7'b0110110);
								// Trace: design.sv:10966:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:10967:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:10970:17
								illegal_insn_o = 1'b1;
						9'b001000001:
							// Trace: design.sv:10974:15
							if (PULP_XPULP) begin
								// Trace: design.sv:10975:17
								alu_operator_o = sv2v_cast_C07C4(7'b0110111);
								// Trace: design.sv:10976:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:10977:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:10980:17
								illegal_insn_o = 1'b1;
						9'b001000010:
							// Trace: design.sv:10984:15
							if (PULP_XPULP) begin
								// Trace: design.sv:10985:17
								alu_operator_o = sv2v_cast_C07C4(7'b0110101);
								// Trace: design.sv:10986:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:10987:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:10990:17
								illegal_insn_o = 1'b1;
						9'b001000011:
							// Trace: design.sv:10994:15
							if (PULP_XPULP) begin
								// Trace: design.sv:10995:17
								alu_operator_o = sv2v_cast_C07C4(7'b0110100);
								// Trace: design.sv:10996:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:10997:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:11000:17
								illegal_insn_o = 1'b1;
						9'b001000100:
							// Trace: design.sv:11004:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11005:17
								alu_operator_o = sv2v_cast_C07C4(7'b0111110);
								// Trace: design.sv:11006:17
								alu_vec_mode_o = cv32e40p_pkg_VEC_MODE16;
								// Trace: design.sv:11007:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:11008:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:11011:17
								illegal_insn_o = 1'b1;
						9'b001000101:
							// Trace: design.sv:11015:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11016:17
								alu_operator_o = sv2v_cast_C07C4(7'b0111111);
								// Trace: design.sv:11017:17
								alu_vec_mode_o = cv32e40p_pkg_VEC_MODE16;
								// Trace: design.sv:11018:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:11019:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:11022:17
								illegal_insn_o = 1'b1;
						9'b001000110:
							// Trace: design.sv:11026:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11027:17
								alu_operator_o = sv2v_cast_C07C4(7'b0111110);
								// Trace: design.sv:11028:17
								alu_vec_mode_o = cv32e40p_pkg_VEC_MODE8;
								// Trace: design.sv:11029:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:11030:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:11033:17
								illegal_insn_o = 1'b1;
						9'b001000111:
							// Trace: design.sv:11037:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11038:17
								alu_operator_o = sv2v_cast_C07C4(7'b0111111);
								// Trace: design.sv:11039:17
								alu_vec_mode_o = cv32e40p_pkg_VEC_MODE8;
								// Trace: design.sv:11040:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:11041:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:11044:17
								illegal_insn_o = 1'b1;
						9'b000010000:
							// Trace: design.sv:11048:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11049:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010100);
								// Trace: design.sv:11050:17
								if (instr_rdata_i[24:20] != 5'b00000)
									// Trace: design.sv:11051:19
									illegal_insn_o = 1'b1;
							end
							else
								// Trace: design.sv:11054:17
								illegal_insn_o = 1'b1;
						9'b001010001:
							// Trace: design.sv:11058:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11059:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010110);
								// Trace: design.sv:11060:17
								alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
								// Trace: design.sv:11061:17
								imm_b_mux_sel_o = cv32e40p_pkg_IMMB_CLIP;
							end
							else
								// Trace: design.sv:11063:17
								illegal_insn_o = 1'b1;
						9'b001010010:
							// Trace: design.sv:11067:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11068:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010111);
								// Trace: design.sv:11069:17
								alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
								// Trace: design.sv:11070:17
								imm_b_mux_sel_o = cv32e40p_pkg_IMMB_CLIP;
							end
							else
								// Trace: design.sv:11072:17
								illegal_insn_o = 1'b1;
						9'b001010101:
							// Trace: design.sv:11076:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11077:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010110);
								// Trace: design.sv:11078:17
								regb_used_o = 1'b1;
							end
							else
								// Trace: design.sv:11080:17
								illegal_insn_o = 1'b1;
						9'b001010110:
							// Trace: design.sv:11084:15
							if (PULP_XPULP) begin
								// Trace: design.sv:11085:17
								alu_operator_o = sv2v_cast_C07C4(7'b0010111);
								// Trace: design.sv:11086:17
								regb_used_o = 1'b1;
							end
							else
								// Trace: design.sv:11088:17
								illegal_insn_o = 1'b1;
						default:
							// Trace: design.sv:11093:15
							illegal_insn_o = 1'b1;
					endcase
				end
			cv32e40p_pkg_OPCODE_OP_FP:
				// Trace: design.sv:11111:9
				if (FPU == 1) begin
					// Trace: design.sv:11114:11
					apu_en = 1'b1;
					// Trace: design.sv:11115:11
					alu_en = 1'b0;
					// Trace: design.sv:11117:11
					rega_used_o = 1'b1;
					// Trace: design.sv:11118:11
					regb_used_o = 1'b1;
					// Trace: design.sv:11119:11
					if (PULP_ZFINX == 0) begin
						// Trace: design.sv:11120:13
						reg_fp_a_o = 1'b1;
						// Trace: design.sv:11121:13
						reg_fp_b_o = 1'b1;
						// Trace: design.sv:11122:13
						reg_fp_d_o = 1'b1;
					end
					else begin
						// Trace: design.sv:11124:13
						reg_fp_a_o = 1'b0;
						// Trace: design.sv:11125:13
						reg_fp_b_o = 1'b0;
						// Trace: design.sv:11126:13
						reg_fp_d_o = 1'b0;
					end
					// Trace: design.sv:11129:11
					check_fprm = 1'b1;
					// Trace: design.sv:11130:11
					fp_rnd_mode_o = instr_rdata_i[14:12];
					(* full_case, parallel_case *)
					case (instr_rdata_i[26:25])
						2'b00:
							// Trace: design.sv:11135:20
							fpu_dst_fmt_o = sv2v_cast_9D6B6('d0);
						2'b01:
							// Trace: design.sv:11137:20
							fpu_dst_fmt_o = sv2v_cast_9D6B6('d1);
						2'b10:
							// Trace: design.sv:11141:15
							if (instr_rdata_i[14:12] == 3'b101)
								// Trace: design.sv:11141:49
								fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
							else
								// Trace: design.sv:11143:20
								fpu_dst_fmt_o = sv2v_cast_9D6B6('d2);
						2'b11:
							// Trace: design.sv:11146:20
							fpu_dst_fmt_o = sv2v_cast_9D6B6('d3);
					endcase
					// Trace: design.sv:11150:11
					fpu_src_fmt_o = fpu_dst_fmt_o;
					(* full_case, parallel_case *)
					case (instr_rdata_i[31:27])
						5'b00000: begin
							// Trace: design.sv:11156:15
							fpu_op = sv2v_cast_A1364(2);
							// Trace: design.sv:11157:15
							fp_op_group = 2'd0;
							// Trace: design.sv:11158:15
							apu_op_o = 2'b00;
							// Trace: design.sv:11159:15
							apu_lat_o = 2'h2;
							// Trace: design.sv:11160:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
							// Trace: design.sv:11161:15
							alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_REGB_OR_FWD;
						end
						5'b00001: begin
							// Trace: design.sv:11165:15
							fpu_op = sv2v_cast_A1364(2);
							// Trace: design.sv:11166:15
							fpu_op_mod = 1'b1;
							// Trace: design.sv:11167:15
							fp_op_group = 2'd0;
							// Trace: design.sv:11168:15
							apu_op_o = 2'b01;
							// Trace: design.sv:11169:15
							apu_lat_o = 2'h2;
							// Trace: design.sv:11170:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
							// Trace: design.sv:11171:15
							alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_REGB_OR_FWD;
						end
						5'b00010: begin
							// Trace: design.sv:11175:15
							fpu_op = sv2v_cast_A1364(3);
							// Trace: design.sv:11176:15
							fp_op_group = 2'd0;
							// Trace: design.sv:11177:15
							apu_lat_o = 2'h2;
						end
						5'b00011: begin
							// Trace: design.sv:11181:15
							fpu_op = sv2v_cast_A1364(4);
							// Trace: design.sv:11182:15
							fp_op_group = 2'd1;
							// Trace: design.sv:11183:15
							apu_lat_o = 2'h3;
						end
						5'b01011: begin
							// Trace: design.sv:11187:15
							regb_used_o = 1'b0;
							// Trace: design.sv:11188:15
							fpu_op = sv2v_cast_A1364(5);
							// Trace: design.sv:11189:15
							fp_op_group = 2'd1;
							// Trace: design.sv:11190:15
							apu_op_o = 1'b1;
							// Trace: design.sv:11191:15
							apu_lat_o = 2'h3;
							// Trace: design.sv:11193:15
							if (instr_rdata_i[24:20] != 5'b00000)
								// Trace: design.sv:11193:53
								illegal_insn_o = 1'b1;
						end
						5'b00100: begin
							// Trace: design.sv:11197:15
							fpu_op = sv2v_cast_A1364(6);
							// Trace: design.sv:11198:15
							fp_op_group = 2'd2;
							// Trace: design.sv:11199:15
							check_fprm = 1'b0;
							// Trace: design.sv:11200:15
							if (cv32e40p_pkg_C_XF16ALT) begin
								// Trace: design.sv:11201:17
								if (!(|{(3'b000 <= instr_rdata_i[14:12]) && (3'b010 >= instr_rdata_i[14:12]), (3'b100 <= instr_rdata_i[14:12]) && (3'b110 >= instr_rdata_i[14:12])}))
									// Trace: design.sv:11202:19
									illegal_insn_o = 1'b1;
								if (instr_rdata_i[14]) begin
									// Trace: design.sv:11206:19
									fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
									// Trace: design.sv:11207:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
								end
								else
									// Trace: design.sv:11209:19
									fp_rnd_mode_o = {1'b0, instr_rdata_i[13:12]};
							end
							else
								// Trace: design.sv:11212:17
								if (!((3'b000 <= instr_rdata_i[14:12]) && (3'b010 >= instr_rdata_i[14:12])))
									// Trace: design.sv:11212:71
									illegal_insn_o = 1'b1;
						end
						5'b00101: begin
							// Trace: design.sv:11217:15
							fpu_op = sv2v_cast_A1364(7);
							// Trace: design.sv:11218:15
							fp_op_group = 2'd2;
							// Trace: design.sv:11219:15
							check_fprm = 1'b0;
							// Trace: design.sv:11220:15
							if (cv32e40p_pkg_C_XF16ALT) begin
								// Trace: design.sv:11221:17
								if (!(|{(3'b000 <= instr_rdata_i[14:12]) && (3'b001 >= instr_rdata_i[14:12]), (3'b100 <= instr_rdata_i[14:12]) && (3'b101 >= instr_rdata_i[14:12])}))
									// Trace: design.sv:11222:19
									illegal_insn_o = 1'b1;
								if (instr_rdata_i[14]) begin
									// Trace: design.sv:11226:19
									fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
									// Trace: design.sv:11227:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
								end
								else
									// Trace: design.sv:11229:19
									fp_rnd_mode_o = {1'b0, instr_rdata_i[13:12]};
							end
							else
								// Trace: design.sv:11232:17
								if (!((3'b000 <= instr_rdata_i[14:12]) && (3'b001 >= instr_rdata_i[14:12])))
									// Trace: design.sv:11232:71
									illegal_insn_o = 1'b1;
						end
						5'b01000: begin
							// Trace: design.sv:11237:15
							regb_used_o = 1'b0;
							// Trace: design.sv:11238:15
							fpu_op = sv2v_cast_A1364(10);
							// Trace: design.sv:11239:15
							fp_op_group = 2'd3;
							// Trace: design.sv:11241:15
							if (instr_rdata_i[24:23])
								// Trace: design.sv:11241:41
								illegal_insn_o = 1'b1;
							(* full_case, parallel_case *)
							case (instr_rdata_i[22:20])
								3'b000: begin
									// Trace: design.sv:11246:19
									if (~cv32e40p_pkg_C_RVF)
										// Trace: design.sv:11246:31
										illegal_insn_o = 1'b1;
									// Trace: design.sv:11247:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d0);
								end
								3'b001: begin
									// Trace: design.sv:11250:19
									if (~cv32e40p_pkg_C_RVD)
										// Trace: design.sv:11250:31
										illegal_insn_o = 1'b1;
									// Trace: design.sv:11251:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d1);
								end
								3'b010: begin
									// Trace: design.sv:11254:19
									if (~cv32e40p_pkg_C_XF16)
										// Trace: design.sv:11254:32
										illegal_insn_o = 1'b1;
									// Trace: design.sv:11255:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d2);
								end
								3'b110: begin
									// Trace: design.sv:11258:19
									if (~cv32e40p_pkg_C_XF16ALT)
										// Trace: design.sv:11258:35
										illegal_insn_o = 1'b1;
									// Trace: design.sv:11259:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
								end
								3'b011: begin
									// Trace: design.sv:11262:19
									if (~cv32e40p_pkg_C_XF8)
										// Trace: design.sv:11262:31
										illegal_insn_o = 1'b1;
									// Trace: design.sv:11263:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d3);
								end
								default:
									// Trace: design.sv:11265:26
									illegal_insn_o = 1'b1;
							endcase
						end
						5'b01001: begin
							// Trace: design.sv:11270:15
							fpu_op = sv2v_cast_A1364(3);
							// Trace: design.sv:11271:15
							fp_op_group = 2'd0;
							// Trace: design.sv:11272:15
							apu_lat_o = 2'h2;
							// Trace: design.sv:11274:15
							fpu_dst_fmt_o = sv2v_cast_9D6B6('d0);
						end
						5'b01010: begin
							// Trace: design.sv:11278:15
							regc_used_o = 1'b1;
							// Trace: design.sv:11279:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:11280:15
							if (PULP_ZFINX == 0)
								// Trace: design.sv:11281:17
								reg_fp_c_o = 1'b1;
							else
								// Trace: design.sv:11283:17
								reg_fp_c_o = 1'b0;
							// Trace: design.sv:11285:15
							fpu_op = sv2v_cast_A1364(0);
							// Trace: design.sv:11286:15
							fp_op_group = 2'd0;
							// Trace: design.sv:11287:15
							apu_lat_o = 2'h2;
							// Trace: design.sv:11289:15
							fpu_dst_fmt_o = sv2v_cast_9D6B6('d0);
						end
						5'b10100: begin
							// Trace: design.sv:11293:15
							fpu_op = sv2v_cast_A1364(8);
							// Trace: design.sv:11294:15
							fp_op_group = 2'd2;
							// Trace: design.sv:11295:15
							reg_fp_d_o = 1'b0;
							// Trace: design.sv:11296:15
							check_fprm = 1'b0;
							// Trace: design.sv:11297:15
							if (cv32e40p_pkg_C_XF16ALT) begin
								// Trace: design.sv:11298:17
								if (!(|{(3'b000 <= instr_rdata_i[14:12]) && (3'b010 >= instr_rdata_i[14:12]), (3'b100 <= instr_rdata_i[14:12]) && (3'b110 >= instr_rdata_i[14:12])}))
									// Trace: design.sv:11299:19
									illegal_insn_o = 1'b1;
								if (instr_rdata_i[14]) begin
									// Trace: design.sv:11303:19
									fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
									// Trace: design.sv:11304:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
								end
								else
									// Trace: design.sv:11306:19
									fp_rnd_mode_o = {1'b0, instr_rdata_i[13:12]};
							end
							else
								// Trace: design.sv:11309:17
								if (!((3'b000 <= instr_rdata_i[14:12]) && (3'b010 >= instr_rdata_i[14:12])))
									// Trace: design.sv:11309:71
									illegal_insn_o = 1'b1;
						end
						5'b11000: begin
							// Trace: design.sv:11314:15
							regb_used_o = 1'b0;
							// Trace: design.sv:11315:15
							reg_fp_d_o = 1'b0;
							// Trace: design.sv:11316:15
							fpu_op = sv2v_cast_A1364(11);
							// Trace: design.sv:11317:15
							fp_op_group = 2'd3;
							// Trace: design.sv:11318:15
							fpu_op_mod = instr_rdata_i[20];
							// Trace: design.sv:11319:15
							apu_op_o = 2'b01;
							// Trace: design.sv:11320:15
							apu_lat_o = 2'h2;
							// Trace: design.sv:11322:15
							(* full_case, parallel_case *)
							case (instr_rdata_i[26:25])
								2'b00:
									// Trace: design.sv:11324:19
									if (~cv32e40p_pkg_C_RVF)
										// Trace: design.sv:11324:31
										illegal_insn_o = 1;
									else
										// Trace: design.sv:11325:24
										fpu_src_fmt_o = sv2v_cast_9D6B6('d0);
								2'b01:
									// Trace: design.sv:11328:19
									if (~cv32e40p_pkg_C_RVD)
										// Trace: design.sv:11328:31
										illegal_insn_o = 1;
									else
										// Trace: design.sv:11329:24
										fpu_src_fmt_o = sv2v_cast_9D6B6('d1);
								2'b10:
									// Trace: design.sv:11332:19
									if (instr_rdata_i[14:12] == 3'b101) begin
										begin
											// Trace: design.sv:11333:21
											if (~cv32e40p_pkg_C_XF16ALT)
												// Trace: design.sv:11333:37
												illegal_insn_o = 1;
											else
												// Trace: design.sv:11334:26
												fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
										end
									end
									else if (~cv32e40p_pkg_C_XF16)
										// Trace: design.sv:11336:21
										illegal_insn_o = 1;
									else
										// Trace: design.sv:11338:21
										fpu_src_fmt_o = sv2v_cast_9D6B6('d2);
								2'b11:
									// Trace: design.sv:11342:19
									if (~cv32e40p_pkg_C_XF8)
										// Trace: design.sv:11342:31
										illegal_insn_o = 1;
									else
										// Trace: design.sv:11343:24
										fpu_src_fmt_o = sv2v_cast_9D6B6('d3);
							endcase
							if (instr_rdata_i[24:21])
								// Trace: design.sv:11347:41
								illegal_insn_o = 1'b1;
						end
						5'b11010: begin
							// Trace: design.sv:11351:15
							regb_used_o = 1'b0;
							// Trace: design.sv:11352:15
							reg_fp_a_o = 1'b0;
							// Trace: design.sv:11353:15
							fpu_op = sv2v_cast_A1364(12);
							// Trace: design.sv:11354:15
							fp_op_group = 2'd3;
							// Trace: design.sv:11355:15
							fpu_op_mod = instr_rdata_i[20];
							// Trace: design.sv:11356:15
							apu_op_o = 2'b00;
							// Trace: design.sv:11357:15
							apu_lat_o = 2'h2;
							// Trace: design.sv:11359:15
							if (instr_rdata_i[24:21])
								// Trace: design.sv:11359:41
								illegal_insn_o = 1'b1;
						end
						5'b11100: begin
							// Trace: design.sv:11363:15
							regb_used_o = 1'b0;
							// Trace: design.sv:11364:15
							reg_fp_d_o = 1'b0;
							// Trace: design.sv:11365:15
							fp_op_group = 2'd2;
							// Trace: design.sv:11366:15
							check_fprm = 1'b0;
							// Trace: design.sv:11368:15
							if ((instr_rdata_i[14:12] == 3'b000) || 1'd0) begin
								// Trace: design.sv:11369:17
								alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
								// Trace: design.sv:11370:17
								fpu_op = sv2v_cast_A1364(6);
								// Trace: design.sv:11371:17
								fpu_op_mod = 1'b1;
								// Trace: design.sv:11372:17
								fp_rnd_mode_o = 3'b011;
								// Trace: design.sv:11374:17
								if (instr_rdata_i[14]) begin
									// Trace: design.sv:11375:19
									fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
									// Trace: design.sv:11376:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
								end
							end
							else if ((instr_rdata_i[14:12] == 3'b001) || 1'd0) begin
								// Trace: design.sv:11380:17
								fpu_op = sv2v_cast_A1364(9);
								// Trace: design.sv:11381:17
								fp_rnd_mode_o = 3'b000;
								// Trace: design.sv:11383:17
								if (instr_rdata_i[14]) begin
									// Trace: design.sv:11384:19
									fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
									// Trace: design.sv:11385:19
									fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
								end
							end
							else
								// Trace: design.sv:11388:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[24:20])
								// Trace: design.sv:11391:41
								illegal_insn_o = 1'b1;
						end
						5'b11110: begin
							// Trace: design.sv:11395:15
							regb_used_o = 1'b0;
							// Trace: design.sv:11396:15
							reg_fp_a_o = 1'b0;
							// Trace: design.sv:11397:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
							// Trace: design.sv:11398:15
							fpu_op = sv2v_cast_A1364(6);
							// Trace: design.sv:11399:15
							fpu_op_mod = 1'b0;
							// Trace: design.sv:11400:15
							fp_op_group = 2'd2;
							// Trace: design.sv:11401:15
							fp_rnd_mode_o = 3'b011;
							// Trace: design.sv:11402:15
							check_fprm = 1'b0;
							// Trace: design.sv:11403:15
							if ((instr_rdata_i[14:12] == 3'b000) || 1'd0) begin
								begin
									// Trace: design.sv:11405:17
									if (instr_rdata_i[14]) begin
										// Trace: design.sv:11406:19
										fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
										// Trace: design.sv:11407:19
										fpu_src_fmt_o = sv2v_cast_9D6B6('d4);
									end
								end
							end
							else
								// Trace: design.sv:11410:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[24:20] != 5'b00000)
								// Trace: design.sv:11413:53
								illegal_insn_o = 1'b1;
						end
						default:
							// Trace: design.sv:11417:15
							illegal_insn_o = 1'b1;
					endcase
					if (~cv32e40p_pkg_C_RVF && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d0)))
						// Trace: design.sv:11422:66
						illegal_insn_o = 1'b1;
					if (~cv32e40p_pkg_C_RVD && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d1)))
						// Trace: design.sv:11423:68
						illegal_insn_o = 1'b1;
					if (~cv32e40p_pkg_C_XF16 && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d2)))
						// Trace: design.sv:11424:69
						illegal_insn_o = 1'b1;
					if (~cv32e40p_pkg_C_XF16ALT && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d4)))
						// Trace: design.sv:11426:13
						illegal_insn_o = 1'b1;
					if (~cv32e40p_pkg_C_XF8 && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d3)))
						// Trace: design.sv:11428:67
						illegal_insn_o = 1'b1;
					if (check_fprm) begin
						begin
							// Trace: design.sv:11432:13
							(* full_case, parallel_case *)
							if ((3'b000 <= instr_rdata_i[14:12]) && (3'b100 >= instr_rdata_i[14:12]))
								;
							else if (instr_rdata_i[14:12] == 3'b101) begin
								// Trace: design.sv:11435:17
								if (~cv32e40p_pkg_C_XF16ALT || (fpu_dst_fmt_o != sv2v_cast_9D6B6('d4)))
									// Trace: design.sv:11435:79
									illegal_insn_o = 1'b1;
								(* full_case, parallel_case *)
								if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
									// Trace: design.sv:11438:37
									fp_rnd_mode_o = frm_i;
								else
									// Trace: design.sv:11439:37
									illegal_insn_o = 1'b1;
							end
							else if (instr_rdata_i[14:12] == 3'b111) begin
								begin
									// Trace: design.sv:11444:17
									(* full_case, parallel_case *)
									if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
										// Trace: design.sv:11445:37
										fp_rnd_mode_o = frm_i;
									else
										// Trace: design.sv:11446:37
										illegal_insn_o = 1'b1;
								end
							end
							else
								// Trace: design.sv:11449:25
								illegal_insn_o = 1'b1;
						end
					end
					case (fp_op_group)
						2'd0:
							// Trace: design.sv:11459:15
							(* full_case, parallel_case *)
							case (fpu_dst_fmt_o)
								sv2v_cast_9D6B6('d0):
									// Trace: design.sv:11460:45
									apu_lat_o = 1;
								sv2v_cast_9D6B6('d1):
									// Trace: design.sv:11461:45
									apu_lat_o = 1;
								sv2v_cast_9D6B6('d2):
									// Trace: design.sv:11462:45
									apu_lat_o = 1;
								sv2v_cast_9D6B6('d4):
									// Trace: design.sv:11463:45
									apu_lat_o = 1;
								sv2v_cast_9D6B6('d3):
									// Trace: design.sv:11464:45
									apu_lat_o = 1;
								default:
									;
							endcase
						2'd1:
							// Trace: design.sv:11469:23
							apu_lat_o = 2'h3;
						2'd2:
							// Trace: design.sv:11471:23
							apu_lat_o = 1;
						2'd3:
							// Trace: design.sv:11473:23
							apu_lat_o = 1;
					endcase
					// Trace: design.sv:11477:11
					apu_op_o = {fpu_vec_op, fpu_op_mod, fpu_op};
				end
				else
					// Trace: design.sv:11482:11
					illegal_insn_o = 1'b1;
			cv32e40p_pkg_OPCODE_OP_FMADD, cv32e40p_pkg_OPCODE_OP_FMSUB, cv32e40p_pkg_OPCODE_OP_FNMSUB, cv32e40p_pkg_OPCODE_OP_FNMADD:
				// Trace: design.sv:11490:9
				if (FPU == 1) begin
					// Trace: design.sv:11492:11
					apu_en = 1'b1;
					// Trace: design.sv:11493:11
					alu_en = 1'b0;
					// Trace: design.sv:11494:11
					apu_lat_o = 2'h3;
					// Trace: design.sv:11496:11
					rega_used_o = 1'b1;
					// Trace: design.sv:11497:11
					regb_used_o = 1'b1;
					// Trace: design.sv:11498:11
					regc_used_o = 1'b1;
					// Trace: design.sv:11499:11
					regc_mux_o = cv32e40p_pkg_REGC_S4;
					// Trace: design.sv:11500:11
					if (PULP_ZFINX == 0) begin
						// Trace: design.sv:11501:13
						reg_fp_a_o = 1'b1;
						// Trace: design.sv:11502:13
						reg_fp_b_o = 1'b1;
						// Trace: design.sv:11503:13
						reg_fp_c_o = 1'b1;
						// Trace: design.sv:11504:13
						reg_fp_d_o = 1'b1;
					end
					else begin
						// Trace: design.sv:11506:13
						reg_fp_a_o = 1'b0;
						// Trace: design.sv:11507:13
						reg_fp_b_o = 1'b0;
						// Trace: design.sv:11508:13
						reg_fp_c_o = 1'b0;
						// Trace: design.sv:11509:13
						reg_fp_d_o = 1'b0;
					end
					// Trace: design.sv:11511:11
					fp_rnd_mode_o = instr_rdata_i[14:12];
					(* full_case, parallel_case *)
					case (instr_rdata_i[26:25])
						2'b00:
							// Trace: design.sv:11516:21
							fpu_dst_fmt_o = sv2v_cast_9D6B6('d0);
						2'b01:
							// Trace: design.sv:11518:21
							fpu_dst_fmt_o = sv2v_cast_9D6B6('d1);
						2'b10:
							// Trace: design.sv:11522:15
							if (instr_rdata_i[14:12] == 3'b101)
								// Trace: design.sv:11522:49
								fpu_dst_fmt_o = sv2v_cast_9D6B6('d4);
							else
								// Trace: design.sv:11523:20
								fpu_dst_fmt_o = sv2v_cast_9D6B6('d2);
						2'b11:
							// Trace: design.sv:11526:21
							fpu_dst_fmt_o = sv2v_cast_9D6B6('d3);
					endcase
					// Trace: design.sv:11530:11
					fpu_src_fmt_o = fpu_dst_fmt_o;
					(* full_case, parallel_case *)
					case (instr_rdata_i[6:0])
						cv32e40p_pkg_OPCODE_OP_FMADD: begin
							// Trace: design.sv:11536:15
							fpu_op = sv2v_cast_A1364(0);
							// Trace: design.sv:11537:15
							apu_op_o = 2'b00;
						end
						cv32e40p_pkg_OPCODE_OP_FMSUB: begin
							// Trace: design.sv:11541:15
							fpu_op = sv2v_cast_A1364(0);
							// Trace: design.sv:11542:15
							fpu_op_mod = 1'b1;
							// Trace: design.sv:11543:15
							apu_op_o = 2'b01;
						end
						cv32e40p_pkg_OPCODE_OP_FNMSUB: begin
							// Trace: design.sv:11547:15
							fpu_op = sv2v_cast_A1364(1);
							// Trace: design.sv:11548:15
							apu_op_o = 2'b10;
						end
						cv32e40p_pkg_OPCODE_OP_FNMADD: begin
							// Trace: design.sv:11552:15
							fpu_op = sv2v_cast_A1364(1);
							// Trace: design.sv:11553:15
							fpu_op_mod = 1'b1;
							// Trace: design.sv:11554:15
							apu_op_o = 2'b11;
						end
					endcase
					if (~cv32e40p_pkg_C_RVF && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d0)))
						// Trace: design.sv:11559:66
						illegal_insn_o = 1'b1;
					if (~cv32e40p_pkg_C_RVD && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d1)))
						// Trace: design.sv:11560:68
						illegal_insn_o = 1'b1;
					if (~cv32e40p_pkg_C_XF16 && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d2)))
						// Trace: design.sv:11561:69
						illegal_insn_o = 1'b1;
					if (~cv32e40p_pkg_C_XF16ALT && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d4)))
						// Trace: design.sv:11563:13
						illegal_insn_o = 1'b1;
					if (~cv32e40p_pkg_C_XF8 && (fpu_dst_fmt_o == sv2v_cast_9D6B6('d3)))
						// Trace: design.sv:11565:67
						illegal_insn_o = 1'b1;
					(* full_case, parallel_case *)
					if ((3'b000 <= instr_rdata_i[14:12]) && (3'b100 >= instr_rdata_i[14:12]))
						;
					else if (instr_rdata_i[14:12] == 3'b101) begin
						// Trace: design.sv:11571:15
						if (~cv32e40p_pkg_C_XF16ALT || (fpu_dst_fmt_o != sv2v_cast_9D6B6('d4)))
							// Trace: design.sv:11571:77
							illegal_insn_o = 1'b1;
						(* full_case, parallel_case *)
						if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
							// Trace: design.sv:11574:35
							fp_rnd_mode_o = frm_i;
						else
							// Trace: design.sv:11575:35
							illegal_insn_o = 1'b1;
					end
					else if (instr_rdata_i[14:12] == 3'b111) begin
						begin
							// Trace: design.sv:11580:15
							(* full_case, parallel_case *)
							if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
								// Trace: design.sv:11581:35
								fp_rnd_mode_o = frm_i;
							else
								// Trace: design.sv:11582:35
								illegal_insn_o = 1'b1;
						end
					end
					else
						// Trace: design.sv:11585:23
						illegal_insn_o = 1'b1;
					(* full_case, parallel_case *)
					case (fpu_dst_fmt_o)
						sv2v_cast_9D6B6('d0):
							// Trace: design.sv:11593:41
							apu_lat_o = 1;
						sv2v_cast_9D6B6('d1):
							// Trace: design.sv:11594:41
							apu_lat_o = 1;
						sv2v_cast_9D6B6('d2):
							// Trace: design.sv:11595:41
							apu_lat_o = 1;
						sv2v_cast_9D6B6('d4):
							// Trace: design.sv:11596:41
							apu_lat_o = 1;
						sv2v_cast_9D6B6('d3):
							// Trace: design.sv:11597:41
							apu_lat_o = 1;
						default:
							;
					endcase
					// Trace: design.sv:11602:11
					apu_op_o = {fpu_vec_op, fpu_op_mod, fpu_op};
				end
				else
					// Trace: design.sv:11606:11
					illegal_insn_o = 1'b1;
			cv32e40p_pkg_OPCODE_STORE_FP:
				// Trace: design.sv:11611:9
				if (FPU == 1) begin
					// Trace: design.sv:11612:11
					data_req = 1'b1;
					// Trace: design.sv:11613:11
					data_we_o = 1'b1;
					// Trace: design.sv:11614:11
					rega_used_o = 1'b1;
					// Trace: design.sv:11615:11
					regb_used_o = 1'b1;
					// Trace: design.sv:11616:11
					alu_operator_o = sv2v_cast_C07C4(7'b0011000);
					// Trace: design.sv:11617:11
					if (PULP_ZFINX == 0)
						// Trace: design.sv:11618:13
						reg_fp_b_o = 1'b1;
					else
						// Trace: design.sv:11620:13
						reg_fp_b_o = 1'b0;
					// Trace: design.sv:11624:11
					imm_b_mux_sel_o = cv32e40p_pkg_IMMB_S;
					// Trace: design.sv:11625:11
					alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
					// Trace: design.sv:11628:11
					alu_op_c_mux_sel_o = cv32e40p_pkg_OP_C_REGB_OR_FWD;
					(* full_case, parallel_case *)
					case (instr_rdata_i[14:12])
						3'b000:
							if (cv32e40p_pkg_C_XF8)
								// Trace: design.sv:11633:33
								data_type_o = 2'b10;
							else
								// Trace: design.sv:11634:27
								illegal_insn_o = 1'b1;
						3'b001:
							if (cv32e40p_pkg_C_XF16 | cv32e40p_pkg_C_XF16ALT)
								// Trace: design.sv:11636:46
								data_type_o = 2'b01;
							else
								// Trace: design.sv:11637:27
								illegal_insn_o = 1'b1;
						3'b010:
							if (cv32e40p_pkg_C_RVF)
								// Trace: design.sv:11639:33
								data_type_o = 2'b00;
							else
								// Trace: design.sv:11640:27
								illegal_insn_o = 1'b1;
						3'b011:
							if (cv32e40p_pkg_C_RVD)
								// Trace: design.sv:11642:33
								data_type_o = 2'b00;
							else
								// Trace: design.sv:11643:27
								illegal_insn_o = 1'b1;
						default:
							// Trace: design.sv:11644:22
							illegal_insn_o = 1'b1;
					endcase
					if (illegal_insn_o) begin
						// Trace: design.sv:11649:13
						data_req = 1'b0;
						// Trace: design.sv:11650:13
						data_we_o = 1'b0;
					end
				end
				else
					// Trace: design.sv:11655:11
					illegal_insn_o = 1'b1;
			cv32e40p_pkg_OPCODE_LOAD_FP:
				// Trace: design.sv:11659:9
				if (FPU == 1) begin
					// Trace: design.sv:11660:11
					data_req = 1'b1;
					// Trace: design.sv:11661:11
					regfile_mem_we = 1'b1;
					// Trace: design.sv:11662:11
					if (PULP_ZFINX == 0)
						// Trace: design.sv:11663:13
						reg_fp_d_o = 1'b1;
					else
						// Trace: design.sv:11665:13
						reg_fp_d_o = 1'b0;
					// Trace: design.sv:11667:11
					rega_used_o = 1'b1;
					// Trace: design.sv:11668:11
					alu_operator_o = sv2v_cast_C07C4(7'b0011000);
					// Trace: design.sv:11671:11
					imm_b_mux_sel_o = cv32e40p_pkg_IMMB_I;
					// Trace: design.sv:11672:11
					alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
					// Trace: design.sv:11675:11
					data_sign_extension_o = 2'b10;
					(* full_case, parallel_case *)
					case (instr_rdata_i[14:12])
						3'b000:
							if (cv32e40p_pkg_C_XF8)
								// Trace: design.sv:11680:33
								data_type_o = 2'b10;
							else
								// Trace: design.sv:11681:27
								illegal_insn_o = 1'b1;
						3'b001:
							if (cv32e40p_pkg_C_XF16 | cv32e40p_pkg_C_XF16ALT)
								// Trace: design.sv:11683:46
								data_type_o = 2'b01;
							else
								// Trace: design.sv:11684:27
								illegal_insn_o = 1'b1;
						3'b010:
							if (cv32e40p_pkg_C_RVF)
								// Trace: design.sv:11686:33
								data_type_o = 2'b00;
							else
								// Trace: design.sv:11687:27
								illegal_insn_o = 1'b1;
						3'b011:
							if (cv32e40p_pkg_C_RVD)
								// Trace: design.sv:11689:33
								data_type_o = 2'b00;
							else
								// Trace: design.sv:11690:27
								illegal_insn_o = 1'b1;
						default:
							// Trace: design.sv:11691:22
							illegal_insn_o = 1'b1;
					endcase
				end
				else
					// Trace: design.sv:11696:11
					illegal_insn_o = 1'b1;
			cv32e40p_pkg_OPCODE_PULP_OP:
				// Trace: design.sv:11700:9
				if (PULP_XPULP) begin
					// Trace: design.sv:11701:11
					regfile_alu_we = 1'b1;
					// Trace: design.sv:11702:11
					rega_used_o = 1'b1;
					// Trace: design.sv:11703:11
					regb_used_o = 1'b1;
					// Trace: design.sv:11705:11
					case (instr_rdata_i[13:12])
						2'b00: begin
							// Trace: design.sv:11707:15
							alu_en = 1'b0;
							// Trace: design.sv:11709:15
							mult_sel_subword_o = instr_rdata_i[30];
							// Trace: design.sv:11710:15
							mult_signed_mode_o = {2 {instr_rdata_i[31]}};
							// Trace: design.sv:11712:15
							mult_imm_mux_o = cv32e40p_pkg_MIMM_S3;
							// Trace: design.sv:11713:15
							regc_mux_o = cv32e40p_pkg_REGC_ZERO;
							// Trace: design.sv:11714:15
							mult_int_en = 1'b1;
							// Trace: design.sv:11716:15
							if (instr_rdata_i[14])
								// Trace: design.sv:11717:17
								mult_operator_o = sv2v_cast_9F558(3'b011);
							else
								// Trace: design.sv:11719:17
								mult_operator_o = sv2v_cast_9F558(3'b010);
						end
						2'b01: begin
							// Trace: design.sv:11723:15
							alu_en = 1'b0;
							// Trace: design.sv:11725:15
							mult_sel_subword_o = instr_rdata_i[30];
							// Trace: design.sv:11726:15
							mult_signed_mode_o = {2 {instr_rdata_i[31]}};
							// Trace: design.sv:11728:15
							regc_used_o = 1'b1;
							// Trace: design.sv:11729:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:11730:15
							mult_imm_mux_o = cv32e40p_pkg_MIMM_S3;
							// Trace: design.sv:11731:15
							mult_int_en = 1'b1;
							// Trace: design.sv:11733:15
							if (instr_rdata_i[14])
								// Trace: design.sv:11734:17
								mult_operator_o = sv2v_cast_9F558(3'b011);
							else
								// Trace: design.sv:11736:17
								mult_operator_o = sv2v_cast_9F558(3'b010);
						end
						2'b10: begin
							// Trace: design.sv:11742:15
							case ({instr_rdata_i[31], instr_rdata_i[14]})
								2'b00:
									// Trace: design.sv:11743:24
									alu_operator_o = sv2v_cast_C07C4(7'b0011000);
								2'b01:
									// Trace: design.sv:11744:24
									alu_operator_o = sv2v_cast_C07C4(7'b0011100);
								2'b10:
									// Trace: design.sv:11745:24
									alu_operator_o = sv2v_cast_C07C4(7'b0011010);
								2'b11:
									// Trace: design.sv:11746:24
									alu_operator_o = sv2v_cast_C07C4(7'b0011110);
							endcase
							// Trace: design.sv:11749:15
							bmask_a_mux_o = cv32e40p_pkg_BMASK_A_ZERO;
							// Trace: design.sv:11750:15
							bmask_b_mux_o = cv32e40p_pkg_BMASK_B_S3;
							if (instr_rdata_i[30]) begin
								// Trace: design.sv:11754:17
								regc_used_o = 1'b1;
								// Trace: design.sv:11755:17
								regc_mux_o = cv32e40p_pkg_REGC_RD;
								// Trace: design.sv:11756:17
								alu_bmask_b_mux_sel_o = cv32e40p_pkg_BMASK_B_REG;
								// Trace: design.sv:11757:17
								alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGC_OR_FWD;
								// Trace: design.sv:11758:17
								alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
								// Trace: design.sv:11759:17
								if (instr_rdata_i[29:25] != 5'b00000)
									// Trace: design.sv:11760:19
									illegal_insn_o = 1'b1;
							end
						end
						2'b11: begin
							// Trace: design.sv:11769:15
							case ({instr_rdata_i[31], instr_rdata_i[14]})
								2'b00:
									// Trace: design.sv:11770:24
									alu_operator_o = sv2v_cast_C07C4(7'b0011001);
								2'b01:
									// Trace: design.sv:11771:24
									alu_operator_o = sv2v_cast_C07C4(7'b0011101);
								2'b10:
									// Trace: design.sv:11772:24
									alu_operator_o = sv2v_cast_C07C4(7'b0011011);
								2'b11:
									// Trace: design.sv:11773:24
									alu_operator_o = sv2v_cast_C07C4(7'b0011111);
							endcase
							// Trace: design.sv:11776:15
							bmask_a_mux_o = cv32e40p_pkg_BMASK_A_ZERO;
							// Trace: design.sv:11777:15
							bmask_b_mux_o = cv32e40p_pkg_BMASK_B_S3;
							if (instr_rdata_i[30]) begin
								// Trace: design.sv:11781:17
								regc_used_o = 1'b1;
								// Trace: design.sv:11782:17
								regc_mux_o = cv32e40p_pkg_REGC_RD;
								// Trace: design.sv:11783:17
								alu_bmask_b_mux_sel_o = cv32e40p_pkg_BMASK_B_REG;
								// Trace: design.sv:11784:17
								alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGC_OR_FWD;
								// Trace: design.sv:11785:17
								alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGA_OR_FWD;
								// Trace: design.sv:11786:17
								if (instr_rdata_i[29:25] != 5'b00000)
									// Trace: design.sv:11787:19
									illegal_insn_o = 1'b1;
							end
						end
					endcase
				end
				else
					// Trace: design.sv:11794:11
					illegal_insn_o = 1'b1;
			cv32e40p_pkg_OPCODE_VECOP:
				// Trace: design.sv:11799:9
				if (PULP_XPULP) begin
					// Trace: design.sv:11800:11
					regfile_alu_we = 1'b1;
					// Trace: design.sv:11801:11
					rega_used_o = 1'b1;
					// Trace: design.sv:11802:11
					imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
					// Trace: design.sv:11805:11
					if (instr_rdata_i[12]) begin
						// Trace: design.sv:11806:13
						alu_vec_mode_o = cv32e40p_pkg_VEC_MODE8;
						// Trace: design.sv:11807:13
						mult_operator_o = sv2v_cast_9F558(3'b100);
					end
					else begin
						// Trace: design.sv:11809:13
						alu_vec_mode_o = cv32e40p_pkg_VEC_MODE16;
						// Trace: design.sv:11810:13
						mult_operator_o = sv2v_cast_9F558(3'b101);
					end
					if (instr_rdata_i[14]) begin
						// Trace: design.sv:11815:13
						scalar_replication_o = 1'b1;
						// Trace: design.sv:11817:13
						if (instr_rdata_i[13])
							// Trace: design.sv:11819:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
						else
							// Trace: design.sv:11822:15
							regb_used_o = 1'b1;
					end
					else
						// Trace: design.sv:11826:13
						regb_used_o = 1'b1;
					(* full_case, parallel_case *)
					case (instr_rdata_i[31:26])
						6'b000000: begin
							// Trace: design.sv:11832:15
							alu_operator_o = sv2v_cast_C07C4(7'b0011000);
							// Trace: design.sv:11833:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11834:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11835:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11838:17
								illegal_insn_o = 1'b1;
						end
						6'b000010: begin
							// Trace: design.sv:11842:15
							alu_operator_o = sv2v_cast_C07C4(7'b0011001);
							// Trace: design.sv:11843:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11844:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11845:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11848:17
								illegal_insn_o = 1'b1;
						end
						6'b000100: begin
							// Trace: design.sv:11852:15
							alu_operator_o = sv2v_cast_C07C4(7'b0011000);
							// Trace: design.sv:11853:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11854:15
							bmask_b_mux_o = cv32e40p_pkg_BMASK_B_ONE;
							// Trace: design.sv:11855:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11856:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11859:17
								illegal_insn_o = 1'b1;
						end
						6'b000110: begin
							// Trace: design.sv:11863:14
							alu_operator_o = sv2v_cast_C07C4(7'b0011010);
							// Trace: design.sv:11864:14
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:11865:14
							bmask_b_mux_o = cv32e40p_pkg_BMASK_B_ONE;
							// Trace: design.sv:11866:14
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11867:16
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11870:16
								illegal_insn_o = 1'b1;
						end
						6'b001000: begin
							// Trace: design.sv:11874:14
							alu_operator_o = sv2v_cast_C07C4(7'b0010000);
							// Trace: design.sv:11875:14
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11876:14
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11877:16
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11880:16
								illegal_insn_o = 1'b1;
						end
						6'b001010: begin
							// Trace: design.sv:11884:15
							alu_operator_o = sv2v_cast_C07C4(7'b0010001);
							// Trace: design.sv:11885:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:11886:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11887:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11890:17
								illegal_insn_o = 1'b1;
						end
						6'b001100: begin
							// Trace: design.sv:11894:15
							alu_operator_o = sv2v_cast_C07C4(7'b0010010);
							// Trace: design.sv:11895:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11896:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11897:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11900:17
								illegal_insn_o = 1'b1;
						end
						6'b001110: begin
							// Trace: design.sv:11904:15
							alu_operator_o = sv2v_cast_C07C4(7'b0010011);
							// Trace: design.sv:11905:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:11906:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11907:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11910:17
								illegal_insn_o = 1'b1;
						end
						6'b010000: begin
							// Trace: design.sv:11914:15
							alu_operator_o = sv2v_cast_C07C4(7'b0100101);
							// Trace: design.sv:11915:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11916:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11917:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11920:17
								illegal_insn_o = 1'b1;
						end
						6'b010010: begin
							// Trace: design.sv:11924:15
							alu_operator_o = sv2v_cast_C07C4(7'b0100100);
							// Trace: design.sv:11925:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11926:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11927:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11930:17
								illegal_insn_o = 1'b1;
						end
						6'b010100: begin
							// Trace: design.sv:11934:15
							alu_operator_o = sv2v_cast_C07C4(7'b0100111);
							// Trace: design.sv:11935:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11936:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11937:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11940:17
								illegal_insn_o = 1'b1;
						end
						6'b010110: begin
							// Trace: design.sv:11944:15
							alu_operator_o = sv2v_cast_C07C4(7'b0101110);
							// Trace: design.sv:11945:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11946:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11947:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11950:17
								illegal_insn_o = 1'b1;
						end
						6'b011000: begin
							// Trace: design.sv:11954:15
							alu_operator_o = sv2v_cast_C07C4(7'b0101111);
							// Trace: design.sv:11955:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11956:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11957:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11960:17
								illegal_insn_o = 1'b1;
						end
						6'b011010: begin
							// Trace: design.sv:11964:15
							alu_operator_o = sv2v_cast_C07C4(7'b0010101);
							// Trace: design.sv:11965:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11966:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:11967:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11970:17
								illegal_insn_o = 1'b1;
						end
						6'b011100: begin
							// Trace: design.sv:11974:15
							alu_operator_o = sv2v_cast_C07C4(7'b0010100);
							// Trace: design.sv:11975:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:11976:15
							if (!((instr_rdata_i[14:12] == 3'b000) || (instr_rdata_i[14:12] == 3'b001)))
								// Trace: design.sv:11977:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[25:20] != 6'b000000)
								// Trace: design.sv:11980:17
								illegal_insn_o = 1'b1;
						end
						6'b110000: begin
							// Trace: design.sv:11984:15
							alu_operator_o = sv2v_cast_C07C4(7'b0111010);
							// Trace: design.sv:11985:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_SHUF;
							// Trace: design.sv:11986:15
							regb_used_o = 1'b1;
							// Trace: design.sv:11987:15
							scalar_replication_o = 1'b0;
							// Trace: design.sv:11988:15
							if ((((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011)) || (instr_rdata_i[14:12] == 3'b100)) || (instr_rdata_i[14:12] == 3'b101))
								// Trace: design.sv:11990:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:11993:17
								illegal_insn_o = 1'b1;
						end
						6'b111010, 6'b111100, 6'b111110: begin
							// Trace: design.sv:11999:15
							alu_operator_o = sv2v_cast_C07C4(7'b0111010);
							// Trace: design.sv:12000:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_SHUF;
							// Trace: design.sv:12001:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12002:15
							scalar_replication_o = 1'b0;
							// Trace: design.sv:12003:15
							if (instr_rdata_i[14:12] != 3'b111)
								// Trace: design.sv:12004:17
								illegal_insn_o = 1'b1;
						end
						6'b110010: begin
							// Trace: design.sv:12008:15
							alu_operator_o = sv2v_cast_C07C4(7'b0111011);
							// Trace: design.sv:12009:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12010:15
							regc_used_o = 1'b1;
							// Trace: design.sv:12011:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:12012:15
							scalar_replication_o = 1'b0;
							// Trace: design.sv:12013:15
							if (!((instr_rdata_i[14:12] == 3'b000) || (instr_rdata_i[14:12] == 3'b001)))
								// Trace: design.sv:12014:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[25] != 1'b0)
								// Trace: design.sv:12017:17
								illegal_insn_o = 1'b1;
						end
						6'b110100: begin
							// Trace: design.sv:12021:15
							alu_operator_o = (instr_rdata_i[25] ? sv2v_cast_C07C4(7'b0111001) : sv2v_cast_C07C4(7'b0111000));
							// Trace: design.sv:12022:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12023:15
							if (instr_rdata_i[14:12] != 3'b000)
								// Trace: design.sv:12024:17
								illegal_insn_o = 1'b1;
						end
						6'b110110: begin
							// Trace: design.sv:12028:15
							alu_operator_o = sv2v_cast_C07C4(7'b0111001);
							// Trace: design.sv:12029:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12030:15
							regc_used_o = 1'b1;
							// Trace: design.sv:12031:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:12032:15
							if (instr_rdata_i[14:12] != 3'b001)
								// Trace: design.sv:12033:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[25] != 1'b0)
								// Trace: design.sv:12036:17
								illegal_insn_o = 1'b1;
						end
						6'b111000: begin
							// Trace: design.sv:12040:15
							alu_operator_o = sv2v_cast_C07C4(7'b0111000);
							// Trace: design.sv:12041:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12042:15
							regc_used_o = 1'b1;
							// Trace: design.sv:12043:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:12044:15
							if (instr_rdata_i[14:12] != 3'b001)
								// Trace: design.sv:12045:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[25] != 1'b0)
								// Trace: design.sv:12048:17
								illegal_insn_o = 1'b1;
						end
						6'b011110: begin
							// Trace: design.sv:12052:15
							alu_operator_o = sv2v_cast_C07C4(7'b0111110);
							// Trace: design.sv:12053:15
							if (!((instr_rdata_i[14:12] == 3'b110) || (instr_rdata_i[14:12] == 3'b111)))
								// Trace: design.sv:12054:17
								illegal_insn_o = 1'b1;
						end
						6'b100100: begin
							// Trace: design.sv:12058:15
							alu_operator_o = sv2v_cast_C07C4(7'b0111111);
							// Trace: design.sv:12059:15
							if (!((instr_rdata_i[14:12] == 3'b110) || (instr_rdata_i[14:12] == 3'b111)))
								// Trace: design.sv:12060:17
								illegal_insn_o = 1'b1;
						end
						6'b101100: begin
							// Trace: design.sv:12064:15
							alu_operator_o = sv2v_cast_C07C4(7'b0101101);
							// Trace: design.sv:12065:15
							regc_used_o = 1'b1;
							// Trace: design.sv:12066:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:12067:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGC_OR_FWD;
							// Trace: design.sv:12068:15
							if (!((instr_rdata_i[14:12] == 3'b110) || (instr_rdata_i[14:12] == 3'b111)))
								// Trace: design.sv:12069:17
								illegal_insn_o = 1'b1;
						end
						6'b100000: begin
							// Trace: design.sv:12073:15
							alu_en = 1'b0;
							// Trace: design.sv:12074:15
							mult_dot_en = 1'b1;
							// Trace: design.sv:12075:15
							mult_dot_signed_o = 2'b00;
							// Trace: design.sv:12076:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:12077:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12078:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12081:17
								illegal_insn_o = 1'b1;
						end
						6'b100010: begin
							// Trace: design.sv:12085:15
							alu_en = 1'b0;
							// Trace: design.sv:12086:15
							mult_dot_en = 1'b1;
							// Trace: design.sv:12087:15
							mult_dot_signed_o = 2'b01;
							// Trace: design.sv:12088:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12089:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12092:17
								illegal_insn_o = 1'b1;
						end
						6'b100110: begin
							// Trace: design.sv:12096:15
							alu_en = 1'b0;
							// Trace: design.sv:12097:15
							mult_dot_en = 1'b1;
							// Trace: design.sv:12098:15
							mult_dot_signed_o = 2'b11;
							// Trace: design.sv:12099:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12100:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12103:17
								illegal_insn_o = 1'b1;
						end
						6'b101000: begin
							// Trace: design.sv:12107:15
							alu_en = 1'b0;
							// Trace: design.sv:12108:15
							mult_dot_en = 1'b1;
							// Trace: design.sv:12109:15
							mult_dot_signed_o = 2'b00;
							// Trace: design.sv:12110:15
							regc_used_o = 1'b1;
							// Trace: design.sv:12111:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:12112:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:12113:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12114:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12117:17
								illegal_insn_o = 1'b1;
						end
						6'b101010: begin
							// Trace: design.sv:12121:15
							alu_en = 1'b0;
							// Trace: design.sv:12122:15
							mult_dot_en = 1'b1;
							// Trace: design.sv:12123:15
							mult_dot_signed_o = 2'b01;
							// Trace: design.sv:12124:15
							regc_used_o = 1'b1;
							// Trace: design.sv:12125:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:12126:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12127:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12130:17
								illegal_insn_o = 1'b1;
						end
						6'b101110: begin
							// Trace: design.sv:12134:15
							alu_en = 1'b0;
							// Trace: design.sv:12135:15
							mult_dot_en = 1'b1;
							// Trace: design.sv:12136:15
							mult_dot_signed_o = 2'b11;
							// Trace: design.sv:12137:15
							regc_used_o = 1'b1;
							// Trace: design.sv:12138:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:12139:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12140:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12143:17
								illegal_insn_o = 1'b1;
						end
						6'b010101: begin
							// Trace: design.sv:12150:15
							alu_en = 1'b0;
							// Trace: design.sv:12151:15
							mult_dot_en = 1'b1;
							// Trace: design.sv:12152:15
							mult_dot_signed_o = 2'b11;
							// Trace: design.sv:12153:15
							is_clpx_o = 1'b1;
							// Trace: design.sv:12154:15
							regc_used_o = 1'b1;
							// Trace: design.sv:12155:15
							regc_mux_o = cv32e40p_pkg_REGC_RD;
							// Trace: design.sv:12156:15
							scalar_replication_o = 1'b0;
							// Trace: design.sv:12157:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGB_OR_FWD;
							// Trace: design.sv:12158:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12159:15
							illegal_insn_o = instr_rdata_i[12];
						end
						6'b011011: begin
							// Trace: design.sv:12163:15
							alu_operator_o = sv2v_cast_C07C4(7'b0011001);
							// Trace: design.sv:12164:15
							is_clpx_o = 1'b1;
							// Trace: design.sv:12165:15
							scalar_replication_o = 1'b0;
							// Trace: design.sv:12166:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGB_OR_FWD;
							// Trace: design.sv:12167:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12168:15
							is_subrot_o = 1'b1;
							// Trace: design.sv:12169:15
							if ((instr_rdata_i[25] != 1'b0) || (instr_rdata_i[12] != 1'b0))
								// Trace: design.sv:12170:17
								illegal_insn_o = 1'b1;
						end
						6'b010111: begin
							// Trace: design.sv:12175:15
							alu_operator_o = sv2v_cast_C07C4(7'b0010100);
							// Trace: design.sv:12176:15
							is_clpx_o = 1'b1;
							// Trace: design.sv:12177:15
							scalar_replication_o = 1'b0;
							// Trace: design.sv:12178:15
							regb_used_o = 1'b0;
							// Trace: design.sv:12179:15
							if (instr_rdata_i[14:12] != 3'b000)
								// Trace: design.sv:12180:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[25:20] != 6'b000000)
								// Trace: design.sv:12183:17
								illegal_insn_o = 1'b1;
						end
						6'b011101: begin
							// Trace: design.sv:12188:15
							alu_operator_o = sv2v_cast_C07C4(7'b0011000);
							// Trace: design.sv:12189:15
							is_clpx_o = 1'b1;
							// Trace: design.sv:12190:15
							scalar_replication_o = 1'b0;
							// Trace: design.sv:12191:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGB_OR_FWD;
							// Trace: design.sv:12192:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12193:15
							if (!(((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b100)) || (instr_rdata_i[14:12] == 3'b110)))
								// Trace: design.sv:12194:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[25] != 1'b0)
								// Trace: design.sv:12197:17
								illegal_insn_o = 1'b1;
						end
						6'b011001: begin
							// Trace: design.sv:12202:15
							alu_operator_o = sv2v_cast_C07C4(7'b0011001);
							// Trace: design.sv:12203:15
							is_clpx_o = 1'b1;
							// Trace: design.sv:12204:15
							scalar_replication_o = 1'b0;
							// Trace: design.sv:12205:15
							alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_REGB_OR_FWD;
							// Trace: design.sv:12206:15
							regb_used_o = 1'b1;
							// Trace: design.sv:12207:15
							if (!(((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b100)) || (instr_rdata_i[14:12] == 3'b110)))
								// Trace: design.sv:12208:17
								illegal_insn_o = 1'b1;
							if (instr_rdata_i[25] != 1'b0)
								// Trace: design.sv:12211:17
								illegal_insn_o = 1'b1;
						end
						6'b000001: begin
							// Trace: design.sv:12217:15
							alu_operator_o = sv2v_cast_C07C4(7'b0001100);
							// Trace: design.sv:12218:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:12219:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12220:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12223:17
								illegal_insn_o = 1'b1;
						end
						6'b000011: begin
							// Trace: design.sv:12227:15
							alu_operator_o = sv2v_cast_C07C4(7'b0001101);
							// Trace: design.sv:12228:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:12229:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12230:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12233:17
								illegal_insn_o = 1'b1;
						end
						6'b000101: begin
							// Trace: design.sv:12237:15
							alu_operator_o = sv2v_cast_C07C4(7'b0001000);
							// Trace: design.sv:12238:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:12239:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12240:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12243:17
								illegal_insn_o = 1'b1;
						end
						6'b000111: begin
							// Trace: design.sv:12247:15
							alu_operator_o = sv2v_cast_C07C4(7'b0001010);
							// Trace: design.sv:12248:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:12249:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12250:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12253:17
								illegal_insn_o = 1'b1;
						end
						6'b001001: begin
							// Trace: design.sv:12257:15
							alu_operator_o = sv2v_cast_C07C4(7'b0000000);
							// Trace: design.sv:12258:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:12259:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12260:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12263:17
								illegal_insn_o = 1'b1;
						end
						6'b001011: begin
							// Trace: design.sv:12267:15
							alu_operator_o = sv2v_cast_C07C4(7'b0000100);
							// Trace: design.sv:12268:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VS;
							// Trace: design.sv:12269:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12270:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12273:17
								illegal_insn_o = 1'b1;
						end
						6'b001101: begin
							// Trace: design.sv:12277:15
							alu_operator_o = sv2v_cast_C07C4(7'b0001001);
							// Trace: design.sv:12278:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:12279:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12280:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12283:17
								illegal_insn_o = 1'b1;
						end
						6'b001111: begin
							// Trace: design.sv:12287:15
							alu_operator_o = sv2v_cast_C07C4(7'b0001011);
							// Trace: design.sv:12288:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:12289:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12290:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12293:17
								illegal_insn_o = 1'b1;
						end
						6'b010001: begin
							// Trace: design.sv:12297:15
							alu_operator_o = sv2v_cast_C07C4(7'b0000001);
							// Trace: design.sv:12298:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:12299:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12300:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12303:17
								illegal_insn_o = 1'b1;
						end
						6'b010011: begin
							// Trace: design.sv:12307:15
							alu_operator_o = sv2v_cast_C07C4(7'b0000101);
							// Trace: design.sv:12308:15
							imm_b_mux_sel_o = cv32e40p_pkg_IMMB_VU;
							// Trace: design.sv:12309:15
							if ((instr_rdata_i[14:12] == 3'b010) || (instr_rdata_i[14:12] == 3'b011))
								// Trace: design.sv:12310:17
								illegal_insn_o = 1'b1;
							if (((instr_rdata_i[14:12] != 3'b110) && (instr_rdata_i[14:12] != 3'b111)) && (instr_rdata_i[25] != 1'b0))
								// Trace: design.sv:12313:17
								illegal_insn_o = 1'b1;
						end
						default:
							// Trace: design.sv:12317:22
							illegal_insn_o = 1'b1;
					endcase
				end
				else
					// Trace: design.sv:12320:11
					illegal_insn_o = 1'b1;
			cv32e40p_pkg_OPCODE_FENCE:
				// Trace: design.sv:12334:9
				(* full_case, parallel_case *)
				case (instr_rdata_i[14:12])
					3'b000:
						// Trace: design.sv:12337:13
						fencei_insn_o = 1'b1;
					3'b001:
						// Trace: design.sv:12342:13
						fencei_insn_o = 1'b1;
					default:
						// Trace: design.sv:12346:13
						illegal_insn_o = 1'b1;
				endcase
			cv32e40p_pkg_OPCODE_SYSTEM:
				// Trace: design.sv:12352:9
				if (instr_rdata_i[14:12] == 3'b000) begin
					begin
						// Trace: design.sv:12355:11
						if ({instr_rdata_i[19:15], instr_rdata_i[11:7]} == {10 {1'sb0}})
							// Trace: design.sv:12357:13
							(* full_case, parallel_case *)
							case (instr_rdata_i[31:20])
								12'h000:
									// Trace: design.sv:12361:17
									ecall_insn_o = 1'b1;
								12'h001:
									// Trace: design.sv:12367:17
									ebrk_insn_o = 1'b1;
								12'h302: begin
									// Trace: design.sv:12372:17
									illegal_insn_o = (PULP_SECURE ? current_priv_lvl_i != 2'b11 : 1'b0);
									// Trace: design.sv:12373:17
									mret_insn_o = ~illegal_insn_o;
									// Trace: design.sv:12374:17
									mret_dec_o = 1'b1;
								end
								12'h002: begin
									// Trace: design.sv:12379:17
									illegal_insn_o = (PULP_SECURE ? 1'b0 : 1'b1);
									// Trace: design.sv:12380:17
									uret_insn_o = ~illegal_insn_o;
									// Trace: design.sv:12381:17
									uret_dec_o = 1'b1;
								end
								12'h7b2: begin
									// Trace: design.sv:12386:17
									illegal_insn_o = !debug_mode_i;
									// Trace: design.sv:12387:17
									dret_insn_o = debug_mode_i;
									// Trace: design.sv:12388:17
									dret_dec_o = 1'b1;
								end
								12'h105: begin
									// Trace: design.sv:12393:17
									wfi_o = 1'b1;
									// Trace: design.sv:12394:17
									if (debug_wfi_no_sleep_i) begin
										// Trace: design.sv:12398:19
										alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
										// Trace: design.sv:12399:19
										imm_b_mux_sel_o = cv32e40p_pkg_IMMB_I;
										// Trace: design.sv:12400:19
										alu_operator_o = sv2v_cast_C07C4(7'b0011000);
									end
								end
								default:
									// Trace: design.sv:12406:17
									illegal_insn_o = 1'b1;
							endcase
						else
							// Trace: design.sv:12409:20
							illegal_insn_o = 1'b1;
					end
				end
				else begin
					// Trace: design.sv:12414:11
					csr_access_o = 1'b1;
					// Trace: design.sv:12415:11
					regfile_alu_we = 1'b1;
					// Trace: design.sv:12416:11
					alu_op_b_mux_sel_o = cv32e40p_pkg_OP_B_IMM;
					// Trace: design.sv:12417:11
					imm_a_mux_sel_o = cv32e40p_pkg_IMMA_Z;
					// Trace: design.sv:12418:11
					imm_b_mux_sel_o = cv32e40p_pkg_IMMB_I;
					// Trace: design.sv:12420:11
					if (instr_rdata_i[14] == 1'b1)
						// Trace: design.sv:12422:13
						alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_IMM;
					else begin
						// Trace: design.sv:12424:13
						rega_used_o = 1'b1;
						// Trace: design.sv:12425:13
						alu_op_a_mux_sel_o = cv32e40p_pkg_OP_A_REGA_OR_FWD;
					end
					(* full_case, parallel_case *)
					case (instr_rdata_i[13:12])
						2'b01:
							// Trace: design.sv:12432:22
							csr_op = sv2v_cast_EB06E(2'b01);
						2'b10:
							// Trace: design.sv:12433:22
							csr_op = (instr_rdata_i[19:15] == 5'b00000 ? sv2v_cast_EB06E(2'b00) : sv2v_cast_EB06E(2'b10));
						2'b11:
							// Trace: design.sv:12434:22
							csr_op = (instr_rdata_i[19:15] == 5'b00000 ? sv2v_cast_EB06E(2'b00) : sv2v_cast_EB06E(2'b11));
						default:
							// Trace: design.sv:12435:22
							csr_illegal = 1'b1;
					endcase
					if (instr_rdata_i[29:28] > current_priv_lvl_i)
						// Trace: design.sv:12440:13
						csr_illegal = 1'b1;
					case (instr_rdata_i[31:20])
						12'h001, 12'h002, 12'h003:
							if (!FPU)
								// Trace: design.sv:12449:26
								csr_illegal = 1'b1;
						12'hf11, 12'hf12, 12'hf13, 12'hf14:
							if (csr_op != sv2v_cast_EB06E(2'b00))
								// Trace: design.sv:12456:43
								csr_illegal = 1'b1;
						12'h300, 12'h341, 12'h305, 12'h342:
							// Trace: design.sv:12464:17
							csr_status_o = 1'b1;
						12'h301, 12'h304, 12'h340, 12'h343, 12'h344:
							;
						12'hb00, 12'hb02, 12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f, 12'hb80, 12'hb82, 12'hb83, 12'hb84, 12'hb85, 12'hb86, 12'hb87, 12'hb88, 12'hb89, 12'hb8a, 12'hb8b, 12'hb8c, 12'hb8d, 12'hb8e, 12'hb8f, 12'hb90, 12'hb91, 12'hb92, 12'hb93, 12'hb94, 12'hb95, 12'hb96, 12'hb97, 12'hb98, 12'hb99, 12'hb9a, 12'hb9b, 12'hb9c, 12'hb9d, 12'hb9e, 12'hb9f, 12'h320, 12'h323, 12'h324, 12'h325, 12'h326, 12'h327, 12'h328, 12'h329, 12'h32a, 12'h32b, 12'h32c, 12'h32d, 12'h32e, 12'h32f, 12'h330, 12'h331, 12'h332, 12'h333, 12'h334, 12'h335, 12'h336, 12'h337, 12'h338, 12'h339, 12'h33a, 12'h33b, 12'h33c, 12'h33d, 12'h33e, 12'h33f:
							// Trace: design.sv:12505:17
							csr_status_o = 1'b1;
						12'hc00, 12'hc02, 12'hc03, 12'hc04, 12'hc05, 12'hc06, 12'hc07, 12'hc08, 12'hc09, 12'hc0a, 12'hc0b, 12'hc0c, 12'hc0d, 12'hc0e, 12'hc0f, 12'hc10, 12'hc11, 12'hc12, 12'hc13, 12'hc14, 12'hc15, 12'hc16, 12'hc17, 12'hc18, 12'hc19, 12'hc1a, 12'hc1b, 12'hc1c, 12'hc1d, 12'hc1e, 12'hc1f, 12'hc80, 12'hc82, 12'hc83, 12'hc84, 12'hc85, 12'hc86, 12'hc87, 12'hc88, 12'hc89, 12'hc8a, 12'hc8b, 12'hc8c, 12'hc8d, 12'hc8e, 12'hc8f, 12'hc90, 12'hc91, 12'hc92, 12'hc93, 12'hc94, 12'hc95, 12'hc96, 12'hc97, 12'hc98, 12'hc99, 12'hc9a, 12'hc9b, 12'hc9c, 12'hc9d, 12'hc9e, 12'hc9f:
							if ((csr_op != sv2v_cast_EB06E(2'b00)) || ((PULP_SECURE && (current_priv_lvl_i != 2'b11)) && !mcounteren_i[instr_rdata_i[24:20]]))
								// Trace: design.sv:12530:19
								csr_illegal = 1'b1;
							else
								// Trace: design.sv:12532:19
								csr_status_o = 1'b1;
						12'h306:
							if (!PULP_SECURE)
								// Trace: design.sv:12538:17
								csr_illegal = 1'b1;
							else
								// Trace: design.sv:12540:17
								csr_status_o = 1'b1;
						12'h7b0, 12'h7b1, 12'h7b2, 12'h7b3:
							if (!debug_mode_i)
								// Trace: design.sv:12549:19
								csr_illegal = 1'b1;
							else
								// Trace: design.sv:12551:17
								csr_status_o = 1'b1;
						12'h7a0, 12'h7a1, 12'h7a2, 12'h7a3, 12'h7a4, 12'h7a8, 12'h7aa:
							if (DEBUG_TRIGGER_EN != 1)
								// Trace: design.sv:12563:19
								csr_illegal = 1'b1;
						12'h800, 12'h801, 12'h802, 12'h804, 12'h805, 12'h806, 12'hcc0:
							if (!PULP_XPULP)
								// Trace: design.sv:12573:33
								csr_illegal = 1'b1;
						12'hcc1:
							if (!PULP_XPULP)
								// Trace: design.sv:12578:17
								csr_illegal = 1'b1;
							else
								// Trace: design.sv:12580:17
								csr_status_o = 1'b1;
						12'h3a0, 12'h3a1, 12'h3a2, 12'h3a3, 12'h3b0, 12'h3b1, 12'h3b2, 12'h3b3, 12'h3b4, 12'h3b5, 12'h3b6, 12'h3b7, 12'h3b8, 12'h3b9, 12'h3ba, 12'h3bb, 12'h3bc, 12'h3bd, 12'h3be, 12'h3bf:
							if (!USE_PMP)
								// Trace: design.sv:12604:30
								csr_illegal = 1'b1;
						12'h000, 12'h041, 12'h005, 12'h042:
							if (!PULP_SECURE)
								// Trace: design.sv:12612:19
								csr_illegal = 1'b1;
							else
								// Trace: design.sv:12614:19
								csr_status_o = 1'b1;
						default:
							// Trace: design.sv:12617:23
							csr_illegal = 1'b1;
					endcase
					// Trace: design.sv:12621:11
					illegal_insn_o = csr_illegal;
				end
			cv32e40p_pkg_OPCODE_HWLOOP:
				// Trace: design.sv:12638:9
				if (PULP_XPULP) begin : HWLOOP_FEATURE_ENABLED
					// Trace: design.sv:12639:11
					hwlp_target_mux_sel_o = 1'b0;
					// Trace: design.sv:12641:11
					(* full_case, parallel_case *)
					case (instr_rdata_i[14:12])
						3'b000: begin
							// Trace: design.sv:12644:15
							hwlp_we[0] = 1'b1;
							// Trace: design.sv:12645:15
							hwlp_start_mux_sel_o = 1'b0;
							// Trace: design.sv:12646:15
							if (instr_rdata_i[19:15] != 5'b00000)
								// Trace: design.sv:12647:17
								illegal_insn_o = 1'b1;
						end
						3'b001: begin
							// Trace: design.sv:12653:15
							hwlp_we[1] = 1'b1;
							// Trace: design.sv:12654:15
							if (instr_rdata_i[19:15] != 5'b00000)
								// Trace: design.sv:12655:17
								illegal_insn_o = 1'b1;
						end
						3'b010: begin
							// Trace: design.sv:12661:15
							hwlp_we[2] = 1'b1;
							// Trace: design.sv:12662:15
							hwlp_cnt_mux_sel_o = 1'b1;
							// Trace: design.sv:12663:15
							rega_used_o = 1'b1;
							// Trace: design.sv:12664:15
							if (instr_rdata_i[31:20] != 12'b000000000000)
								// Trace: design.sv:12665:17
								illegal_insn_o = 1'b1;
						end
						3'b011: begin
							// Trace: design.sv:12671:15
							hwlp_we[2] = 1'b1;
							// Trace: design.sv:12672:15
							hwlp_cnt_mux_sel_o = 1'b0;
							// Trace: design.sv:12673:15
							if (instr_rdata_i[19:15] != 5'b00000)
								// Trace: design.sv:12674:17
								illegal_insn_o = 1'b1;
						end
						3'b100: begin
							// Trace: design.sv:12681:15
							hwlp_we = 3'b111;
							// Trace: design.sv:12682:15
							hwlp_start_mux_sel_o = 1'b1;
							// Trace: design.sv:12683:15
							hwlp_cnt_mux_sel_o = 1'b1;
							// Trace: design.sv:12684:15
							rega_used_o = 1'b1;
						end
						3'b101: begin
							// Trace: design.sv:12690:15
							hwlp_we = 3'b111;
							// Trace: design.sv:12691:15
							hwlp_target_mux_sel_o = 1'b1;
							// Trace: design.sv:12692:15
							hwlp_start_mux_sel_o = 1'b1;
							// Trace: design.sv:12693:15
							hwlp_cnt_mux_sel_o = 1'b0;
						end
						default:
							// Trace: design.sv:12697:15
							illegal_insn_o = 1'b1;
					endcase
					if (instr_rdata_i[11:8] != 4'b0000)
						// Trace: design.sv:12702:13
						illegal_insn_o = 1'b1;
				end
				else
					// Trace: design.sv:12708:11
					illegal_insn_o = 1'b1;
			default:
				// Trace: design.sv:12713:9
				illegal_insn_o = 1'b1;
		endcase
		if (illegal_c_insn_i)
			// Trace: design.sv:12720:7
			illegal_insn_o = 1'b1;
	end
	// Trace: design.sv:12726:3
	assign alu_en_o = (deassert_we_i ? 1'b0 : alu_en);
	// Trace: design.sv:12727:3
	assign apu_en_o = (deassert_we_i ? 1'b0 : apu_en);
	// Trace: design.sv:12728:3
	assign mult_int_en_o = (deassert_we_i ? 1'b0 : mult_int_en);
	// Trace: design.sv:12729:3
	assign mult_dot_en_o = (deassert_we_i ? 1'b0 : mult_dot_en);
	// Trace: design.sv:12730:3
	assign regfile_mem_we_o = (deassert_we_i ? 1'b0 : regfile_mem_we);
	// Trace: design.sv:12731:3
	assign regfile_alu_we_o = (deassert_we_i ? 1'b0 : regfile_alu_we);
	// Trace: design.sv:12732:3
	assign data_req_o = (deassert_we_i ? 1'b0 : data_req);
	// Trace: design.sv:12733:3
	assign hwlp_we_o = (deassert_we_i ? 3'b000 : hwlp_we);
	// Trace: design.sv:12734:3
	assign csr_op_o = (deassert_we_i ? sv2v_cast_EB06E(2'b00) : csr_op);
	// Trace: design.sv:12735:3
	assign ctrl_transfer_insn_in_id_o = (deassert_we_i ? cv32e40p_pkg_BRANCH_NONE : ctrl_transfer_insn);
	// Trace: design.sv:12737:3
	assign ctrl_transfer_insn_in_dec_o = ctrl_transfer_insn;
	// Trace: design.sv:12738:3
	assign regfile_alu_we_dec_o = regfile_alu_we;
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_int_controller (
	clk,
	rst_n,
	irq_i,
	irq_sec_i,
	irq_req_ctrl_o,
	irq_sec_ctrl_o,
	irq_id_ctrl_o,
	irq_wu_ctrl_o,
	mie_bypass_i,
	mip_o,
	m_ie_i,
	u_ie_i,
	current_priv_lvl_i
);
	reg _sv2v_0;
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:12767:15
	parameter PULP_SECURE = 0;
	// Trace: design.sv:12769:5
	input wire clk;
	// Trace: design.sv:12770:5
	input wire rst_n;
	// Trace: design.sv:12773:5
	input wire [31:0] irq_i;
	// Trace: design.sv:12774:5
	input wire irq_sec_i;
	// Trace: design.sv:12777:5
	output wire irq_req_ctrl_o;
	// Trace: design.sv:12778:5
	output wire irq_sec_ctrl_o;
	// Trace: design.sv:12779:5
	output reg [4:0] irq_id_ctrl_o;
	// Trace: design.sv:12780:5
	output wire irq_wu_ctrl_o;
	// Trace: design.sv:12783:5
	input wire [31:0] mie_bypass_i;
	// Trace: design.sv:12784:5
	output wire [31:0] mip_o;
	// Trace: design.sv:12785:5
	input wire m_ie_i;
	// Trace: design.sv:12786:5
	input wire u_ie_i;
	// Trace: design.sv:12787:5
	// removed localparam type cv32e40p_pkg_PrivLvl_t
	input wire [1:0] current_priv_lvl_i;
	// Trace: design.sv:12790:3
	wire global_irq_enable;
	// Trace: design.sv:12791:3
	wire [31:0] irq_local_qual;
	// Trace: design.sv:12792:3
	reg [31:0] irq_q;
	// Trace: design.sv:12793:3
	reg irq_sec_q;
	// Trace: design.sv:12799:3
	localparam cv32e40p_pkg_IRQ_MASK = 32'hffff0888;
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:12800:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:12801:7
			irq_q <= 1'sb0;
			// Trace: design.sv:12802:7
			irq_sec_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:12804:7
			irq_q <= irq_i & cv32e40p_pkg_IRQ_MASK;
			// Trace: design.sv:12805:7
			irq_sec_q <= irq_sec_i;
		end
	// Trace: design.sv:12810:3
	assign mip_o = irq_q;
	// Trace: design.sv:12813:3
	assign irq_local_qual = irq_q & mie_bypass_i;
	// Trace: design.sv:12816:3
	assign irq_wu_ctrl_o = |(irq_i & mie_bypass_i);
	// Trace: design.sv:12819:3
	generate
		if (PULP_SECURE) begin : gen_pulp_secure
			// Trace: design.sv:12821:7
			assign global_irq_enable = ((u_ie_i || irq_sec_i) && (current_priv_lvl_i == 2'b00)) || (m_ie_i && (current_priv_lvl_i == 2'b11));
		end
		else begin : gen_no_pulp_secure
			// Trace: design.sv:12823:7
			assign global_irq_enable = m_ie_i;
		end
	endgenerate
	// Trace: design.sv:12828:3
	assign irq_req_ctrl_o = |irq_local_qual && global_irq_enable;
	// Trace: design.sv:12835:3
	localparam [31:0] cv32e40p_pkg_CSR_MEIX_BIT = 11;
	localparam [31:0] cv32e40p_pkg_CSR_MSIX_BIT = 3;
	localparam [31:0] cv32e40p_pkg_CSR_MTIX_BIT = 7;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:12836:5
		if (irq_local_qual[31])
			// Trace: design.sv:12836:29
			irq_id_ctrl_o = 5'd31;
		else if (irq_local_qual[30])
			// Trace: design.sv:12837:34
			irq_id_ctrl_o = 5'd30;
		else if (irq_local_qual[29])
			// Trace: design.sv:12838:34
			irq_id_ctrl_o = 5'd29;
		else if (irq_local_qual[28])
			// Trace: design.sv:12839:34
			irq_id_ctrl_o = 5'd28;
		else if (irq_local_qual[27])
			// Trace: design.sv:12840:34
			irq_id_ctrl_o = 5'd27;
		else if (irq_local_qual[26])
			// Trace: design.sv:12841:34
			irq_id_ctrl_o = 5'd26;
		else if (irq_local_qual[25])
			// Trace: design.sv:12842:34
			irq_id_ctrl_o = 5'd25;
		else if (irq_local_qual[24])
			// Trace: design.sv:12843:34
			irq_id_ctrl_o = 5'd24;
		else if (irq_local_qual[23])
			// Trace: design.sv:12844:34
			irq_id_ctrl_o = 5'd23;
		else if (irq_local_qual[22])
			// Trace: design.sv:12845:34
			irq_id_ctrl_o = 5'd22;
		else if (irq_local_qual[21])
			// Trace: design.sv:12846:34
			irq_id_ctrl_o = 5'd21;
		else if (irq_local_qual[20])
			// Trace: design.sv:12847:34
			irq_id_ctrl_o = 5'd20;
		else if (irq_local_qual[19])
			// Trace: design.sv:12848:34
			irq_id_ctrl_o = 5'd19;
		else if (irq_local_qual[18])
			// Trace: design.sv:12849:34
			irq_id_ctrl_o = 5'd18;
		else if (irq_local_qual[17])
			// Trace: design.sv:12850:34
			irq_id_ctrl_o = 5'd17;
		else if (irq_local_qual[16])
			// Trace: design.sv:12851:34
			irq_id_ctrl_o = 5'd16;
		else if (irq_local_qual[15])
			// Trace: design.sv:12854:7
			irq_id_ctrl_o = 5'd15;
		else if (irq_local_qual[14])
			// Trace: design.sv:12856:7
			irq_id_ctrl_o = 5'd14;
		else if (irq_local_qual[13])
			// Trace: design.sv:12858:7
			irq_id_ctrl_o = 5'd13;
		else if (irq_local_qual[12])
			// Trace: design.sv:12860:7
			irq_id_ctrl_o = 5'd12;
		else if (irq_local_qual[cv32e40p_pkg_CSR_MEIX_BIT])
			// Trace: design.sv:12862:44
			irq_id_ctrl_o = cv32e40p_pkg_CSR_MEIX_BIT;
		else if (irq_local_qual[cv32e40p_pkg_CSR_MSIX_BIT])
			// Trace: design.sv:12863:44
			irq_id_ctrl_o = cv32e40p_pkg_CSR_MSIX_BIT;
		else if (irq_local_qual[cv32e40p_pkg_CSR_MTIX_BIT])
			// Trace: design.sv:12864:44
			irq_id_ctrl_o = cv32e40p_pkg_CSR_MTIX_BIT;
		else if (irq_local_qual[10])
			// Trace: design.sv:12867:7
			irq_id_ctrl_o = 5'd10;
		else if (irq_local_qual[2])
			// Trace: design.sv:12869:7
			irq_id_ctrl_o = 5'd2;
		else if (irq_local_qual[6])
			// Trace: design.sv:12871:7
			irq_id_ctrl_o = 5'd6;
		else if (irq_local_qual[9])
			// Trace: design.sv:12874:7
			irq_id_ctrl_o = 5'd9;
		else if (irq_local_qual[1])
			// Trace: design.sv:12876:7
			irq_id_ctrl_o = 5'd1;
		else if (irq_local_qual[5])
			// Trace: design.sv:12878:7
			irq_id_ctrl_o = 5'd5;
		else if (irq_local_qual[8])
			// Trace: design.sv:12881:7
			irq_id_ctrl_o = 5'd8;
		else if (irq_local_qual[0])
			// Trace: design.sv:12883:7
			irq_id_ctrl_o = 5'd0;
		else if (irq_local_qual[4])
			// Trace: design.sv:12885:7
			irq_id_ctrl_o = 5'd4;
		else
			// Trace: design.sv:12887:10
			irq_id_ctrl_o = cv32e40p_pkg_CSR_MTIX_BIT;
	end
	// Trace: design.sv:12890:3
	assign irq_sec_ctrl_o = irq_sec_q;
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_ex_stage (
	clk,
	rst_n,
	alu_operator_i,
	alu_operand_a_i,
	alu_operand_b_i,
	alu_operand_c_i,
	alu_en_i,
	bmask_a_i,
	bmask_b_i,
	imm_vec_ext_i,
	alu_vec_mode_i,
	alu_is_clpx_i,
	alu_is_subrot_i,
	alu_clpx_shift_i,
	mult_operator_i,
	mult_operand_a_i,
	mult_operand_b_i,
	mult_operand_c_i,
	mult_en_i,
	mult_sel_subword_i,
	mult_signed_mode_i,
	mult_imm_i,
	mult_dot_op_a_i,
	mult_dot_op_b_i,
	mult_dot_op_c_i,
	mult_dot_signed_i,
	mult_is_clpx_i,
	mult_clpx_shift_i,
	mult_clpx_img_i,
	mult_multicycle_o,
	fpu_fflags_we_o,
	apu_en_i,
	apu_op_i,
	apu_lat_i,
	apu_operands_i,
	apu_waddr_i,
	apu_flags_i,
	apu_read_regs_i,
	apu_read_regs_valid_i,
	apu_read_dep_o,
	apu_write_regs_i,
	apu_write_regs_valid_i,
	apu_write_dep_o,
	apu_perf_type_o,
	apu_perf_cont_o,
	apu_perf_wb_o,
	apu_busy_o,
	apu_ready_wb_o,
	apu_req_o,
	apu_gnt_i,
	apu_operands_o,
	apu_op_o,
	apu_rvalid_i,
	apu_result_i,
	lsu_en_i,
	lsu_rdata_i,
	branch_in_ex_i,
	regfile_alu_waddr_i,
	regfile_alu_we_i,
	regfile_we_i,
	regfile_waddr_i,
	csr_access_i,
	csr_rdata_i,
	regfile_waddr_wb_o,
	regfile_we_wb_o,
	regfile_wdata_wb_o,
	regfile_alu_waddr_fw_o,
	regfile_alu_we_fw_o,
	regfile_alu_wdata_fw_o,
	jump_target_o,
	branch_decision_o,
	is_decoding_i,
	lsu_ready_ex_i,
	lsu_err_i,
	ex_ready_o,
	ex_valid_o,
	wb_ready_i
);
	reg _sv2v_0;
	// removed import cv32e40p_pkg::*;
	// removed import cv32e40p_apu_core_pkg::*;
	// Trace: design.sv:12928:15
	parameter FPU = 0;
	// Trace: design.sv:12929:15
	parameter APU_NARGS_CPU = 3;
	// Trace: design.sv:12930:15
	parameter APU_WOP_CPU = 6;
	// Trace: design.sv:12931:15
	parameter APU_NDSFLAGS_CPU = 15;
	// Trace: design.sv:12932:15
	parameter APU_NUSFLAGS_CPU = 5;
	// Trace: design.sv:12934:5
	input wire clk;
	// Trace: design.sv:12935:5
	input wire rst_n;
	// Trace: design.sv:12938:5
	localparam cv32e40p_pkg_ALU_OP_WIDTH = 7;
	// removed localparam type cv32e40p_pkg_alu_opcode_e
	input wire [6:0] alu_operator_i;
	// Trace: design.sv:12939:5
	input wire [31:0] alu_operand_a_i;
	// Trace: design.sv:12940:5
	input wire [31:0] alu_operand_b_i;
	// Trace: design.sv:12941:5
	input wire [31:0] alu_operand_c_i;
	// Trace: design.sv:12942:5
	input wire alu_en_i;
	// Trace: design.sv:12943:5
	input wire [4:0] bmask_a_i;
	// Trace: design.sv:12944:5
	input wire [4:0] bmask_b_i;
	// Trace: design.sv:12945:5
	input wire [1:0] imm_vec_ext_i;
	// Trace: design.sv:12946:5
	input wire [1:0] alu_vec_mode_i;
	// Trace: design.sv:12947:5
	input wire alu_is_clpx_i;
	// Trace: design.sv:12948:5
	input wire alu_is_subrot_i;
	// Trace: design.sv:12949:5
	input wire [1:0] alu_clpx_shift_i;
	// Trace: design.sv:12952:5
	localparam cv32e40p_pkg_MUL_OP_WIDTH = 3;
	// removed localparam type cv32e40p_pkg_mul_opcode_e
	input wire [2:0] mult_operator_i;
	// Trace: design.sv:12953:5
	input wire [31:0] mult_operand_a_i;
	// Trace: design.sv:12954:5
	input wire [31:0] mult_operand_b_i;
	// Trace: design.sv:12955:5
	input wire [31:0] mult_operand_c_i;
	// Trace: design.sv:12956:5
	input wire mult_en_i;
	// Trace: design.sv:12957:5
	input wire mult_sel_subword_i;
	// Trace: design.sv:12958:5
	input wire [1:0] mult_signed_mode_i;
	// Trace: design.sv:12959:5
	input wire [4:0] mult_imm_i;
	// Trace: design.sv:12961:5
	input wire [31:0] mult_dot_op_a_i;
	// Trace: design.sv:12962:5
	input wire [31:0] mult_dot_op_b_i;
	// Trace: design.sv:12963:5
	input wire [31:0] mult_dot_op_c_i;
	// Trace: design.sv:12964:5
	input wire [1:0] mult_dot_signed_i;
	// Trace: design.sv:12965:5
	input wire mult_is_clpx_i;
	// Trace: design.sv:12966:5
	input wire [1:0] mult_clpx_shift_i;
	// Trace: design.sv:12967:5
	input wire mult_clpx_img_i;
	// Trace: design.sv:12969:5
	output wire mult_multicycle_o;
	// Trace: design.sv:12972:5
	output wire fpu_fflags_we_o;
	// Trace: design.sv:12975:5
	input wire apu_en_i;
	// Trace: design.sv:12976:5
	input wire [APU_WOP_CPU - 1:0] apu_op_i;
	// Trace: design.sv:12977:5
	input wire [1:0] apu_lat_i;
	// Trace: design.sv:12978:5
	input wire [(APU_NARGS_CPU * 32) - 1:0] apu_operands_i;
	// Trace: design.sv:12979:5
	input wire [5:0] apu_waddr_i;
	// Trace: design.sv:12980:5
	input wire [APU_NDSFLAGS_CPU - 1:0] apu_flags_i;
	// Trace: design.sv:12982:5
	input wire [17:0] apu_read_regs_i;
	// Trace: design.sv:12983:5
	input wire [2:0] apu_read_regs_valid_i;
	// Trace: design.sv:12984:5
	output wire apu_read_dep_o;
	// Trace: design.sv:12985:5
	input wire [11:0] apu_write_regs_i;
	// Trace: design.sv:12986:5
	input wire [1:0] apu_write_regs_valid_i;
	// Trace: design.sv:12987:5
	output wire apu_write_dep_o;
	// Trace: design.sv:12989:5
	output wire apu_perf_type_o;
	// Trace: design.sv:12990:5
	output wire apu_perf_cont_o;
	// Trace: design.sv:12991:5
	output wire apu_perf_wb_o;
	// Trace: design.sv:12993:5
	output wire apu_busy_o;
	// Trace: design.sv:12994:5
	output wire apu_ready_wb_o;
	// Trace: design.sv:12998:5
	output wire apu_req_o;
	// Trace: design.sv:12999:5
	input wire apu_gnt_i;
	// Trace: design.sv:13001:5
	output wire [(APU_NARGS_CPU * 32) - 1:0] apu_operands_o;
	// Trace: design.sv:13002:5
	output wire [APU_WOP_CPU - 1:0] apu_op_o;
	// Trace: design.sv:13004:5
	input wire apu_rvalid_i;
	// Trace: design.sv:13005:5
	input wire [31:0] apu_result_i;
	// Trace: design.sv:13007:5
	input wire lsu_en_i;
	// Trace: design.sv:13008:5
	input wire [31:0] lsu_rdata_i;
	// Trace: design.sv:13011:5
	input wire branch_in_ex_i;
	// Trace: design.sv:13012:5
	input wire [5:0] regfile_alu_waddr_i;
	// Trace: design.sv:13013:5
	input wire regfile_alu_we_i;
	// Trace: design.sv:13016:5
	input wire regfile_we_i;
	// Trace: design.sv:13017:5
	input wire [5:0] regfile_waddr_i;
	// Trace: design.sv:13020:5
	input wire csr_access_i;
	// Trace: design.sv:13021:5
	input wire [31:0] csr_rdata_i;
	// Trace: design.sv:13024:5
	output reg [5:0] regfile_waddr_wb_o;
	// Trace: design.sv:13025:5
	output reg regfile_we_wb_o;
	// Trace: design.sv:13026:5
	output reg [31:0] regfile_wdata_wb_o;
	// Trace: design.sv:13029:5
	output reg [5:0] regfile_alu_waddr_fw_o;
	// Trace: design.sv:13030:5
	output reg regfile_alu_we_fw_o;
	// Trace: design.sv:13031:5
	output reg [31:0] regfile_alu_wdata_fw_o;
	// Trace: design.sv:13034:5
	output wire [31:0] jump_target_o;
	// Trace: design.sv:13035:5
	output wire branch_decision_o;
	// Trace: design.sv:13038:5
	input wire is_decoding_i;
	// Trace: design.sv:13039:5
	input wire lsu_ready_ex_i;
	// Trace: design.sv:13040:5
	input wire lsu_err_i;
	// Trace: design.sv:13042:5
	output wire ex_ready_o;
	// Trace: design.sv:13043:5
	output wire ex_valid_o;
	// Trace: design.sv:13044:5
	input wire wb_ready_i;
	// Trace: design.sv:13047:3
	wire [31:0] alu_result;
	// Trace: design.sv:13048:3
	wire [31:0] mult_result;
	// Trace: design.sv:13049:3
	wire alu_cmp_result;
	// Trace: design.sv:13051:3
	reg regfile_we_lsu;
	// Trace: design.sv:13052:3
	reg [5:0] regfile_waddr_lsu;
	// Trace: design.sv:13054:3
	reg wb_contention;
	// Trace: design.sv:13055:3
	reg wb_contention_lsu;
	// Trace: design.sv:13057:3
	wire alu_ready;
	// Trace: design.sv:13058:3
	wire mult_ready;
	// Trace: design.sv:13061:3
	wire apu_valid;
	// Trace: design.sv:13062:3
	wire [5:0] apu_waddr;
	// Trace: design.sv:13063:3
	wire [31:0] apu_result;
	// Trace: design.sv:13064:3
	wire apu_stall;
	// Trace: design.sv:13065:3
	wire apu_active;
	// Trace: design.sv:13066:3
	wire apu_singlecycle;
	// Trace: design.sv:13067:3
	wire apu_multicycle;
	// Trace: design.sv:13068:3
	wire apu_req;
	// Trace: design.sv:13069:3
	wire apu_gnt;
	// Trace: design.sv:13072:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:13073:5
		regfile_alu_wdata_fw_o = 1'sb0;
		// Trace: design.sv:13074:5
		regfile_alu_waddr_fw_o = 1'sb0;
		// Trace: design.sv:13075:5
		regfile_alu_we_fw_o = 1'sb0;
		// Trace: design.sv:13076:5
		wb_contention = 1'b0;
		// Trace: design.sv:13079:5
		if (apu_valid & (apu_singlecycle | apu_multicycle)) begin
			// Trace: design.sv:13080:7
			regfile_alu_we_fw_o = 1'b1;
			// Trace: design.sv:13081:7
			regfile_alu_waddr_fw_o = apu_waddr;
			// Trace: design.sv:13082:7
			regfile_alu_wdata_fw_o = apu_result;
			// Trace: design.sv:13084:7
			if (regfile_alu_we_i & ~apu_en_i)
				// Trace: design.sv:13085:9
				wb_contention = 1'b1;
		end
		else begin
			// Trace: design.sv:13088:7
			regfile_alu_we_fw_o = regfile_alu_we_i & ~apu_en_i;
			// Trace: design.sv:13089:7
			regfile_alu_waddr_fw_o = regfile_alu_waddr_i;
			// Trace: design.sv:13090:7
			if (alu_en_i)
				// Trace: design.sv:13090:21
				regfile_alu_wdata_fw_o = alu_result;
			if (mult_en_i)
				// Trace: design.sv:13091:22
				regfile_alu_wdata_fw_o = mult_result;
			if (csr_access_i)
				// Trace: design.sv:13092:25
				regfile_alu_wdata_fw_o = csr_rdata_i;
		end
	end
	// Trace: design.sv:13097:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:13098:5
		regfile_we_wb_o = 1'b0;
		// Trace: design.sv:13099:5
		regfile_waddr_wb_o = regfile_waddr_lsu;
		// Trace: design.sv:13100:5
		regfile_wdata_wb_o = lsu_rdata_i;
		// Trace: design.sv:13101:5
		wb_contention_lsu = 1'b0;
		// Trace: design.sv:13103:5
		if (regfile_we_lsu) begin
			// Trace: design.sv:13104:7
			regfile_we_wb_o = 1'b1;
			// Trace: design.sv:13105:7
			if (apu_valid & (!apu_singlecycle & !apu_multicycle))
				// Trace: design.sv:13106:9
				wb_contention_lsu = 1'b1;
		end
		else if (apu_valid & (!apu_singlecycle & !apu_multicycle)) begin
			// Trace: design.sv:13110:7
			regfile_we_wb_o = 1'b1;
			// Trace: design.sv:13111:7
			regfile_waddr_wb_o = apu_waddr;
			// Trace: design.sv:13112:7
			regfile_wdata_wb_o = apu_result;
		end
	end
	// Trace: design.sv:13117:3
	assign branch_decision_o = alu_cmp_result;
	// Trace: design.sv:13118:3
	assign jump_target_o = alu_operand_c_i;
	// Trace: design.sv:13130:3
	cv32e40p_alu alu_i(
		.clk(clk),
		.rst_n(rst_n),
		.enable_i(alu_en_i),
		.operator_i(alu_operator_i),
		.operand_a_i(alu_operand_a_i),
		.operand_b_i(alu_operand_b_i),
		.operand_c_i(alu_operand_c_i),
		.vector_mode_i(alu_vec_mode_i),
		.bmask_a_i(bmask_a_i),
		.bmask_b_i(bmask_b_i),
		.imm_vec_ext_i(imm_vec_ext_i),
		.is_clpx_i(alu_is_clpx_i),
		.clpx_shift_i(alu_clpx_shift_i),
		.is_subrot_i(alu_is_subrot_i),
		.result_o(alu_result),
		.comparison_result_o(alu_cmp_result),
		.ready_o(alu_ready),
		.ex_ready_i(ex_ready_o)
	);
	// Trace: design.sv:13165:3
	cv32e40p_mult mult_i(
		.clk(clk),
		.rst_n(rst_n),
		.enable_i(mult_en_i),
		.operator_i(mult_operator_i),
		.short_subword_i(mult_sel_subword_i),
		.short_signed_i(mult_signed_mode_i),
		.op_a_i(mult_operand_a_i),
		.op_b_i(mult_operand_b_i),
		.op_c_i(mult_operand_c_i),
		.imm_i(mult_imm_i),
		.dot_op_a_i(mult_dot_op_a_i),
		.dot_op_b_i(mult_dot_op_b_i),
		.dot_op_c_i(mult_dot_op_c_i),
		.dot_signed_i(mult_dot_signed_i),
		.is_clpx_i(mult_is_clpx_i),
		.clpx_shift_i(mult_clpx_shift_i),
		.clpx_img_i(mult_clpx_img_i),
		.result_o(mult_result),
		.multicycle_o(mult_multicycle_o),
		.ready_o(mult_ready),
		.ex_ready_i(ex_ready_o)
	);
	// Trace: design.sv:13195:3
	generate
		if (FPU == 1) begin : gen_apu
			// Trace: design.sv:13206:7
			cv32e40p_apu_disp apu_disp_i(
				.clk_i(clk),
				.rst_ni(rst_n),
				.enable_i(apu_en_i),
				.apu_lat_i(apu_lat_i),
				.apu_waddr_i(apu_waddr_i),
				.apu_waddr_o(apu_waddr),
				.apu_multicycle_o(apu_multicycle),
				.apu_singlecycle_o(apu_singlecycle),
				.active_o(apu_active),
				.stall_o(apu_stall),
				.is_decoding_i(is_decoding_i),
				.read_regs_i(apu_read_regs_i),
				.read_regs_valid_i(apu_read_regs_valid_i),
				.read_dep_o(apu_read_dep_o),
				.write_regs_i(apu_write_regs_i),
				.write_regs_valid_i(apu_write_regs_valid_i),
				.write_dep_o(apu_write_dep_o),
				.perf_type_o(apu_perf_type_o),
				.perf_cont_o(apu_perf_cont_o),
				.apu_req_o(apu_req),
				.apu_gnt_i(apu_gnt),
				.apu_rvalid_i(apu_valid)
			);
			// Trace: design.sv:13240:7
			assign apu_perf_wb_o = wb_contention | wb_contention_lsu;
			// Trace: design.sv:13241:7
			assign apu_ready_wb_o = ~((apu_active | apu_en_i) | apu_stall) | apu_valid;
			// Trace: design.sv:13243:7
			assign apu_req_o = apu_req;
			// Trace: design.sv:13244:7
			assign apu_gnt = apu_gnt_i;
			// Trace: design.sv:13245:7
			assign apu_valid = apu_rvalid_i;
			// Trace: design.sv:13246:7
			assign apu_operands_o = apu_operands_i;
			// Trace: design.sv:13247:7
			assign apu_op_o = apu_op_i;
			// Trace: design.sv:13248:7
			assign apu_result = apu_result_i;
			// Trace: design.sv:13249:7
			assign fpu_fflags_we_o = apu_valid;
		end
		else begin : gen_no_apu
			// Trace: design.sv:13252:7
			assign apu_req_o = 1'sb0;
			// Trace: design.sv:13253:7
			assign apu_operands_o[0+:32] = 1'sb0;
			// Trace: design.sv:13254:7
			assign apu_operands_o[32+:32] = 1'sb0;
			// Trace: design.sv:13255:7
			assign apu_operands_o[64+:32] = 1'sb0;
			// Trace: design.sv:13256:7
			assign apu_op_o = 1'sb0;
			// Trace: design.sv:13257:7
			assign apu_req = 1'b0;
			// Trace: design.sv:13258:7
			assign apu_gnt = 1'b0;
			// Trace: design.sv:13259:7
			assign apu_result = 32'b00000000000000000000000000000000;
			// Trace: design.sv:13260:7
			assign apu_valid = 1'b0;
			// Trace: design.sv:13261:7
			assign apu_waddr = 6'b000000;
			// Trace: design.sv:13262:7
			assign apu_stall = 1'b0;
			// Trace: design.sv:13263:7
			assign apu_active = 1'b0;
			// Trace: design.sv:13264:7
			assign apu_ready_wb_o = 1'b1;
			// Trace: design.sv:13265:7
			assign apu_perf_wb_o = 1'b0;
			// Trace: design.sv:13266:7
			assign apu_perf_cont_o = 1'b0;
			// Trace: design.sv:13267:7
			assign apu_perf_type_o = 1'b0;
			// Trace: design.sv:13268:7
			assign apu_singlecycle = 1'b0;
			// Trace: design.sv:13269:7
			assign apu_multicycle = 1'b0;
			// Trace: design.sv:13270:7
			assign apu_read_dep_o = 1'b0;
			// Trace: design.sv:13271:7
			assign apu_write_dep_o = 1'b0;
			// Trace: design.sv:13272:7
			assign fpu_fflags_we_o = 1'b0;
		end
	endgenerate
	// Trace: design.sv:13277:3
	assign apu_busy_o = apu_active;
	// Trace: design.sv:13282:3
	always @(posedge clk or negedge rst_n) begin : EX_WB_Pipeline_Register
		// Trace: design.sv:13283:5
		if (~rst_n) begin
			// Trace: design.sv:13284:7
			regfile_waddr_lsu <= 1'sb0;
			// Trace: design.sv:13285:7
			regfile_we_lsu <= 1'b0;
		end
		else
			// Trace: design.sv:13287:7
			if (ex_valid_o) begin
				// Trace: design.sv:13289:9
				regfile_we_lsu <= regfile_we_i & ~lsu_err_i;
				// Trace: design.sv:13290:9
				if (regfile_we_i & ~lsu_err_i)
					// Trace: design.sv:13291:11
					regfile_waddr_lsu <= regfile_waddr_i;
			end
			else if (wb_ready_i)
				// Trace: design.sv:13296:9
				regfile_we_lsu <= 1'b0;
	end
	// Trace: design.sv:13304:3
	assign ex_ready_o = (((((~apu_stall & alu_ready) & mult_ready) & lsu_ready_ex_i) & wb_ready_i) & ~wb_contention) | branch_in_ex_i;
	// Trace: design.sv:13306:3
	assign ex_valid_o = ((((apu_valid | alu_en_i) | mult_en_i) | csr_access_i) | lsu_en_i) & (((alu_ready & mult_ready) & lsu_ready_ex_i) & wb_ready_i);
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_hwloop_regs (
	clk,
	rst_n,
	hwlp_start_data_i,
	hwlp_end_data_i,
	hwlp_cnt_data_i,
	hwlp_we_i,
	hwlp_regid_i,
	valid_i,
	hwlp_dec_cnt_i,
	hwlp_start_addr_o,
	hwlp_end_addr_o,
	hwlp_counter_o
);
	// Trace: design.sv:13335:15
	parameter N_REGS = 2;
	// Trace: design.sv:13336:15
	parameter N_REG_BITS = $clog2(N_REGS);
	// Trace: design.sv:13338:5
	input wire clk;
	// Trace: design.sv:13339:5
	input wire rst_n;
	// Trace: design.sv:13342:5
	input wire [31:0] hwlp_start_data_i;
	// Trace: design.sv:13343:5
	input wire [31:0] hwlp_end_data_i;
	// Trace: design.sv:13344:5
	input wire [31:0] hwlp_cnt_data_i;
	// Trace: design.sv:13345:5
	input wire [2:0] hwlp_we_i;
	// Trace: design.sv:13346:5
	input wire [N_REG_BITS - 1:0] hwlp_regid_i;
	// Trace: design.sv:13349:5
	input wire valid_i;
	// Trace: design.sv:13352:5
	input wire [N_REGS - 1:0] hwlp_dec_cnt_i;
	// Trace: design.sv:13355:5
	output wire [(N_REGS * 32) - 1:0] hwlp_start_addr_o;
	// Trace: design.sv:13356:5
	output wire [(N_REGS * 32) - 1:0] hwlp_end_addr_o;
	// Trace: design.sv:13357:5
	output wire [(N_REGS * 32) - 1:0] hwlp_counter_o;
	// Trace: design.sv:13361:3
	reg [(N_REGS * 32) - 1:0] hwlp_start_q;
	// Trace: design.sv:13362:3
	reg [(N_REGS * 32) - 1:0] hwlp_end_q;
	// Trace: design.sv:13363:3
	reg [(N_REGS * 32) - 1:0] hwlp_counter_q;
	wire [(N_REGS * 32) - 1:0] hwlp_counter_n;
	// Trace: design.sv:13365:3
	reg [31:0] i;
	// Trace: design.sv:13368:3
	assign hwlp_start_addr_o = hwlp_start_q;
	// Trace: design.sv:13369:3
	assign hwlp_end_addr_o = hwlp_end_q;
	// Trace: design.sv:13370:3
	assign hwlp_counter_o = hwlp_counter_q;
	// Trace: design.sv:13376:3
	always @(posedge clk or negedge rst_n) begin : HWLOOP_REGS_START
		// Trace: design.sv:13377:5
		if (rst_n == 1'b0)
			// Trace: design.sv:13378:7
			hwlp_start_q <= {N_REGS {32'b00000000000000000000000000000000}};
		else if (hwlp_we_i[0] == 1'b1)
			// Trace: design.sv:13380:7
			hwlp_start_q[hwlp_regid_i * 32+:32] <= hwlp_start_data_i;
	end
	// Trace: design.sv:13388:3
	always @(posedge clk or negedge rst_n) begin : HWLOOP_REGS_END
		// Trace: design.sv:13389:5
		if (rst_n == 1'b0)
			// Trace: design.sv:13390:7
			hwlp_end_q <= {N_REGS {32'b00000000000000000000000000000000}};
		else if (hwlp_we_i[1] == 1'b1)
			// Trace: design.sv:13392:7
			hwlp_end_q[hwlp_regid_i * 32+:32] <= hwlp_end_data_i;
	end
	// Trace: design.sv:13400:3
	genvar _gv_k_3;
	// Trace: design.sv:13401:3
	generate
		for (_gv_k_3 = 0; _gv_k_3 < N_REGS; _gv_k_3 = _gv_k_3 + 1) begin : genblk1
			localparam k = _gv_k_3;
			// Trace: design.sv:13402:5
			assign hwlp_counter_n[k * 32+:32] = hwlp_counter_q[k * 32+:32] - 1;
		end
	endgenerate
	// Trace: design.sv:13405:3
	always @(posedge clk or negedge rst_n) begin : HWLOOP_REGS_COUNTER
		// Trace: design.sv:13406:5
		if (rst_n == 1'b0)
			// Trace: design.sv:13407:7
			hwlp_counter_q <= {N_REGS {32'b00000000000000000000000000000000}};
		else
			// Trace: design.sv:13409:7
			for (i = 0; i < N_REGS; i = i + 1)
				begin
					// Trace: design.sv:13410:9
					if ((hwlp_we_i[2] == 1'b1) && (i == hwlp_regid_i))
						// Trace: design.sv:13411:11
						hwlp_counter_q[i * 32+:32] <= hwlp_cnt_data_i;
					else
						// Trace: design.sv:13413:11
						if (hwlp_dec_cnt_i[i] && valid_i)
							// Trace: design.sv:13413:45
							hwlp_counter_q[i * 32+:32] <= hwlp_counter_n[i * 32+:32];
				end
	end
endmodule
module cv32e40p_id_stage (
	clk,
	clk_ungated_i,
	rst_n,
	scan_cg_en_i,
	fetch_enable_i,
	ctrl_busy_o,
	is_decoding_o,
	instr_valid_i,
	instr_rdata_i,
	instr_req_o,
	is_compressed_i,
	illegal_c_insn_i,
	branch_in_ex_o,
	branch_decision_i,
	jump_target_o,
	clear_instr_valid_o,
	pc_set_o,
	pc_mux_o,
	exc_pc_mux_o,
	trap_addr_mux_o,
	is_fetch_failed_i,
	pc_id_i,
	halt_if_o,
	id_ready_o,
	ex_ready_i,
	wb_ready_i,
	id_valid_o,
	ex_valid_i,
	pc_ex_o,
	alu_operand_a_ex_o,
	alu_operand_b_ex_o,
	alu_operand_c_ex_o,
	bmask_a_ex_o,
	bmask_b_ex_o,
	imm_vec_ext_ex_o,
	alu_vec_mode_ex_o,
	regfile_waddr_ex_o,
	regfile_we_ex_o,
	regfile_alu_waddr_ex_o,
	regfile_alu_we_ex_o,
	alu_en_ex_o,
	alu_operator_ex_o,
	alu_is_clpx_ex_o,
	alu_is_subrot_ex_o,
	alu_clpx_shift_ex_o,
	mult_operator_ex_o,
	mult_operand_a_ex_o,
	mult_operand_b_ex_o,
	mult_operand_c_ex_o,
	mult_en_ex_o,
	mult_sel_subword_ex_o,
	mult_signed_mode_ex_o,
	mult_imm_ex_o,
	mult_dot_op_a_ex_o,
	mult_dot_op_b_ex_o,
	mult_dot_op_c_ex_o,
	mult_dot_signed_ex_o,
	mult_is_clpx_ex_o,
	mult_clpx_shift_ex_o,
	mult_clpx_img_ex_o,
	apu_en_ex_o,
	apu_op_ex_o,
	apu_lat_ex_o,
	apu_operands_ex_o,
	apu_flags_ex_o,
	apu_waddr_ex_o,
	apu_read_regs_o,
	apu_read_regs_valid_o,
	apu_read_dep_i,
	apu_write_regs_o,
	apu_write_regs_valid_o,
	apu_write_dep_i,
	apu_perf_dep_o,
	apu_busy_i,
	frm_i,
	csr_access_ex_o,
	csr_op_ex_o,
	current_priv_lvl_i,
	csr_irq_sec_o,
	csr_cause_o,
	csr_save_if_o,
	csr_save_id_o,
	csr_save_ex_o,
	csr_restore_mret_id_o,
	csr_restore_uret_id_o,
	csr_restore_dret_id_o,
	csr_save_cause_o,
	hwlp_start_o,
	hwlp_end_o,
	hwlp_cnt_o,
	hwlp_jump_o,
	hwlp_target_o,
	csr_hwlp_regid_i,
	csr_hwlp_we_i,
	csr_hwlp_data_i,
	data_req_ex_o,
	data_we_ex_o,
	data_type_ex_o,
	data_sign_ext_ex_o,
	data_reg_offset_ex_o,
	data_load_event_ex_o,
	data_misaligned_ex_o,
	prepost_useincr_ex_o,
	data_misaligned_i,
	data_err_i,
	data_err_ack_o,
	atop_ex_o,
	irq_i,
	irq_sec_i,
	mie_bypass_i,
	mip_o,
	m_irq_enable_i,
	u_irq_enable_i,
	irq_ack_o,
	irq_id_o,
	exc_cause_o,
	debug_mode_o,
	debug_cause_o,
	debug_csr_save_o,
	debug_req_i,
	debug_single_step_i,
	debug_ebreakm_i,
	debug_ebreaku_i,
	trigger_match_i,
	debug_p_elw_no_sleep_o,
	debug_havereset_o,
	debug_running_o,
	debug_halted_o,
	wake_from_sleep_o,
	regfile_waddr_wb_i,
	regfile_we_wb_i,
	regfile_wdata_wb_i,
	regfile_alu_waddr_fw_i,
	regfile_alu_we_fw_i,
	regfile_alu_wdata_fw_i,
	mult_multicycle_i,
	mhpmevent_minstret_o,
	mhpmevent_load_o,
	mhpmevent_store_o,
	mhpmevent_jump_o,
	mhpmevent_branch_o,
	mhpmevent_branch_taken_o,
	mhpmevent_compressed_o,
	mhpmevent_jr_stall_o,
	mhpmevent_imiss_o,
	mhpmevent_ld_stall_o,
	mhpmevent_pipe_stall_o,
	perf_imiss_i,
	mcounteren_i
);
	reg _sv2v_0;
	// removed import cv32e40p_pkg::*;
	// removed import cv32e40p_apu_core_pkg::*;
	// Trace: design.sv:13460:15
	parameter PULP_XPULP = 1;
	// Trace: design.sv:13461:15
	parameter PULP_CLUSTER = 0;
	// Trace: design.sv:13462:15
	parameter N_HWLP = 2;
	// Trace: design.sv:13463:15
	parameter N_HWLP_BITS = $clog2(N_HWLP);
	// Trace: design.sv:13464:15
	parameter PULP_SECURE = 0;
	// Trace: design.sv:13465:15
	parameter USE_PMP = 0;
	// Trace: design.sv:13466:15
	parameter A_EXTENSION = 0;
	// Trace: design.sv:13467:15
	parameter APU = 0;
	// Trace: design.sv:13468:15
	parameter FPU = 0;
	// Trace: design.sv:13469:15
	parameter PULP_ZFINX = 0;
	// Trace: design.sv:13470:15
	parameter APU_NARGS_CPU = 3;
	// Trace: design.sv:13471:15
	parameter APU_WOP_CPU = 6;
	// Trace: design.sv:13472:15
	parameter APU_NDSFLAGS_CPU = 15;
	// Trace: design.sv:13473:15
	parameter APU_NUSFLAGS_CPU = 5;
	// Trace: design.sv:13474:15
	parameter DEBUG_TRIGGER_EN = 1;
	// Trace: design.sv:13476:5
	input wire clk;
	// Trace: design.sv:13477:5
	input wire clk_ungated_i;
	// Trace: design.sv:13478:5
	input wire rst_n;
	// Trace: design.sv:13480:5
	input wire scan_cg_en_i;
	// Trace: design.sv:13482:5
	input wire fetch_enable_i;
	// Trace: design.sv:13483:5
	output wire ctrl_busy_o;
	// Trace: design.sv:13484:5
	output wire is_decoding_o;
	// Trace: design.sv:13487:5
	input wire instr_valid_i;
	// Trace: design.sv:13488:5
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:13489:5
	output wire instr_req_o;
	// Trace: design.sv:13490:5
	input wire is_compressed_i;
	// Trace: design.sv:13491:5
	input wire illegal_c_insn_i;
	// Trace: design.sv:13494:5
	output reg branch_in_ex_o;
	// Trace: design.sv:13495:5
	input wire branch_decision_i;
	// Trace: design.sv:13496:5
	output wire [31:0] jump_target_o;
	// Trace: design.sv:13499:5
	output wire clear_instr_valid_o;
	// Trace: design.sv:13500:5
	output wire pc_set_o;
	// Trace: design.sv:13501:5
	output wire [3:0] pc_mux_o;
	// Trace: design.sv:13502:5
	output wire [2:0] exc_pc_mux_o;
	// Trace: design.sv:13503:5
	output wire [1:0] trap_addr_mux_o;
	// Trace: design.sv:13506:5
	input wire is_fetch_failed_i;
	// Trace: design.sv:13508:5
	input wire [31:0] pc_id_i;
	// Trace: design.sv:13511:5
	output wire halt_if_o;
	// Trace: design.sv:13513:5
	output wire id_ready_o;
	// Trace: design.sv:13514:5
	input wire ex_ready_i;
	// Trace: design.sv:13515:5
	input wire wb_ready_i;
	// Trace: design.sv:13517:5
	output wire id_valid_o;
	// Trace: design.sv:13518:5
	input wire ex_valid_i;
	// Trace: design.sv:13521:5
	output reg [31:0] pc_ex_o;
	// Trace: design.sv:13523:5
	output reg [31:0] alu_operand_a_ex_o;
	// Trace: design.sv:13524:5
	output reg [31:0] alu_operand_b_ex_o;
	// Trace: design.sv:13525:5
	output reg [31:0] alu_operand_c_ex_o;
	// Trace: design.sv:13526:5
	output reg [4:0] bmask_a_ex_o;
	// Trace: design.sv:13527:5
	output reg [4:0] bmask_b_ex_o;
	// Trace: design.sv:13528:5
	output reg [1:0] imm_vec_ext_ex_o;
	// Trace: design.sv:13529:5
	output reg [1:0] alu_vec_mode_ex_o;
	// Trace: design.sv:13531:5
	output reg [5:0] regfile_waddr_ex_o;
	// Trace: design.sv:13532:5
	output reg regfile_we_ex_o;
	// Trace: design.sv:13534:5
	output reg [5:0] regfile_alu_waddr_ex_o;
	// Trace: design.sv:13535:5
	output reg regfile_alu_we_ex_o;
	// Trace: design.sv:13538:5
	output reg alu_en_ex_o;
	// Trace: design.sv:13539:5
	localparam cv32e40p_pkg_ALU_OP_WIDTH = 7;
	// removed localparam type cv32e40p_pkg_alu_opcode_e
	output reg [6:0] alu_operator_ex_o;
	// Trace: design.sv:13540:5
	output reg alu_is_clpx_ex_o;
	// Trace: design.sv:13541:5
	output reg alu_is_subrot_ex_o;
	// Trace: design.sv:13542:5
	output reg [1:0] alu_clpx_shift_ex_o;
	// Trace: design.sv:13545:5
	localparam cv32e40p_pkg_MUL_OP_WIDTH = 3;
	// removed localparam type cv32e40p_pkg_mul_opcode_e
	output reg [2:0] mult_operator_ex_o;
	// Trace: design.sv:13546:5
	output reg [31:0] mult_operand_a_ex_o;
	// Trace: design.sv:13547:5
	output reg [31:0] mult_operand_b_ex_o;
	// Trace: design.sv:13548:5
	output reg [31:0] mult_operand_c_ex_o;
	// Trace: design.sv:13549:5
	output reg mult_en_ex_o;
	// Trace: design.sv:13550:5
	output reg mult_sel_subword_ex_o;
	// Trace: design.sv:13551:5
	output reg [1:0] mult_signed_mode_ex_o;
	// Trace: design.sv:13552:5
	output reg [4:0] mult_imm_ex_o;
	// Trace: design.sv:13554:5
	output reg [31:0] mult_dot_op_a_ex_o;
	// Trace: design.sv:13555:5
	output reg [31:0] mult_dot_op_b_ex_o;
	// Trace: design.sv:13556:5
	output reg [31:0] mult_dot_op_c_ex_o;
	// Trace: design.sv:13557:5
	output reg [1:0] mult_dot_signed_ex_o;
	// Trace: design.sv:13558:5
	output reg mult_is_clpx_ex_o;
	// Trace: design.sv:13559:5
	output reg [1:0] mult_clpx_shift_ex_o;
	// Trace: design.sv:13560:5
	output reg mult_clpx_img_ex_o;
	// Trace: design.sv:13563:5
	output reg apu_en_ex_o;
	// Trace: design.sv:13564:5
	output reg [APU_WOP_CPU - 1:0] apu_op_ex_o;
	// Trace: design.sv:13565:5
	output reg [1:0] apu_lat_ex_o;
	// Trace: design.sv:13566:5
	output reg [(APU_NARGS_CPU * 32) - 1:0] apu_operands_ex_o;
	// Trace: design.sv:13567:5
	output reg [APU_NDSFLAGS_CPU - 1:0] apu_flags_ex_o;
	// Trace: design.sv:13568:5
	output reg [5:0] apu_waddr_ex_o;
	// Trace: design.sv:13570:5
	output wire [17:0] apu_read_regs_o;
	// Trace: design.sv:13571:5
	output wire [2:0] apu_read_regs_valid_o;
	// Trace: design.sv:13572:5
	input wire apu_read_dep_i;
	// Trace: design.sv:13573:5
	output wire [11:0] apu_write_regs_o;
	// Trace: design.sv:13574:5
	output wire [1:0] apu_write_regs_valid_o;
	// Trace: design.sv:13575:5
	input wire apu_write_dep_i;
	// Trace: design.sv:13576:5
	output wire apu_perf_dep_o;
	// Trace: design.sv:13577:5
	input wire apu_busy_i;
	// Trace: design.sv:13578:5
	localparam cv32e40p_pkg_C_RM = 3;
	input wire [2:0] frm_i;
	// Trace: design.sv:13581:5
	output reg csr_access_ex_o;
	// Trace: design.sv:13582:5
	localparam cv32e40p_pkg_CSR_OP_WIDTH = 2;
	// removed localparam type cv32e40p_pkg_csr_opcode_e
	output reg [1:0] csr_op_ex_o;
	// Trace: design.sv:13583:5
	// removed localparam type cv32e40p_pkg_PrivLvl_t
	input wire [1:0] current_priv_lvl_i;
	// Trace: design.sv:13584:5
	output wire csr_irq_sec_o;
	// Trace: design.sv:13585:5
	output wire [5:0] csr_cause_o;
	// Trace: design.sv:13586:5
	output wire csr_save_if_o;
	// Trace: design.sv:13587:5
	output wire csr_save_id_o;
	// Trace: design.sv:13588:5
	output wire csr_save_ex_o;
	// Trace: design.sv:13589:5
	output wire csr_restore_mret_id_o;
	// Trace: design.sv:13590:5
	output wire csr_restore_uret_id_o;
	// Trace: design.sv:13591:5
	output wire csr_restore_dret_id_o;
	// Trace: design.sv:13592:5
	output wire csr_save_cause_o;
	// Trace: design.sv:13595:5
	output wire [(N_HWLP * 32) - 1:0] hwlp_start_o;
	// Trace: design.sv:13596:5
	output wire [(N_HWLP * 32) - 1:0] hwlp_end_o;
	// Trace: design.sv:13597:5
	output wire [(N_HWLP * 32) - 1:0] hwlp_cnt_o;
	// Trace: design.sv:13598:5
	output wire hwlp_jump_o;
	// Trace: design.sv:13599:5
	output wire [31:0] hwlp_target_o;
	// Trace: design.sv:13602:5
	input wire [N_HWLP_BITS - 1:0] csr_hwlp_regid_i;
	// Trace: design.sv:13603:5
	input wire [2:0] csr_hwlp_we_i;
	// Trace: design.sv:13604:5
	input wire [31:0] csr_hwlp_data_i;
	// Trace: design.sv:13607:5
	output reg data_req_ex_o;
	// Trace: design.sv:13608:5
	output reg data_we_ex_o;
	// Trace: design.sv:13609:5
	output reg [1:0] data_type_ex_o;
	// Trace: design.sv:13610:5
	output reg [1:0] data_sign_ext_ex_o;
	// Trace: design.sv:13611:5
	output reg [1:0] data_reg_offset_ex_o;
	// Trace: design.sv:13612:5
	output reg data_load_event_ex_o;
	// Trace: design.sv:13614:5
	output reg data_misaligned_ex_o;
	// Trace: design.sv:13616:5
	output reg prepost_useincr_ex_o;
	// Trace: design.sv:13617:5
	input wire data_misaligned_i;
	// Trace: design.sv:13618:5
	input wire data_err_i;
	// Trace: design.sv:13619:5
	output wire data_err_ack_o;
	// Trace: design.sv:13621:5
	output reg [5:0] atop_ex_o;
	// Trace: design.sv:13624:5
	input wire [31:0] irq_i;
	// Trace: design.sv:13625:5
	input wire irq_sec_i;
	// Trace: design.sv:13626:5
	input wire [31:0] mie_bypass_i;
	// Trace: design.sv:13627:5
	output wire [31:0] mip_o;
	// Trace: design.sv:13628:5
	input wire m_irq_enable_i;
	// Trace: design.sv:13629:5
	input wire u_irq_enable_i;
	// Trace: design.sv:13630:5
	output wire irq_ack_o;
	// Trace: design.sv:13631:5
	output wire [4:0] irq_id_o;
	// Trace: design.sv:13632:5
	output wire [4:0] exc_cause_o;
	// Trace: design.sv:13635:5
	output wire debug_mode_o;
	// Trace: design.sv:13636:5
	output wire [2:0] debug_cause_o;
	// Trace: design.sv:13637:5
	output wire debug_csr_save_o;
	// Trace: design.sv:13638:5
	input wire debug_req_i;
	// Trace: design.sv:13639:5
	input wire debug_single_step_i;
	// Trace: design.sv:13640:5
	input wire debug_ebreakm_i;
	// Trace: design.sv:13641:5
	input wire debug_ebreaku_i;
	// Trace: design.sv:13642:5
	input wire trigger_match_i;
	// Trace: design.sv:13643:5
	output wire debug_p_elw_no_sleep_o;
	// Trace: design.sv:13644:5
	output wire debug_havereset_o;
	// Trace: design.sv:13645:5
	output wire debug_running_o;
	// Trace: design.sv:13646:5
	output wire debug_halted_o;
	// Trace: design.sv:13649:5
	output wire wake_from_sleep_o;
	// Trace: design.sv:13652:5
	input wire [5:0] regfile_waddr_wb_i;
	// Trace: design.sv:13653:5
	input wire regfile_we_wb_i;
	// Trace: design.sv:13654:5
	input wire [31:0] regfile_wdata_wb_i;
	// Trace: design.sv:13656:5
	input wire [5:0] regfile_alu_waddr_fw_i;
	// Trace: design.sv:13657:5
	input wire regfile_alu_we_fw_i;
	// Trace: design.sv:13658:5
	input wire [31:0] regfile_alu_wdata_fw_i;
	// Trace: design.sv:13661:5
	input wire mult_multicycle_i;
	// Trace: design.sv:13664:5
	output reg mhpmevent_minstret_o;
	// Trace: design.sv:13665:5
	output reg mhpmevent_load_o;
	// Trace: design.sv:13666:5
	output reg mhpmevent_store_o;
	// Trace: design.sv:13667:5
	output reg mhpmevent_jump_o;
	// Trace: design.sv:13668:5
	output reg mhpmevent_branch_o;
	// Trace: design.sv:13669:5
	output reg mhpmevent_branch_taken_o;
	// Trace: design.sv:13670:5
	output reg mhpmevent_compressed_o;
	// Trace: design.sv:13671:5
	output reg mhpmevent_jr_stall_o;
	// Trace: design.sv:13672:5
	output reg mhpmevent_imiss_o;
	// Trace: design.sv:13673:5
	output reg mhpmevent_ld_stall_o;
	// Trace: design.sv:13674:5
	output reg mhpmevent_pipe_stall_o;
	// Trace: design.sv:13676:5
	input wire perf_imiss_i;
	// Trace: design.sv:13677:5
	input wire [31:0] mcounteren_i;
	// Trace: design.sv:13681:3
	localparam REG_S1_MSB = 19;
	// Trace: design.sv:13682:3
	localparam REG_S1_LSB = 15;
	// Trace: design.sv:13684:3
	localparam REG_S2_MSB = 24;
	// Trace: design.sv:13685:3
	localparam REG_S2_LSB = 20;
	// Trace: design.sv:13687:3
	localparam REG_S4_MSB = 31;
	// Trace: design.sv:13688:3
	localparam REG_S4_LSB = 27;
	// Trace: design.sv:13690:3
	localparam REG_D_MSB = 11;
	// Trace: design.sv:13691:3
	localparam REG_D_LSB = 7;
	// Trace: design.sv:13693:3
	wire [31:0] instr;
	// Trace: design.sv:13697:3
	wire deassert_we;
	// Trace: design.sv:13699:3
	wire illegal_insn_dec;
	// Trace: design.sv:13700:3
	wire ebrk_insn_dec;
	// Trace: design.sv:13701:3
	wire mret_insn_dec;
	// Trace: design.sv:13702:3
	wire uret_insn_dec;
	// Trace: design.sv:13704:3
	wire dret_insn_dec;
	// Trace: design.sv:13706:3
	wire ecall_insn_dec;
	// Trace: design.sv:13707:3
	wire wfi_insn_dec;
	// Trace: design.sv:13709:3
	wire fencei_insn_dec;
	// Trace: design.sv:13711:3
	wire rega_used_dec;
	// Trace: design.sv:13712:3
	wire regb_used_dec;
	// Trace: design.sv:13713:3
	wire regc_used_dec;
	// Trace: design.sv:13715:3
	wire branch_taken_ex;
	// Trace: design.sv:13716:3
	wire [1:0] ctrl_transfer_insn_in_id;
	// Trace: design.sv:13717:3
	wire [1:0] ctrl_transfer_insn_in_dec;
	// Trace: design.sv:13719:3
	wire misaligned_stall;
	// Trace: design.sv:13720:3
	wire jr_stall;
	// Trace: design.sv:13721:3
	wire load_stall;
	// Trace: design.sv:13722:3
	wire csr_apu_stall;
	// Trace: design.sv:13723:3
	wire hwlp_mask;
	// Trace: design.sv:13724:3
	wire halt_id;
	// Trace: design.sv:13725:3
	wire halt_if;
	// Trace: design.sv:13727:3
	wire debug_wfi_no_sleep;
	// Trace: design.sv:13730:3
	wire [31:0] imm_i_type;
	// Trace: design.sv:13731:3
	wire [31:0] imm_iz_type;
	// Trace: design.sv:13732:3
	wire [31:0] imm_s_type;
	// Trace: design.sv:13733:3
	wire [31:0] imm_sb_type;
	// Trace: design.sv:13734:3
	wire [31:0] imm_u_type;
	// Trace: design.sv:13735:3
	wire [31:0] imm_uj_type;
	// Trace: design.sv:13736:3
	wire [31:0] imm_z_type;
	// Trace: design.sv:13737:3
	wire [31:0] imm_s2_type;
	// Trace: design.sv:13738:3
	wire [31:0] imm_bi_type;
	// Trace: design.sv:13739:3
	wire [31:0] imm_s3_type;
	// Trace: design.sv:13740:3
	wire [31:0] imm_vs_type;
	// Trace: design.sv:13741:3
	wire [31:0] imm_vu_type;
	// Trace: design.sv:13742:3
	wire [31:0] imm_shuffleb_type;
	// Trace: design.sv:13743:3
	wire [31:0] imm_shuffleh_type;
	// Trace: design.sv:13744:3
	reg [31:0] imm_shuffle_type;
	// Trace: design.sv:13745:3
	wire [31:0] imm_clip_type;
	// Trace: design.sv:13747:3
	reg [31:0] imm_a;
	// Trace: design.sv:13748:3
	reg [31:0] imm_b;
	// Trace: design.sv:13750:3
	reg [31:0] jump_target;
	// Trace: design.sv:13753:3
	wire irq_req_ctrl;
	// Trace: design.sv:13754:3
	wire irq_sec_ctrl;
	// Trace: design.sv:13755:3
	wire irq_wu_ctrl;
	// Trace: design.sv:13756:3
	wire [4:0] irq_id_ctrl;
	// Trace: design.sv:13759:3
	wire [5:0] regfile_addr_ra_id;
	// Trace: design.sv:13760:3
	wire [5:0] regfile_addr_rb_id;
	// Trace: design.sv:13761:3
	reg [5:0] regfile_addr_rc_id;
	// Trace: design.sv:13763:3
	wire regfile_fp_a;
	// Trace: design.sv:13764:3
	wire regfile_fp_b;
	// Trace: design.sv:13765:3
	wire regfile_fp_c;
	// Trace: design.sv:13766:3
	wire regfile_fp_d;
	// Trace: design.sv:13768:3
	wire [5:0] regfile_waddr_id;
	// Trace: design.sv:13769:3
	wire [5:0] regfile_alu_waddr_id;
	// Trace: design.sv:13770:3
	wire regfile_alu_we_id;
	wire regfile_alu_we_dec_id;
	// Trace: design.sv:13772:3
	wire [31:0] regfile_data_ra_id;
	// Trace: design.sv:13773:3
	wire [31:0] regfile_data_rb_id;
	// Trace: design.sv:13774:3
	wire [31:0] regfile_data_rc_id;
	// Trace: design.sv:13777:3
	wire alu_en;
	// Trace: design.sv:13778:3
	wire [6:0] alu_operator;
	// Trace: design.sv:13779:3
	wire [2:0] alu_op_a_mux_sel;
	// Trace: design.sv:13780:3
	wire [2:0] alu_op_b_mux_sel;
	// Trace: design.sv:13781:3
	wire [1:0] alu_op_c_mux_sel;
	// Trace: design.sv:13782:3
	wire [1:0] regc_mux;
	// Trace: design.sv:13784:3
	wire [0:0] imm_a_mux_sel;
	// Trace: design.sv:13785:3
	wire [3:0] imm_b_mux_sel;
	// Trace: design.sv:13786:3
	wire [1:0] ctrl_transfer_target_mux_sel;
	// Trace: design.sv:13789:3
	wire [2:0] mult_operator;
	// Trace: design.sv:13790:3
	wire mult_en;
	// Trace: design.sv:13791:3
	wire mult_int_en;
	// Trace: design.sv:13792:3
	wire mult_sel_subword;
	// Trace: design.sv:13793:3
	wire [1:0] mult_signed_mode;
	// Trace: design.sv:13794:3
	wire mult_dot_en;
	// Trace: design.sv:13795:3
	wire [1:0] mult_dot_signed;
	// Trace: design.sv:13798:3
	localparam [31:0] cv32e40p_fpu_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] cv32e40p_fpu_pkg_FP_FORMAT_BITS = 3;
	wire [2:0] fpu_src_fmt;
	// Trace: design.sv:13799:3
	wire [2:0] fpu_dst_fmt;
	// Trace: design.sv:13800:3
	localparam [31:0] cv32e40p_fpu_pkg_NUM_INT_FORMATS = 4;
	localparam [31:0] cv32e40p_fpu_pkg_INT_FORMAT_BITS = 2;
	wire [1:0] fpu_int_fmt;
	// Trace: design.sv:13803:3
	wire apu_en;
	// Trace: design.sv:13804:3
	wire [APU_WOP_CPU - 1:0] apu_op;
	// Trace: design.sv:13805:3
	wire [1:0] apu_lat;
	// Trace: design.sv:13806:3
	wire [(APU_NARGS_CPU * 32) - 1:0] apu_operands;
	// Trace: design.sv:13807:3
	wire [APU_NDSFLAGS_CPU - 1:0] apu_flags;
	// Trace: design.sv:13808:3
	wire [5:0] apu_waddr;
	// Trace: design.sv:13810:3
	reg [17:0] apu_read_regs;
	// Trace: design.sv:13811:3
	reg [2:0] apu_read_regs_valid;
	// Trace: design.sv:13812:3
	wire [11:0] apu_write_regs;
	// Trace: design.sv:13813:3
	wire [1:0] apu_write_regs_valid;
	// Trace: design.sv:13815:3
	wire apu_stall;
	// Trace: design.sv:13816:3
	wire [2:0] fp_rnd_mode;
	// Trace: design.sv:13819:3
	wire regfile_we_id;
	// Trace: design.sv:13820:3
	wire regfile_alu_waddr_mux_sel;
	// Trace: design.sv:13823:3
	wire data_we_id;
	// Trace: design.sv:13824:3
	wire [1:0] data_type_id;
	// Trace: design.sv:13825:3
	wire [1:0] data_sign_ext_id;
	// Trace: design.sv:13826:3
	wire [1:0] data_reg_offset_id;
	// Trace: design.sv:13827:3
	wire data_req_id;
	// Trace: design.sv:13828:3
	wire data_load_event_id;
	// Trace: design.sv:13831:3
	wire [5:0] atop_id;
	// Trace: design.sv:13834:3
	wire [N_HWLP_BITS - 1:0] hwlp_regid;
	wire [N_HWLP_BITS - 1:0] hwlp_regid_int;
	// Trace: design.sv:13835:3
	wire [2:0] hwlp_we;
	wire [2:0] hwlp_we_int;
	wire [2:0] hwlp_we_masked;
	// Trace: design.sv:13836:3
	wire hwlp_target_mux_sel;
	// Trace: design.sv:13837:3
	wire hwlp_start_mux_sel;
	// Trace: design.sv:13838:3
	wire hwlp_cnt_mux_sel;
	// Trace: design.sv:13840:3
	reg [31:0] hwlp_target;
	// Trace: design.sv:13841:3
	wire [31:0] hwlp_start;
	reg [31:0] hwlp_start_int;
	// Trace: design.sv:13842:3
	wire [31:0] hwlp_end;
	// Trace: design.sv:13843:3
	wire [31:0] hwlp_cnt;
	reg [31:0] hwlp_cnt_int;
	// Trace: design.sv:13844:3
	wire [N_HWLP - 1:0] hwlp_dec_cnt;
	// Trace: design.sv:13845:3
	wire hwlp_valid;
	// Trace: design.sv:13848:3
	wire csr_access;
	// Trace: design.sv:13849:3
	wire [1:0] csr_op;
	// Trace: design.sv:13850:3
	wire csr_status;
	// Trace: design.sv:13852:3
	wire prepost_useincr;
	// Trace: design.sv:13855:3
	wire [1:0] operand_a_fw_mux_sel;
	// Trace: design.sv:13856:3
	wire [1:0] operand_b_fw_mux_sel;
	// Trace: design.sv:13857:3
	wire [1:0] operand_c_fw_mux_sel;
	// Trace: design.sv:13858:3
	reg [31:0] operand_a_fw_id;
	// Trace: design.sv:13859:3
	reg [31:0] operand_b_fw_id;
	// Trace: design.sv:13860:3
	reg [31:0] operand_c_fw_id;
	// Trace: design.sv:13862:3
	reg [31:0] operand_b;
	reg [31:0] operand_b_vec;
	// Trace: design.sv:13863:3
	reg [31:0] operand_c;
	reg [31:0] operand_c_vec;
	// Trace: design.sv:13865:3
	reg [31:0] alu_operand_a;
	// Trace: design.sv:13866:3
	wire [31:0] alu_operand_b;
	// Trace: design.sv:13867:3
	wire [31:0] alu_operand_c;
	// Trace: design.sv:13870:3
	wire [0:0] bmask_a_mux;
	// Trace: design.sv:13871:3
	wire [1:0] bmask_b_mux;
	// Trace: design.sv:13872:3
	wire alu_bmask_a_mux_sel;
	// Trace: design.sv:13873:3
	wire alu_bmask_b_mux_sel;
	// Trace: design.sv:13874:3
	wire [0:0] mult_imm_mux;
	// Trace: design.sv:13876:3
	reg [4:0] bmask_a_id_imm;
	// Trace: design.sv:13877:3
	reg [4:0] bmask_b_id_imm;
	// Trace: design.sv:13878:3
	reg [4:0] bmask_a_id;
	// Trace: design.sv:13879:3
	reg [4:0] bmask_b_id;
	// Trace: design.sv:13880:3
	wire [1:0] imm_vec_ext_id;
	// Trace: design.sv:13881:3
	reg [4:0] mult_imm_id;
	// Trace: design.sv:13883:3
	wire [1:0] alu_vec_mode;
	// Trace: design.sv:13884:3
	wire scalar_replication;
	// Trace: design.sv:13885:3
	wire scalar_replication_c;
	// Trace: design.sv:13888:3
	wire reg_d_ex_is_reg_a_id;
	// Trace: design.sv:13889:3
	wire reg_d_ex_is_reg_b_id;
	// Trace: design.sv:13890:3
	wire reg_d_ex_is_reg_c_id;
	// Trace: design.sv:13891:3
	wire reg_d_wb_is_reg_a_id;
	// Trace: design.sv:13892:3
	wire reg_d_wb_is_reg_b_id;
	// Trace: design.sv:13893:3
	wire reg_d_wb_is_reg_c_id;
	// Trace: design.sv:13894:3
	wire reg_d_alu_is_reg_a_id;
	// Trace: design.sv:13895:3
	wire reg_d_alu_is_reg_b_id;
	// Trace: design.sv:13896:3
	wire reg_d_alu_is_reg_c_id;
	// Trace: design.sv:13898:3
	wire is_clpx;
	wire is_subrot;
	// Trace: design.sv:13900:3
	wire mret_dec;
	// Trace: design.sv:13901:3
	wire uret_dec;
	// Trace: design.sv:13902:3
	wire dret_dec;
	// Trace: design.sv:13905:3
	reg id_valid_q;
	// Trace: design.sv:13906:3
	wire minstret;
	// Trace: design.sv:13907:3
	wire perf_pipeline_stall;
	// Trace: design.sv:13909:3
	assign instr = instr_rdata_i;
	// Trace: design.sv:13913:3
	assign imm_i_type = {{20 {instr[31]}}, instr[31:20]};
	// Trace: design.sv:13914:3
	assign imm_iz_type = {20'b00000000000000000000, instr[31:20]};
	// Trace: design.sv:13915:3
	assign imm_s_type = {{20 {instr[31]}}, instr[31:25], instr[11:7]};
	// Trace: design.sv:13916:3
	assign imm_sb_type = {{19 {instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
	// Trace: design.sv:13917:3
	assign imm_u_type = {instr[31:12], 12'b000000000000};
	// Trace: design.sv:13918:3
	assign imm_uj_type = {{12 {instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};
	// Trace: design.sv:13921:3
	assign imm_z_type = {27'b000000000000000000000000000, instr[REG_S1_MSB:REG_S1_LSB]};
	// Trace: design.sv:13923:3
	assign imm_s2_type = {27'b000000000000000000000000000, instr[24:20]};
	// Trace: design.sv:13924:3
	assign imm_bi_type = {{27 {instr[24]}}, instr[24:20]};
	// Trace: design.sv:13925:3
	assign imm_s3_type = {27'b000000000000000000000000000, instr[29:25]};
	// Trace: design.sv:13926:3
	assign imm_vs_type = {{26 {instr[24]}}, instr[24:20], instr[25]};
	// Trace: design.sv:13927:3
	assign imm_vu_type = {26'b00000000000000000000000000, instr[24:20], instr[25]};
	// Trace: design.sv:13930:3
	assign imm_shuffleb_type = {6'b000000, instr[28:27], 6'b000000, instr[24:23], 6'b000000, instr[22:21], 6'b000000, instr[20], instr[25]};
	// Trace: design.sv:13933:3
	assign imm_shuffleh_type = {15'h0000, instr[20], 15'h0000, instr[25]};
	// Trace: design.sv:13938:3
	assign imm_clip_type = (32'h00000001 << instr[24:20]) - 1;
	// Trace: design.sv:13943:3
	assign regfile_addr_ra_id = {regfile_fp_a, instr[REG_S1_MSB:REG_S1_LSB]};
	// Trace: design.sv:13944:3
	assign regfile_addr_rb_id = {regfile_fp_b, instr[REG_S2_MSB:REG_S2_LSB]};
	// Trace: design.sv:13947:3
	localparam cv32e40p_pkg_REGC_RD = 2'b01;
	localparam cv32e40p_pkg_REGC_S1 = 2'b10;
	localparam cv32e40p_pkg_REGC_S4 = 2'b00;
	localparam cv32e40p_pkg_REGC_ZERO = 2'b11;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:13948:5
		(* full_case, parallel_case *)
		case (regc_mux)
			cv32e40p_pkg_REGC_ZERO:
				// Trace: design.sv:13949:18
				regfile_addr_rc_id = 1'sb0;
			cv32e40p_pkg_REGC_RD:
				// Trace: design.sv:13950:18
				regfile_addr_rc_id = {regfile_fp_c, instr[REG_D_MSB:REG_D_LSB]};
			cv32e40p_pkg_REGC_S1:
				// Trace: design.sv:13951:18
				regfile_addr_rc_id = {regfile_fp_c, instr[REG_S1_MSB:REG_S1_LSB]};
			cv32e40p_pkg_REGC_S4:
				// Trace: design.sv:13952:18
				regfile_addr_rc_id = {regfile_fp_c, instr[REG_S4_MSB:REG_S4_LSB]};
		endcase
	end
	// Trace: design.sv:13959:3
	assign regfile_waddr_id = {regfile_fp_d, instr[REG_D_MSB:REG_D_LSB]};
	// Trace: design.sv:13963:3
	assign regfile_alu_waddr_id = (regfile_alu_waddr_mux_sel ? regfile_waddr_id : regfile_addr_ra_id);
	// Trace: design.sv:13966:3
	assign reg_d_ex_is_reg_a_id = ((regfile_waddr_ex_o == regfile_addr_ra_id) && (rega_used_dec == 1'b1)) && (regfile_addr_ra_id != {6 {1'sb0}});
	// Trace: design.sv:13967:3
	assign reg_d_ex_is_reg_b_id = ((regfile_waddr_ex_o == regfile_addr_rb_id) && (regb_used_dec == 1'b1)) && (regfile_addr_rb_id != {6 {1'sb0}});
	// Trace: design.sv:13968:3
	assign reg_d_ex_is_reg_c_id = ((regfile_waddr_ex_o == regfile_addr_rc_id) && (regc_used_dec == 1'b1)) && (regfile_addr_rc_id != {6 {1'sb0}});
	// Trace: design.sv:13969:3
	assign reg_d_wb_is_reg_a_id = ((regfile_waddr_wb_i == regfile_addr_ra_id) && (rega_used_dec == 1'b1)) && (regfile_addr_ra_id != {6 {1'sb0}});
	// Trace: design.sv:13970:3
	assign reg_d_wb_is_reg_b_id = ((regfile_waddr_wb_i == regfile_addr_rb_id) && (regb_used_dec == 1'b1)) && (regfile_addr_rb_id != {6 {1'sb0}});
	// Trace: design.sv:13971:3
	assign reg_d_wb_is_reg_c_id = ((regfile_waddr_wb_i == regfile_addr_rc_id) && (regc_used_dec == 1'b1)) && (regfile_addr_rc_id != {6 {1'sb0}});
	// Trace: design.sv:13972:3
	assign reg_d_alu_is_reg_a_id = ((regfile_alu_waddr_fw_i == regfile_addr_ra_id) && (rega_used_dec == 1'b1)) && (regfile_addr_ra_id != {6 {1'sb0}});
	// Trace: design.sv:13973:3
	assign reg_d_alu_is_reg_b_id = ((regfile_alu_waddr_fw_i == regfile_addr_rb_id) && (regb_used_dec == 1'b1)) && (regfile_addr_rb_id != {6 {1'sb0}});
	// Trace: design.sv:13974:3
	assign reg_d_alu_is_reg_c_id = ((regfile_alu_waddr_fw_i == regfile_addr_rc_id) && (regc_used_dec == 1'b1)) && (regfile_addr_rc_id != {6 {1'sb0}});
	// Trace: design.sv:13979:3
	assign clear_instr_valid_o = (id_ready_o | halt_id) | branch_taken_ex;
	// Trace: design.sv:13981:3
	assign branch_taken_ex = branch_in_ex_o && branch_decision_i;
	// Trace: design.sv:13984:3
	assign mult_en = mult_int_en | mult_dot_en;
	// Trace: design.sv:13996:3
	localparam cv32e40p_pkg_JT_COND = 2'b11;
	localparam cv32e40p_pkg_JT_JAL = 2'b01;
	localparam cv32e40p_pkg_JT_JALR = 2'b10;
	always @(*) begin : jump_target_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:13997:5
		(* full_case, parallel_case *)
		case (ctrl_transfer_target_mux_sel)
			cv32e40p_pkg_JT_JAL:
				// Trace: design.sv:13998:16
				jump_target = pc_id_i + imm_uj_type;
			cv32e40p_pkg_JT_COND:
				// Trace: design.sv:13999:16
				jump_target = pc_id_i + imm_sb_type;
			cv32e40p_pkg_JT_JALR:
				// Trace: design.sv:14002:16
				jump_target = regfile_data_ra_id + imm_i_type;
			default:
				// Trace: design.sv:14003:16
				jump_target = regfile_data_ra_id + imm_i_type;
		endcase
	end
	// Trace: design.sv:14007:3
	assign jump_target_o = jump_target;
	// Trace: design.sv:14020:3
	localparam cv32e40p_pkg_OP_A_CURRPC = 3'b001;
	localparam cv32e40p_pkg_OP_A_IMM = 3'b010;
	localparam cv32e40p_pkg_OP_A_REGA_OR_FWD = 3'b000;
	localparam cv32e40p_pkg_OP_A_REGB_OR_FWD = 3'b011;
	localparam cv32e40p_pkg_OP_A_REGC_OR_FWD = 3'b100;
	always @(*) begin : alu_operand_a_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:14021:5
		case (alu_op_a_mux_sel)
			cv32e40p_pkg_OP_A_REGA_OR_FWD:
				// Trace: design.sv:14022:25
				alu_operand_a = operand_a_fw_id;
			cv32e40p_pkg_OP_A_REGB_OR_FWD:
				// Trace: design.sv:14023:25
				alu_operand_a = operand_b_fw_id;
			cv32e40p_pkg_OP_A_REGC_OR_FWD:
				// Trace: design.sv:14024:25
				alu_operand_a = operand_c_fw_id;
			cv32e40p_pkg_OP_A_CURRPC:
				// Trace: design.sv:14025:25
				alu_operand_a = pc_id_i;
			cv32e40p_pkg_OP_A_IMM:
				// Trace: design.sv:14026:25
				alu_operand_a = imm_a;
			default:
				// Trace: design.sv:14027:25
				alu_operand_a = operand_a_fw_id;
		endcase
	end
	// Trace: design.sv:14032:3
	localparam cv32e40p_pkg_IMMA_Z = 1'b0;
	localparam cv32e40p_pkg_IMMA_ZERO = 1'b1;
	always @(*) begin : immediate_a_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:14033:5
		(* full_case, parallel_case *)
		case (imm_a_mux_sel)
			cv32e40p_pkg_IMMA_Z:
				// Trace: design.sv:14034:18
				imm_a = imm_z_type;
			cv32e40p_pkg_IMMA_ZERO:
				// Trace: design.sv:14035:18
				imm_a = 1'sb0;
		endcase
	end
	// Trace: design.sv:14040:3
	localparam cv32e40p_pkg_SEL_FW_EX = 2'b01;
	localparam cv32e40p_pkg_SEL_FW_WB = 2'b10;
	localparam cv32e40p_pkg_SEL_REGFILE = 2'b00;
	always @(*) begin : operand_a_fw_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:14041:5
		case (operand_a_fw_mux_sel)
			cv32e40p_pkg_SEL_FW_EX:
				// Trace: design.sv:14042:20
				operand_a_fw_id = regfile_alu_wdata_fw_i;
			cv32e40p_pkg_SEL_FW_WB:
				// Trace: design.sv:14043:20
				operand_a_fw_id = regfile_wdata_wb_i;
			cv32e40p_pkg_SEL_REGFILE:
				// Trace: design.sv:14044:20
				operand_a_fw_id = regfile_data_ra_id;
			default:
				// Trace: design.sv:14045:20
				operand_a_fw_id = regfile_data_ra_id;
		endcase
	end
	// Trace: design.sv:14060:3
	localparam cv32e40p_pkg_IMMB_BI = 4'b1011;
	localparam cv32e40p_pkg_IMMB_CLIP = 4'b1001;
	localparam cv32e40p_pkg_IMMB_I = 4'b0000;
	localparam cv32e40p_pkg_IMMB_PCINCR = 4'b0011;
	localparam cv32e40p_pkg_IMMB_S = 4'b0001;
	localparam cv32e40p_pkg_IMMB_S2 = 4'b0100;
	localparam cv32e40p_pkg_IMMB_S3 = 4'b0101;
	localparam cv32e40p_pkg_IMMB_SHUF = 4'b1000;
	localparam cv32e40p_pkg_IMMB_U = 4'b0010;
	localparam cv32e40p_pkg_IMMB_VS = 4'b0110;
	localparam cv32e40p_pkg_IMMB_VU = 4'b0111;
	always @(*) begin : immediate_b_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:14061:5
		(* full_case, parallel_case *)
		case (imm_b_mux_sel)
			cv32e40p_pkg_IMMB_I:
				// Trace: design.sv:14062:20
				imm_b = imm_i_type;
			cv32e40p_pkg_IMMB_S:
				// Trace: design.sv:14063:20
				imm_b = imm_s_type;
			cv32e40p_pkg_IMMB_U:
				// Trace: design.sv:14064:20
				imm_b = imm_u_type;
			cv32e40p_pkg_IMMB_PCINCR:
				// Trace: design.sv:14065:20
				imm_b = (is_compressed_i ? 32'h00000002 : 32'h00000004);
			cv32e40p_pkg_IMMB_S2:
				// Trace: design.sv:14066:20
				imm_b = imm_s2_type;
			cv32e40p_pkg_IMMB_BI:
				// Trace: design.sv:14067:20
				imm_b = imm_bi_type;
			cv32e40p_pkg_IMMB_S3:
				// Trace: design.sv:14068:20
				imm_b = imm_s3_type;
			cv32e40p_pkg_IMMB_VS:
				// Trace: design.sv:14069:20
				imm_b = imm_vs_type;
			cv32e40p_pkg_IMMB_VU:
				// Trace: design.sv:14070:20
				imm_b = imm_vu_type;
			cv32e40p_pkg_IMMB_SHUF:
				// Trace: design.sv:14071:20
				imm_b = imm_shuffle_type;
			cv32e40p_pkg_IMMB_CLIP:
				// Trace: design.sv:14072:20
				imm_b = {1'b0, imm_clip_type[31:1]};
			default:
				// Trace: design.sv:14073:20
				imm_b = imm_i_type;
		endcase
	end
	// Trace: design.sv:14078:3
	localparam cv32e40p_pkg_OP_B_BMASK = 3'b100;
	localparam cv32e40p_pkg_OP_B_IMM = 3'b010;
	localparam cv32e40p_pkg_OP_B_REGA_OR_FWD = 3'b011;
	localparam cv32e40p_pkg_OP_B_REGB_OR_FWD = 3'b000;
	localparam cv32e40p_pkg_OP_B_REGC_OR_FWD = 3'b001;
	always @(*) begin : alu_operand_b_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:14079:5
		case (alu_op_b_mux_sel)
			cv32e40p_pkg_OP_B_REGA_OR_FWD:
				// Trace: design.sv:14080:25
				operand_b = operand_a_fw_id;
			cv32e40p_pkg_OP_B_REGB_OR_FWD:
				// Trace: design.sv:14081:25
				operand_b = operand_b_fw_id;
			cv32e40p_pkg_OP_B_REGC_OR_FWD:
				// Trace: design.sv:14082:25
				operand_b = operand_c_fw_id;
			cv32e40p_pkg_OP_B_IMM:
				// Trace: design.sv:14083:25
				operand_b = imm_b;
			cv32e40p_pkg_OP_B_BMASK:
				// Trace: design.sv:14084:25
				operand_b = $unsigned(operand_b_fw_id[4:0]);
			default:
				// Trace: design.sv:14085:25
				operand_b = operand_b_fw_id;
		endcase
	end
	// Trace: design.sv:14091:3
	localparam cv32e40p_pkg_VEC_MODE8 = 2'b11;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:14092:5
		if (alu_vec_mode == cv32e40p_pkg_VEC_MODE8) begin
			// Trace: design.sv:14093:7
			operand_b_vec = {4 {operand_b[7:0]}};
			// Trace: design.sv:14094:7
			imm_shuffle_type = imm_shuffleb_type;
		end
		else begin
			// Trace: design.sv:14096:7
			operand_b_vec = {2 {operand_b[15:0]}};
			// Trace: design.sv:14097:7
			imm_shuffle_type = imm_shuffleh_type;
		end
	end
	// Trace: design.sv:14102:3
	assign alu_operand_b = (scalar_replication == 1'b1 ? operand_b_vec : operand_b);
	// Trace: design.sv:14106:3
	always @(*) begin : operand_b_fw_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:14107:5
		case (operand_b_fw_mux_sel)
			cv32e40p_pkg_SEL_FW_EX:
				// Trace: design.sv:14108:20
				operand_b_fw_id = regfile_alu_wdata_fw_i;
			cv32e40p_pkg_SEL_FW_WB:
				// Trace: design.sv:14109:20
				operand_b_fw_id = regfile_wdata_wb_i;
			cv32e40p_pkg_SEL_REGFILE:
				// Trace: design.sv:14110:20
				operand_b_fw_id = regfile_data_rb_id;
			default:
				// Trace: design.sv:14111:20
				operand_b_fw_id = regfile_data_rb_id;
		endcase
	end
	// Trace: design.sv:14127:3
	localparam cv32e40p_pkg_OP_C_JT = 2'b10;
	localparam cv32e40p_pkg_OP_C_REGB_OR_FWD = 2'b01;
	localparam cv32e40p_pkg_OP_C_REGC_OR_FWD = 2'b00;
	always @(*) begin : alu_operand_c_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:14128:5
		case (alu_op_c_mux_sel)
			cv32e40p_pkg_OP_C_REGC_OR_FWD:
				// Trace: design.sv:14129:25
				operand_c = operand_c_fw_id;
			cv32e40p_pkg_OP_C_REGB_OR_FWD:
				// Trace: design.sv:14130:25
				operand_c = operand_b_fw_id;
			cv32e40p_pkg_OP_C_JT:
				// Trace: design.sv:14131:25
				operand_c = jump_target;
			default:
				// Trace: design.sv:14132:25
				operand_c = operand_c_fw_id;
		endcase
	end
	// Trace: design.sv:14138:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:14139:5
		if (alu_vec_mode == cv32e40p_pkg_VEC_MODE8)
			// Trace: design.sv:14140:7
			operand_c_vec = {4 {operand_c[7:0]}};
		else
			// Trace: design.sv:14142:7
			operand_c_vec = {2 {operand_c[15:0]}};
	end
	// Trace: design.sv:14147:3
	assign alu_operand_c = (scalar_replication_c == 1'b1 ? operand_c_vec : operand_c);
	// Trace: design.sv:14151:3
	always @(*) begin : operand_c_fw_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:14152:5
		case (operand_c_fw_mux_sel)
			cv32e40p_pkg_SEL_FW_EX:
				// Trace: design.sv:14153:20
				operand_c_fw_id = regfile_alu_wdata_fw_i;
			cv32e40p_pkg_SEL_FW_WB:
				// Trace: design.sv:14154:20
				operand_c_fw_id = regfile_wdata_wb_i;
			cv32e40p_pkg_SEL_REGFILE:
				// Trace: design.sv:14155:20
				operand_c_fw_id = regfile_data_rc_id;
			default:
				// Trace: design.sv:14156:20
				operand_c_fw_id = regfile_data_rc_id;
		endcase
	end
	// Trace: design.sv:14171:3
	localparam cv32e40p_pkg_BMASK_A_S3 = 1'b1;
	localparam cv32e40p_pkg_BMASK_A_ZERO = 1'b0;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:14172:5
		(* full_case, parallel_case *)
		case (bmask_a_mux)
			cv32e40p_pkg_BMASK_A_ZERO:
				// Trace: design.sv:14173:21
				bmask_a_id_imm = 1'sb0;
			cv32e40p_pkg_BMASK_A_S3:
				// Trace: design.sv:14174:21
				bmask_a_id_imm = imm_s3_type[4:0];
		endcase
	end
	// Trace: design.sv:14177:3
	localparam cv32e40p_pkg_BMASK_B_ONE = 2'b11;
	localparam cv32e40p_pkg_BMASK_B_S2 = 2'b00;
	localparam cv32e40p_pkg_BMASK_B_S3 = 2'b01;
	localparam cv32e40p_pkg_BMASK_B_ZERO = 2'b10;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:14178:5
		(* full_case, parallel_case *)
		case (bmask_b_mux)
			cv32e40p_pkg_BMASK_B_ZERO:
				// Trace: design.sv:14179:21
				bmask_b_id_imm = 1'sb0;
			cv32e40p_pkg_BMASK_B_ONE:
				// Trace: design.sv:14180:21
				bmask_b_id_imm = 5'd1;
			cv32e40p_pkg_BMASK_B_S2:
				// Trace: design.sv:14181:21
				bmask_b_id_imm = imm_s2_type[4:0];
			cv32e40p_pkg_BMASK_B_S3:
				// Trace: design.sv:14182:21
				bmask_b_id_imm = imm_s3_type[4:0];
		endcase
	end
	// Trace: design.sv:14186:3
	localparam cv32e40p_pkg_BMASK_A_IMM = 1'b1;
	localparam cv32e40p_pkg_BMASK_A_REG = 1'b0;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:14187:5
		(* full_case, parallel_case *)
		case (alu_bmask_a_mux_sel)
			cv32e40p_pkg_BMASK_A_IMM:
				// Trace: design.sv:14188:20
				bmask_a_id = bmask_a_id_imm;
			cv32e40p_pkg_BMASK_A_REG:
				// Trace: design.sv:14189:20
				bmask_a_id = operand_b_fw_id[9:5];
		endcase
	end
	// Trace: design.sv:14192:3
	localparam cv32e40p_pkg_BMASK_B_IMM = 1'b1;
	localparam cv32e40p_pkg_BMASK_B_REG = 1'b0;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:14193:5
		(* full_case, parallel_case *)
		case (alu_bmask_b_mux_sel)
			cv32e40p_pkg_BMASK_B_IMM:
				// Trace: design.sv:14194:20
				bmask_b_id = bmask_b_id_imm;
			cv32e40p_pkg_BMASK_B_REG:
				// Trace: design.sv:14195:20
				bmask_b_id = operand_b_fw_id[4:0];
		endcase
	end
	// Trace: design.sv:14199:3
	assign imm_vec_ext_id = imm_vu_type[1:0];
	// Trace: design.sv:14202:3
	localparam cv32e40p_pkg_MIMM_S3 = 1'b1;
	localparam cv32e40p_pkg_MIMM_ZERO = 1'b0;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:14203:5
		(* full_case, parallel_case *)
		case (mult_imm_mux)
			cv32e40p_pkg_MIMM_ZERO:
				// Trace: design.sv:14204:18
				mult_imm_id = 1'sb0;
			cv32e40p_pkg_MIMM_S3:
				// Trace: design.sv:14205:18
				mult_imm_id = imm_s3_type[4:0];
		endcase
	end
	// Trace: design.sv:14213:3
	generate
		if (APU == 1) begin : gen_apu
			if (APU_NARGS_CPU >= 1) begin : genblk1
				// Trace: design.sv:14216:31
				assign apu_operands[0+:32] = alu_operand_a;
			end
			if (APU_NARGS_CPU >= 2) begin : genblk2
				// Trace: design.sv:14217:31
				assign apu_operands[32+:32] = alu_operand_b;
			end
			if (APU_NARGS_CPU >= 3) begin : genblk3
				// Trace: design.sv:14218:31
				assign apu_operands[64+:32] = alu_operand_c;
			end
			// Trace: design.sv:14221:7
			assign apu_waddr = regfile_alu_waddr_id;
			// Trace: design.sv:14224:7
			assign apu_flags = (FPU == 1 ? {fpu_int_fmt, fpu_src_fmt, fpu_dst_fmt, fp_rnd_mode} : {APU_NDSFLAGS_CPU {1'sb0}});
			// Trace: design.sv:14227:7
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:14228:9
				(* full_case, parallel_case *)
				case (alu_op_a_mux_sel)
					cv32e40p_pkg_OP_A_REGA_OR_FWD: begin
						// Trace: design.sv:14230:13
						apu_read_regs[0+:6] = regfile_addr_ra_id;
						// Trace: design.sv:14231:13
						apu_read_regs_valid[0] = 1'b1;
					end
					cv32e40p_pkg_OP_A_REGB_OR_FWD: begin
						// Trace: design.sv:14234:13
						apu_read_regs[0+:6] = regfile_addr_rb_id;
						// Trace: design.sv:14235:13
						apu_read_regs_valid[0] = 1'b1;
					end
					default: begin
						// Trace: design.sv:14238:13
						apu_read_regs[0+:6] = regfile_addr_ra_id;
						// Trace: design.sv:14239:13
						apu_read_regs_valid[0] = 1'b0;
					end
				endcase
			end
			// Trace: design.sv:14244:7
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:14245:9
				(* full_case, parallel_case *)
				case (alu_op_b_mux_sel)
					cv32e40p_pkg_OP_B_REGA_OR_FWD: begin
						// Trace: design.sv:14247:13
						apu_read_regs[6+:6] = regfile_addr_ra_id;
						// Trace: design.sv:14248:13
						apu_read_regs_valid[1] = 1'b1;
					end
					cv32e40p_pkg_OP_B_REGB_OR_FWD: begin
						// Trace: design.sv:14251:13
						apu_read_regs[6+:6] = regfile_addr_rb_id;
						// Trace: design.sv:14252:13
						apu_read_regs_valid[1] = 1'b1;
					end
					cv32e40p_pkg_OP_B_REGC_OR_FWD: begin
						// Trace: design.sv:14255:13
						apu_read_regs[6+:6] = regfile_addr_rc_id;
						// Trace: design.sv:14256:13
						apu_read_regs_valid[1] = 1'b1;
					end
					default: begin
						// Trace: design.sv:14259:13
						apu_read_regs[6+:6] = regfile_addr_rb_id;
						// Trace: design.sv:14260:13
						apu_read_regs_valid[1] = 1'b0;
					end
				endcase
			end
			// Trace: design.sv:14265:7
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:14266:9
				(* full_case, parallel_case *)
				case (alu_op_c_mux_sel)
					cv32e40p_pkg_OP_C_REGB_OR_FWD: begin
						// Trace: design.sv:14268:13
						apu_read_regs[12+:6] = regfile_addr_rb_id;
						// Trace: design.sv:14269:13
						apu_read_regs_valid[2] = 1'b1;
					end
					cv32e40p_pkg_OP_C_REGC_OR_FWD: begin
						// Trace: design.sv:14272:13
						apu_read_regs[12+:6] = regfile_addr_rc_id;
						// Trace: design.sv:14273:13
						apu_read_regs_valid[2] = 1'b1;
					end
					default: begin
						// Trace: design.sv:14276:13
						apu_read_regs[12+:6] = regfile_addr_rc_id;
						// Trace: design.sv:14277:13
						apu_read_regs_valid[2] = 1'b0;
					end
				endcase
			end
			// Trace: design.sv:14282:7
			assign apu_write_regs[0+:6] = regfile_alu_waddr_id;
			// Trace: design.sv:14283:7
			assign apu_write_regs_valid[0] = regfile_alu_we_id;
			// Trace: design.sv:14285:7
			assign apu_write_regs[6+:6] = regfile_waddr_id;
			// Trace: design.sv:14286:7
			assign apu_write_regs_valid[1] = regfile_we_id;
			// Trace: design.sv:14288:7
			assign apu_read_regs_o = apu_read_regs;
			// Trace: design.sv:14289:7
			assign apu_read_regs_valid_o = apu_read_regs_valid;
			// Trace: design.sv:14291:7
			assign apu_write_regs_o = apu_write_regs;
			// Trace: design.sv:14292:7
			assign apu_write_regs_valid_o = apu_write_regs_valid;
		end
		else begin : gen_no_apu
			genvar _gv_i_2;
			for (_gv_i_2 = 0; _gv_i_2 < APU_NARGS_CPU; _gv_i_2 = _gv_i_2 + 1) begin : gen_apu_tie_off
				localparam i = _gv_i_2;
				// Trace: design.sv:14295:9
				assign apu_operands[i * 32+:32] = 1'sb0;
			end
			// Trace: design.sv:14298:7
			wire [18:1] sv2v_tmp_B43AF;
			assign sv2v_tmp_B43AF = 1'sb0;
			always @(*) apu_read_regs = sv2v_tmp_B43AF;
			// Trace: design.sv:14299:7
			wire [3:1] sv2v_tmp_093B8;
			assign sv2v_tmp_093B8 = 1'sb0;
			always @(*) apu_read_regs_valid = sv2v_tmp_093B8;
			// Trace: design.sv:14300:7
			assign apu_write_regs = 1'sb0;
			// Trace: design.sv:14301:7
			assign apu_write_regs_valid = 1'sb0;
			// Trace: design.sv:14302:7
			assign apu_waddr = 1'sb0;
			// Trace: design.sv:14303:7
			assign apu_flags = 1'sb0;
			// Trace: design.sv:14304:7
			assign apu_write_regs_o = 1'sb0;
			// Trace: design.sv:14305:7
			assign apu_read_regs_o = 1'sb0;
			// Trace: design.sv:14306:7
			assign apu_write_regs_valid_o = 1'sb0;
			// Trace: design.sv:14307:7
			assign apu_read_regs_valid_o = 1'sb0;
		end
	endgenerate
	// Trace: design.sv:14311:3
	assign apu_perf_dep_o = apu_stall;
	// Trace: design.sv:14313:3
	assign csr_apu_stall = csr_access & ((apu_en_ex_o & (apu_lat_ex_o[1] == 1'b1)) | apu_busy_i);
	// Trace: design.sv:14324:3
	cv32e40p_register_file #(
		.ADDR_WIDTH(6),
		.DATA_WIDTH(32),
		.FPU(FPU),
		.PULP_ZFINX(PULP_ZFINX)
	) register_file_i(
		.clk(clk),
		.rst_n(rst_n),
		.scan_cg_en_i(scan_cg_en_i),
		.raddr_a_i(regfile_addr_ra_id),
		.rdata_a_o(regfile_data_ra_id),
		.raddr_b_i(regfile_addr_rb_id),
		.rdata_b_o(regfile_data_rb_id),
		.raddr_c_i(regfile_addr_rc_id),
		.rdata_c_o(regfile_data_rc_id),
		.waddr_a_i(regfile_waddr_wb_i),
		.wdata_a_i(regfile_wdata_wb_i),
		.we_a_i(regfile_we_wb_i),
		.waddr_b_i(regfile_alu_waddr_fw_i),
		.wdata_b_i(regfile_alu_wdata_fw_i),
		.we_b_i(regfile_alu_we_fw_i)
	);
	// Trace: design.sv:14368:3
	cv32e40p_decoder #(
		.PULP_XPULP(PULP_XPULP),
		.PULP_CLUSTER(PULP_CLUSTER),
		.A_EXTENSION(A_EXTENSION),
		.FPU(FPU),
		.PULP_ZFINX(PULP_ZFINX),
		.PULP_SECURE(PULP_SECURE),
		.USE_PMP(USE_PMP),
		.APU_WOP_CPU(APU_WOP_CPU),
		.DEBUG_TRIGGER_EN(DEBUG_TRIGGER_EN)
	) decoder_i(
		.deassert_we_i(deassert_we),
		.illegal_insn_o(illegal_insn_dec),
		.ebrk_insn_o(ebrk_insn_dec),
		.mret_insn_o(mret_insn_dec),
		.uret_insn_o(uret_insn_dec),
		.dret_insn_o(dret_insn_dec),
		.mret_dec_o(mret_dec),
		.uret_dec_o(uret_dec),
		.dret_dec_o(dret_dec),
		.ecall_insn_o(ecall_insn_dec),
		.wfi_o(wfi_insn_dec),
		.fencei_insn_o(fencei_insn_dec),
		.rega_used_o(rega_used_dec),
		.regb_used_o(regb_used_dec),
		.regc_used_o(regc_used_dec),
		.reg_fp_a_o(regfile_fp_a),
		.reg_fp_b_o(regfile_fp_b),
		.reg_fp_c_o(regfile_fp_c),
		.reg_fp_d_o(regfile_fp_d),
		.bmask_a_mux_o(bmask_a_mux),
		.bmask_b_mux_o(bmask_b_mux),
		.alu_bmask_a_mux_sel_o(alu_bmask_a_mux_sel),
		.alu_bmask_b_mux_sel_o(alu_bmask_b_mux_sel),
		.instr_rdata_i(instr),
		.illegal_c_insn_i(illegal_c_insn_i),
		.alu_en_o(alu_en),
		.alu_operator_o(alu_operator),
		.alu_op_a_mux_sel_o(alu_op_a_mux_sel),
		.alu_op_b_mux_sel_o(alu_op_b_mux_sel),
		.alu_op_c_mux_sel_o(alu_op_c_mux_sel),
		.alu_vec_mode_o(alu_vec_mode),
		.scalar_replication_o(scalar_replication),
		.scalar_replication_c_o(scalar_replication_c),
		.imm_a_mux_sel_o(imm_a_mux_sel),
		.imm_b_mux_sel_o(imm_b_mux_sel),
		.regc_mux_o(regc_mux),
		.is_clpx_o(is_clpx),
		.is_subrot_o(is_subrot),
		.mult_operator_o(mult_operator),
		.mult_int_en_o(mult_int_en),
		.mult_sel_subword_o(mult_sel_subword),
		.mult_signed_mode_o(mult_signed_mode),
		.mult_imm_mux_o(mult_imm_mux),
		.mult_dot_en_o(mult_dot_en),
		.mult_dot_signed_o(mult_dot_signed),
		.frm_i(frm_i),
		.fpu_src_fmt_o(fpu_src_fmt),
		.fpu_dst_fmt_o(fpu_dst_fmt),
		.fpu_int_fmt_o(fpu_int_fmt),
		.apu_en_o(apu_en),
		.apu_op_o(apu_op),
		.apu_lat_o(apu_lat),
		.fp_rnd_mode_o(fp_rnd_mode),
		.regfile_mem_we_o(regfile_we_id),
		.regfile_alu_we_o(regfile_alu_we_id),
		.regfile_alu_we_dec_o(regfile_alu_we_dec_id),
		.regfile_alu_waddr_sel_o(regfile_alu_waddr_mux_sel),
		.csr_access_o(csr_access),
		.csr_status_o(csr_status),
		.csr_op_o(csr_op),
		.current_priv_lvl_i(current_priv_lvl_i),
		.data_req_o(data_req_id),
		.data_we_o(data_we_id),
		.prepost_useincr_o(prepost_useincr),
		.data_type_o(data_type_id),
		.data_sign_extension_o(data_sign_ext_id),
		.data_reg_offset_o(data_reg_offset_id),
		.data_load_event_o(data_load_event_id),
		.atop_o(atop_id),
		.hwlp_we_o(hwlp_we_int),
		.hwlp_target_mux_sel_o(hwlp_target_mux_sel),
		.hwlp_start_mux_sel_o(hwlp_start_mux_sel),
		.hwlp_cnt_mux_sel_o(hwlp_cnt_mux_sel),
		.debug_mode_i(debug_mode_o),
		.debug_wfi_no_sleep_i(debug_wfi_no_sleep),
		.ctrl_transfer_insn_in_dec_o(ctrl_transfer_insn_in_dec),
		.ctrl_transfer_insn_in_id_o(ctrl_transfer_insn_in_id),
		.ctrl_transfer_target_mux_sel_o(ctrl_transfer_target_mux_sel),
		.mcounteren_i(mcounteren_i)
	);
	// Trace: design.sv:14503:3
	cv32e40p_controller #(
		.PULP_CLUSTER(PULP_CLUSTER),
		.PULP_XPULP(PULP_XPULP)
	) controller_i(
		.clk(clk),
		.clk_ungated_i(clk_ungated_i),
		.rst_n(rst_n),
		.fetch_enable_i(fetch_enable_i),
		.ctrl_busy_o(ctrl_busy_o),
		.is_decoding_o(is_decoding_o),
		.is_fetch_failed_i(is_fetch_failed_i),
		.deassert_we_o(deassert_we),
		.illegal_insn_i(illegal_insn_dec),
		.ecall_insn_i(ecall_insn_dec),
		.mret_insn_i(mret_insn_dec),
		.uret_insn_i(uret_insn_dec),
		.dret_insn_i(dret_insn_dec),
		.mret_dec_i(mret_dec),
		.uret_dec_i(uret_dec),
		.dret_dec_i(dret_dec),
		.wfi_i(wfi_insn_dec),
		.ebrk_insn_i(ebrk_insn_dec),
		.fencei_insn_i(fencei_insn_dec),
		.csr_status_i(csr_status),
		.hwlp_mask_o(hwlp_mask),
		.instr_valid_i(instr_valid_i),
		.instr_req_o(instr_req_o),
		.pc_set_o(pc_set_o),
		.pc_mux_o(pc_mux_o),
		.exc_pc_mux_o(exc_pc_mux_o),
		.exc_cause_o(exc_cause_o),
		.trap_addr_mux_o(trap_addr_mux_o),
		.pc_id_i(pc_id_i),
		.is_compressed_i(is_compressed_i),
		.hwlp_start_addr_i(hwlp_start_o),
		.hwlp_end_addr_i(hwlp_end_o),
		.hwlp_counter_i(hwlp_cnt_o),
		.hwlp_dec_cnt_o(hwlp_dec_cnt),
		.hwlp_jump_o(hwlp_jump_o),
		.hwlp_targ_addr_o(hwlp_target_o),
		.data_req_ex_i(data_req_ex_o),
		.data_we_ex_i(data_we_ex_o),
		.data_misaligned_i(data_misaligned_i),
		.data_load_event_i(data_load_event_id),
		.data_err_i(data_err_i),
		.data_err_ack_o(data_err_ack_o),
		.mult_multicycle_i(mult_multicycle_i),
		.apu_en_i(apu_en),
		.apu_read_dep_i(apu_read_dep_i),
		.apu_write_dep_i(apu_write_dep_i),
		.apu_stall_o(apu_stall),
		.branch_taken_ex_i(branch_taken_ex),
		.ctrl_transfer_insn_in_id_i(ctrl_transfer_insn_in_id),
		.ctrl_transfer_insn_in_dec_i(ctrl_transfer_insn_in_dec),
		.irq_wu_ctrl_i(irq_wu_ctrl),
		.irq_req_ctrl_i(irq_req_ctrl),
		.irq_sec_ctrl_i(irq_sec_ctrl),
		.irq_id_ctrl_i(irq_id_ctrl),
		.current_priv_lvl_i(current_priv_lvl_i),
		.irq_ack_o(irq_ack_o),
		.irq_id_o(irq_id_o),
		.debug_mode_o(debug_mode_o),
		.debug_cause_o(debug_cause_o),
		.debug_csr_save_o(debug_csr_save_o),
		.debug_req_i(debug_req_i),
		.debug_single_step_i(debug_single_step_i),
		.debug_ebreakm_i(debug_ebreakm_i),
		.debug_ebreaku_i(debug_ebreaku_i),
		.trigger_match_i(trigger_match_i),
		.debug_p_elw_no_sleep_o(debug_p_elw_no_sleep_o),
		.debug_wfi_no_sleep_o(debug_wfi_no_sleep),
		.debug_havereset_o(debug_havereset_o),
		.debug_running_o(debug_running_o),
		.debug_halted_o(debug_halted_o),
		.wake_from_sleep_o(wake_from_sleep_o),
		.csr_save_cause_o(csr_save_cause_o),
		.csr_cause_o(csr_cause_o),
		.csr_save_if_o(csr_save_if_o),
		.csr_save_id_o(csr_save_id_o),
		.csr_save_ex_o(csr_save_ex_o),
		.csr_restore_mret_id_o(csr_restore_mret_id_o),
		.csr_restore_uret_id_o(csr_restore_uret_id_o),
		.csr_restore_dret_id_o(csr_restore_dret_id_o),
		.csr_irq_sec_o(csr_irq_sec_o),
		.regfile_we_id_i(regfile_alu_we_dec_id),
		.regfile_alu_waddr_id_i(regfile_alu_waddr_id),
		.regfile_we_ex_i(regfile_we_ex_o),
		.regfile_waddr_ex_i(regfile_waddr_ex_o),
		.regfile_we_wb_i(regfile_we_wb_i),
		.regfile_alu_we_fw_i(regfile_alu_we_fw_i),
		.reg_d_ex_is_reg_a_i(reg_d_ex_is_reg_a_id),
		.reg_d_ex_is_reg_b_i(reg_d_ex_is_reg_b_id),
		.reg_d_ex_is_reg_c_i(reg_d_ex_is_reg_c_id),
		.reg_d_wb_is_reg_a_i(reg_d_wb_is_reg_a_id),
		.reg_d_wb_is_reg_b_i(reg_d_wb_is_reg_b_id),
		.reg_d_wb_is_reg_c_i(reg_d_wb_is_reg_c_id),
		.reg_d_alu_is_reg_a_i(reg_d_alu_is_reg_a_id),
		.reg_d_alu_is_reg_b_i(reg_d_alu_is_reg_b_id),
		.reg_d_alu_is_reg_c_i(reg_d_alu_is_reg_c_id),
		.operand_a_fw_mux_sel_o(operand_a_fw_mux_sel),
		.operand_b_fw_mux_sel_o(operand_b_fw_mux_sel),
		.operand_c_fw_mux_sel_o(operand_c_fw_mux_sel),
		.halt_if_o(halt_if),
		.halt_id_o(halt_id),
		.misaligned_stall_o(misaligned_stall),
		.jr_stall_o(jr_stall),
		.load_stall_o(load_stall),
		.id_ready_i(id_ready_o),
		.id_valid_i(id_valid_o),
		.ex_valid_i(ex_valid_i),
		.wb_ready_i(wb_ready_i),
		.perf_pipeline_stall_o(perf_pipeline_stall)
	);
	// Trace: design.sv:14684:3
	cv32e40p_int_controller #(.PULP_SECURE(PULP_SECURE)) int_controller_i(
		.clk(clk),
		.rst_n(rst_n),
		.irq_i(irq_i),
		.irq_sec_i(irq_sec_i),
		.irq_req_ctrl_o(irq_req_ctrl),
		.irq_sec_ctrl_o(irq_sec_ctrl),
		.irq_id_ctrl_o(irq_id_ctrl),
		.irq_wu_ctrl_o(irq_wu_ctrl),
		.mie_bypass_i(mie_bypass_i),
		.mip_o(mip_o),
		.m_ie_i(m_irq_enable_i),
		.u_ie_i(u_irq_enable_i),
		.current_priv_lvl_i(current_priv_lvl_i)
	);
	// Trace: design.sv:14708:3
	generate
		if (PULP_XPULP) begin : gen_hwloop_regs
			// Trace: design.sv:14721:7
			cv32e40p_hwloop_regs #(.N_REGS(N_HWLP)) hwloop_regs_i(
				.clk(clk),
				.rst_n(rst_n),
				.hwlp_start_data_i(hwlp_start),
				.hwlp_end_data_i(hwlp_end),
				.hwlp_cnt_data_i(hwlp_cnt),
				.hwlp_we_i(hwlp_we),
				.hwlp_regid_i(hwlp_regid),
				.valid_i(hwlp_valid),
				.hwlp_start_addr_o(hwlp_start_o),
				.hwlp_end_addr_o(hwlp_end_o),
				.hwlp_counter_o(hwlp_cnt_o),
				.hwlp_dec_cnt_i(hwlp_dec_cnt)
			);
			// Trace: design.sv:14746:7
			assign hwlp_valid = instr_valid_i & clear_instr_valid_o;
			// Trace: design.sv:14749:7
			assign hwlp_regid_int = instr[7];
			// Trace: design.sv:14752:7
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:14753:9
				case (hwlp_target_mux_sel)
					1'b0:
						// Trace: design.sv:14754:17
						hwlp_target = pc_id_i + {imm_iz_type[30:0], 1'b0};
					1'b1:
						// Trace: design.sv:14755:17
						hwlp_target = pc_id_i + {imm_z_type[30:0], 1'b0};
				endcase
			end
			// Trace: design.sv:14760:7
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:14761:9
				case (hwlp_start_mux_sel)
					1'b0:
						// Trace: design.sv:14762:17
						hwlp_start_int = hwlp_target;
					1'b1:
						// Trace: design.sv:14763:17
						hwlp_start_int = pc_id_i + 4;
				endcase
			end
			// Trace: design.sv:14769:7
			always @(*) begin : hwlp_cnt_mux
				if (_sv2v_0)
					;
				// Trace: design.sv:14770:9
				case (hwlp_cnt_mux_sel)
					1'b0:
						// Trace: design.sv:14771:17
						hwlp_cnt_int = imm_iz_type;
					1'b1:
						// Trace: design.sv:14772:17
						hwlp_cnt_int = operand_a_fw_id;
				endcase
			end
			// Trace: design.sv:14784:7
			assign hwlp_we_masked = (hwlp_we_int & ~{3 {hwlp_mask}}) & {3 {id_ready_o}};
			// Trace: design.sv:14787:7
			assign hwlp_start = (hwlp_we_masked[0] ? hwlp_start_int : csr_hwlp_data_i);
			// Trace: design.sv:14788:7
			assign hwlp_end = (hwlp_we_masked[1] ? hwlp_target : csr_hwlp_data_i);
			// Trace: design.sv:14789:7
			assign hwlp_cnt = (hwlp_we_masked[2] ? hwlp_cnt_int : csr_hwlp_data_i);
			// Trace: design.sv:14790:7
			assign hwlp_regid = (|hwlp_we_masked ? hwlp_regid_int : csr_hwlp_regid_i);
			// Trace: design.sv:14791:7
			assign hwlp_we = (|hwlp_we_masked ? hwlp_we_masked : csr_hwlp_we_i);
		end
		else begin : gen_no_hwloop_regs
			// Trace: design.sv:14795:7
			assign hwlp_start_o = 'b0;
			// Trace: design.sv:14796:7
			assign hwlp_end_o = 'b0;
			// Trace: design.sv:14797:7
			assign hwlp_cnt_o = 'b0;
			// Trace: design.sv:14798:7
			assign hwlp_valid = 'b0;
			// Trace: design.sv:14799:7
			assign hwlp_regid_int = 'b0;
			// Trace: design.sv:14800:7
			wire [32:1] sv2v_tmp_18A71;
			assign sv2v_tmp_18A71 = 'b0;
			always @(*) hwlp_target = sv2v_tmp_18A71;
			// Trace: design.sv:14801:7
			wire [32:1] sv2v_tmp_B96B9;
			assign sv2v_tmp_B96B9 = 'b0;
			always @(*) hwlp_start_int = sv2v_tmp_B96B9;
			// Trace: design.sv:14802:7
			wire [32:1] sv2v_tmp_658E6;
			assign sv2v_tmp_658E6 = 'b0;
			always @(*) hwlp_cnt_int = sv2v_tmp_658E6;
			// Trace: design.sv:14803:7
			assign hwlp_we_masked = 'b0;
			// Trace: design.sv:14804:7
			assign hwlp_start = 'b0;
			// Trace: design.sv:14805:7
			assign hwlp_end = 'b0;
			// Trace: design.sv:14806:7
			assign hwlp_cnt = 'b0;
			// Trace: design.sv:14807:7
			assign hwlp_regid = 'b0;
			// Trace: design.sv:14808:7
			assign hwlp_we = 'b0;
		end
	endgenerate
	// Trace: design.sv:14823:3
	localparam cv32e40p_pkg_BRANCH_COND = 2'b11;
	function automatic [6:0] sv2v_cast_C07C4;
		input reg [6:0] inp;
		sv2v_cast_C07C4 = inp;
	endfunction
	function automatic [2:0] sv2v_cast_9F558;
		input reg [2:0] inp;
		sv2v_cast_9F558 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_EB06E;
		input reg [1:0] inp;
		sv2v_cast_EB06E = inp;
	endfunction
	always @(posedge clk or negedge rst_n) begin : ID_EX_PIPE_REGISTERS
		// Trace: design.sv:14824:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:14825:7
			alu_en_ex_o <= 1'sb0;
			// Trace: design.sv:14826:7
			alu_operator_ex_o <= sv2v_cast_C07C4(7'b0000011);
			// Trace: design.sv:14827:7
			alu_operand_a_ex_o <= 1'sb0;
			// Trace: design.sv:14828:7
			alu_operand_b_ex_o <= 1'sb0;
			// Trace: design.sv:14829:7
			alu_operand_c_ex_o <= 1'sb0;
			// Trace: design.sv:14830:7
			bmask_a_ex_o <= 1'sb0;
			// Trace: design.sv:14831:7
			bmask_b_ex_o <= 1'sb0;
			// Trace: design.sv:14832:7
			imm_vec_ext_ex_o <= 1'sb0;
			// Trace: design.sv:14833:7
			alu_vec_mode_ex_o <= 1'sb0;
			// Trace: design.sv:14834:7
			alu_clpx_shift_ex_o <= 2'b00;
			// Trace: design.sv:14835:7
			alu_is_clpx_ex_o <= 1'b0;
			// Trace: design.sv:14836:7
			alu_is_subrot_ex_o <= 1'b0;
			// Trace: design.sv:14838:7
			mult_operator_ex_o <= sv2v_cast_9F558(3'b000);
			// Trace: design.sv:14839:7
			mult_operand_a_ex_o <= 1'sb0;
			// Trace: design.sv:14840:7
			mult_operand_b_ex_o <= 1'sb0;
			// Trace: design.sv:14841:7
			mult_operand_c_ex_o <= 1'sb0;
			// Trace: design.sv:14842:7
			mult_en_ex_o <= 1'b0;
			// Trace: design.sv:14843:7
			mult_sel_subword_ex_o <= 1'b0;
			// Trace: design.sv:14844:7
			mult_signed_mode_ex_o <= 2'b00;
			// Trace: design.sv:14845:7
			mult_imm_ex_o <= 1'sb0;
			// Trace: design.sv:14847:7
			mult_dot_op_a_ex_o <= 1'sb0;
			// Trace: design.sv:14848:7
			mult_dot_op_b_ex_o <= 1'sb0;
			// Trace: design.sv:14849:7
			mult_dot_op_c_ex_o <= 1'sb0;
			// Trace: design.sv:14850:7
			mult_dot_signed_ex_o <= 1'sb0;
			// Trace: design.sv:14851:7
			mult_is_clpx_ex_o <= 1'b0;
			// Trace: design.sv:14852:7
			mult_clpx_shift_ex_o <= 2'b00;
			// Trace: design.sv:14853:7
			mult_clpx_img_ex_o <= 1'b0;
			// Trace: design.sv:14855:7
			apu_en_ex_o <= 1'sb0;
			// Trace: design.sv:14856:7
			apu_op_ex_o <= 1'sb0;
			// Trace: design.sv:14857:7
			apu_lat_ex_o <= 1'sb0;
			// Trace: design.sv:14858:7
			apu_operands_ex_o[0+:32] <= 1'sb0;
			// Trace: design.sv:14859:7
			apu_operands_ex_o[32+:32] <= 1'sb0;
			// Trace: design.sv:14860:7
			apu_operands_ex_o[64+:32] <= 1'sb0;
			// Trace: design.sv:14861:7
			apu_flags_ex_o <= 1'sb0;
			// Trace: design.sv:14862:7
			apu_waddr_ex_o <= 1'sb0;
			// Trace: design.sv:14865:7
			regfile_waddr_ex_o <= 6'b000000;
			// Trace: design.sv:14866:7
			regfile_we_ex_o <= 1'b0;
			// Trace: design.sv:14868:7
			regfile_alu_waddr_ex_o <= 6'b000000;
			// Trace: design.sv:14869:7
			regfile_alu_we_ex_o <= 1'b0;
			// Trace: design.sv:14870:7
			prepost_useincr_ex_o <= 1'b0;
			// Trace: design.sv:14872:7
			csr_access_ex_o <= 1'b0;
			// Trace: design.sv:14873:7
			csr_op_ex_o <= sv2v_cast_EB06E(2'b00);
			// Trace: design.sv:14875:7
			data_we_ex_o <= 1'b0;
			// Trace: design.sv:14876:7
			data_type_ex_o <= 2'b00;
			// Trace: design.sv:14877:7
			data_sign_ext_ex_o <= 2'b00;
			// Trace: design.sv:14878:7
			data_reg_offset_ex_o <= 2'b00;
			// Trace: design.sv:14879:7
			data_req_ex_o <= 1'b0;
			// Trace: design.sv:14880:7
			data_load_event_ex_o <= 1'b0;
			// Trace: design.sv:14881:7
			atop_ex_o <= 5'b00000;
			// Trace: design.sv:14883:7
			data_misaligned_ex_o <= 1'b0;
			// Trace: design.sv:14885:7
			pc_ex_o <= 1'sb0;
			// Trace: design.sv:14887:7
			branch_in_ex_o <= 1'b0;
		end
		else if (data_misaligned_i) begin
			begin
				// Trace: design.sv:14891:7
				if (ex_ready_i) begin
					// Trace: design.sv:14896:9
					if (prepost_useincr_ex_o == 1'b1)
						// Trace: design.sv:14897:11
						alu_operand_a_ex_o <= operand_a_fw_id;
					// Trace: design.sv:14900:9
					alu_operand_b_ex_o <= 32'h00000004;
					// Trace: design.sv:14901:9
					regfile_alu_we_ex_o <= 1'b0;
					// Trace: design.sv:14902:9
					prepost_useincr_ex_o <= 1'b1;
					// Trace: design.sv:14904:9
					data_misaligned_ex_o <= 1'b1;
				end
			end
		end
		else if (mult_multicycle_i)
			// Trace: design.sv:14907:7
			mult_operand_c_ex_o <= operand_c_fw_id;
		else
			// Trace: design.sv:14911:7
			if (id_valid_o) begin
				// Trace: design.sv:14912:9
				alu_en_ex_o <= alu_en;
				// Trace: design.sv:14913:9
				if (alu_en) begin
					// Trace: design.sv:14914:11
					alu_operator_ex_o <= alu_operator;
					// Trace: design.sv:14915:11
					alu_operand_a_ex_o <= alu_operand_a;
					// Trace: design.sv:14916:11
					alu_operand_b_ex_o <= alu_operand_b;
					// Trace: design.sv:14917:11
					alu_operand_c_ex_o <= alu_operand_c;
					// Trace: design.sv:14918:11
					bmask_a_ex_o <= bmask_a_id;
					// Trace: design.sv:14919:11
					bmask_b_ex_o <= bmask_b_id;
					// Trace: design.sv:14920:11
					imm_vec_ext_ex_o <= imm_vec_ext_id;
					// Trace: design.sv:14921:11
					alu_vec_mode_ex_o <= alu_vec_mode;
					// Trace: design.sv:14922:11
					alu_is_clpx_ex_o <= is_clpx;
					// Trace: design.sv:14923:11
					alu_clpx_shift_ex_o <= instr[14:13];
					// Trace: design.sv:14924:11
					alu_is_subrot_ex_o <= is_subrot;
				end
				// Trace: design.sv:14927:9
				mult_en_ex_o <= mult_en;
				if (mult_int_en) begin
					// Trace: design.sv:14929:11
					mult_operator_ex_o <= mult_operator;
					// Trace: design.sv:14930:11
					mult_sel_subword_ex_o <= mult_sel_subword;
					// Trace: design.sv:14931:11
					mult_signed_mode_ex_o <= mult_signed_mode;
					// Trace: design.sv:14932:11
					mult_operand_a_ex_o <= alu_operand_a;
					// Trace: design.sv:14933:11
					mult_operand_b_ex_o <= alu_operand_b;
					// Trace: design.sv:14934:11
					mult_operand_c_ex_o <= alu_operand_c;
					// Trace: design.sv:14935:11
					mult_imm_ex_o <= mult_imm_id;
				end
				if (mult_dot_en) begin
					// Trace: design.sv:14938:11
					mult_operator_ex_o <= mult_operator;
					// Trace: design.sv:14939:11
					mult_dot_signed_ex_o <= mult_dot_signed;
					// Trace: design.sv:14940:11
					mult_dot_op_a_ex_o <= alu_operand_a;
					// Trace: design.sv:14941:11
					mult_dot_op_b_ex_o <= alu_operand_b;
					// Trace: design.sv:14942:11
					mult_dot_op_c_ex_o <= alu_operand_c;
					// Trace: design.sv:14943:11
					mult_is_clpx_ex_o <= is_clpx;
					// Trace: design.sv:14944:11
					mult_clpx_shift_ex_o <= instr[14:13];
					// Trace: design.sv:14945:11
					mult_clpx_img_ex_o <= instr[25];
				end
				// Trace: design.sv:14949:9
				apu_en_ex_o <= apu_en;
				if (apu_en) begin
					// Trace: design.sv:14951:11
					apu_op_ex_o <= apu_op;
					// Trace: design.sv:14952:11
					apu_lat_ex_o <= apu_lat;
					// Trace: design.sv:14953:11
					apu_operands_ex_o <= apu_operands;
					// Trace: design.sv:14954:11
					apu_flags_ex_o <= apu_flags;
					// Trace: design.sv:14955:11
					apu_waddr_ex_o <= apu_waddr;
				end
				// Trace: design.sv:14958:9
				regfile_we_ex_o <= regfile_we_id;
				if (regfile_we_id)
					// Trace: design.sv:14960:11
					regfile_waddr_ex_o <= regfile_waddr_id;
				// Trace: design.sv:14963:9
				regfile_alu_we_ex_o <= regfile_alu_we_id;
				if (regfile_alu_we_id)
					// Trace: design.sv:14965:11
					regfile_alu_waddr_ex_o <= regfile_alu_waddr_id;
				// Trace: design.sv:14968:9
				prepost_useincr_ex_o <= prepost_useincr;
				// Trace: design.sv:14970:9
				csr_access_ex_o <= csr_access;
				// Trace: design.sv:14971:9
				csr_op_ex_o <= csr_op;
				// Trace: design.sv:14973:9
				data_req_ex_o <= data_req_id;
				if (data_req_id) begin
					// Trace: design.sv:14975:11
					data_we_ex_o <= data_we_id;
					// Trace: design.sv:14976:11
					data_type_ex_o <= data_type_id;
					// Trace: design.sv:14977:11
					data_sign_ext_ex_o <= data_sign_ext_id;
					// Trace: design.sv:14978:11
					data_reg_offset_ex_o <= data_reg_offset_id;
					// Trace: design.sv:14979:11
					data_load_event_ex_o <= data_load_event_id;
					// Trace: design.sv:14980:11
					atop_ex_o <= atop_id;
				end
				else
					// Trace: design.sv:14982:11
					data_load_event_ex_o <= 1'b0;
				// Trace: design.sv:14985:9
				data_misaligned_ex_o <= 1'b0;
				if ((ctrl_transfer_insn_in_id == cv32e40p_pkg_BRANCH_COND) || data_req_id)
					// Trace: design.sv:14988:11
					pc_ex_o <= pc_id_i;
				// Trace: design.sv:14991:9
				branch_in_ex_o <= ctrl_transfer_insn_in_id == cv32e40p_pkg_BRANCH_COND;
			end
			else if (ex_ready_i) begin
				// Trace: design.sv:14996:9
				regfile_we_ex_o <= 1'b0;
				// Trace: design.sv:14998:9
				regfile_alu_we_ex_o <= 1'b0;
				// Trace: design.sv:15000:9
				csr_op_ex_o <= sv2v_cast_EB06E(2'b00);
				// Trace: design.sv:15002:9
				data_req_ex_o <= 1'b0;
				// Trace: design.sv:15004:9
				data_load_event_ex_o <= 1'b0;
				// Trace: design.sv:15006:9
				data_misaligned_ex_o <= 1'b0;
				// Trace: design.sv:15008:9
				branch_in_ex_o <= 1'b0;
				// Trace: design.sv:15010:9
				apu_en_ex_o <= 1'b0;
				// Trace: design.sv:15012:9
				alu_operator_ex_o <= sv2v_cast_C07C4(7'b0000011);
				// Trace: design.sv:15014:9
				mult_en_ex_o <= 1'b0;
				// Trace: design.sv:15016:9
				alu_en_ex_o <= 1'b1;
			end
			else if (csr_access_ex_o)
				// Trace: design.sv:15022:9
				regfile_alu_we_ex_o <= 1'b0;
	end
	// Trace: design.sv:15032:3
	assign minstret = (id_valid_o && is_decoding_o) && !((illegal_insn_dec || ebrk_insn_dec) || ecall_insn_dec);
	// Trace: design.sv:15034:3
	localparam cv32e40p_pkg_BRANCH_JAL = 2'b01;
	localparam cv32e40p_pkg_BRANCH_JALR = 2'b10;
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:15035:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:15036:7
			id_valid_q <= 1'b0;
			// Trace: design.sv:15037:7
			mhpmevent_minstret_o <= 1'b0;
			// Trace: design.sv:15038:7
			mhpmevent_load_o <= 1'b0;
			// Trace: design.sv:15039:7
			mhpmevent_store_o <= 1'b0;
			// Trace: design.sv:15040:7
			mhpmevent_jump_o <= 1'b0;
			// Trace: design.sv:15041:7
			mhpmevent_branch_o <= 1'b0;
			// Trace: design.sv:15042:7
			mhpmevent_compressed_o <= 1'b0;
			// Trace: design.sv:15043:7
			mhpmevent_branch_taken_o <= 1'b0;
			// Trace: design.sv:15044:7
			mhpmevent_jr_stall_o <= 1'b0;
			// Trace: design.sv:15045:7
			mhpmevent_imiss_o <= 1'b0;
			// Trace: design.sv:15046:7
			mhpmevent_ld_stall_o <= 1'b0;
			// Trace: design.sv:15047:7
			mhpmevent_pipe_stall_o <= 1'b0;
		end
		else begin
			// Trace: design.sv:15050:7
			id_valid_q <= id_valid_o;
			// Trace: design.sv:15052:7
			mhpmevent_minstret_o <= minstret;
			// Trace: design.sv:15053:7
			mhpmevent_load_o <= (minstret && data_req_id) && !data_we_id;
			// Trace: design.sv:15054:7
			mhpmevent_store_o <= (minstret && data_req_id) && data_we_id;
			// Trace: design.sv:15055:7
			mhpmevent_jump_o <= minstret && ((ctrl_transfer_insn_in_id == cv32e40p_pkg_BRANCH_JAL) || (ctrl_transfer_insn_in_id == cv32e40p_pkg_BRANCH_JALR));
			// Trace: design.sv:15056:7
			mhpmevent_branch_o <= minstret && (ctrl_transfer_insn_in_id == cv32e40p_pkg_BRANCH_COND);
			// Trace: design.sv:15057:7
			mhpmevent_compressed_o <= minstret && is_compressed_i;
			// Trace: design.sv:15059:7
			mhpmevent_branch_taken_o <= mhpmevent_branch_o && branch_decision_i;
			// Trace: design.sv:15061:7
			mhpmevent_imiss_o <= perf_imiss_i;
			// Trace: design.sv:15063:7
			mhpmevent_jr_stall_o <= (jr_stall && !halt_id) && id_valid_q;
			// Trace: design.sv:15065:7
			mhpmevent_ld_stall_o <= (load_stall && !halt_id) && id_valid_q;
			// Trace: design.sv:15067:7
			mhpmevent_pipe_stall_o <= perf_pipeline_stall;
		end
	// Trace: design.sv:15072:3
	assign id_ready_o = ((((~misaligned_stall & ~jr_stall) & ~load_stall) & ~apu_stall) & ~csr_apu_stall) & ex_ready_i;
	// Trace: design.sv:15073:3
	assign id_valid_o = ~halt_id & id_ready_o;
	// Trace: design.sv:15074:3
	assign halt_if_o = halt_if;
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_if_stage (
	clk,
	rst_n,
	m_trap_base_addr_i,
	u_trap_base_addr_i,
	trap_addr_mux_i,
	boot_addr_i,
	dm_exception_addr_i,
	dm_halt_addr_i,
	req_i,
	instr_req_o,
	instr_addr_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_rdata_i,
	instr_err_i,
	instr_err_pmp_i,
	instr_valid_id_o,
	instr_rdata_id_o,
	is_compressed_id_o,
	illegal_c_insn_id_o,
	pc_if_o,
	pc_id_o,
	is_fetch_failed_o,
	clear_instr_valid_i,
	pc_set_i,
	mepc_i,
	uepc_i,
	depc_i,
	pc_mux_i,
	exc_pc_mux_i,
	m_exc_vec_pc_mux_i,
	u_exc_vec_pc_mux_i,
	csr_mtvec_init_o,
	jump_target_id_i,
	jump_target_ex_i,
	hwlp_jump_i,
	hwlp_target_i,
	halt_if_i,
	id_ready_i,
	if_busy_o,
	perf_imiss_o
);
	reg _sv2v_0;
	// Trace: design.sv:15258:15
	parameter PULP_XPULP = 0;
	// Trace: design.sv:15259:15
	parameter PULP_OBI = 0;
	// Trace: design.sv:15260:15
	parameter PULP_SECURE = 0;
	// Trace: design.sv:15261:15
	parameter FPU = 0;
	// Trace: design.sv:15263:5
	input wire clk;
	// Trace: design.sv:15264:5
	input wire rst_n;
	// Trace: design.sv:15267:5
	input wire [23:0] m_trap_base_addr_i;
	// Trace: design.sv:15268:5
	input wire [23:0] u_trap_base_addr_i;
	// Trace: design.sv:15269:5
	input wire [1:0] trap_addr_mux_i;
	// Trace: design.sv:15271:5
	input wire [31:0] boot_addr_i;
	// Trace: design.sv:15272:5
	input wire [31:0] dm_exception_addr_i;
	// Trace: design.sv:15275:5
	input wire [31:0] dm_halt_addr_i;
	// Trace: design.sv:15278:5
	input wire req_i;
	// Trace: design.sv:15281:5
	output wire instr_req_o;
	// Trace: design.sv:15282:5
	output wire [31:0] instr_addr_o;
	// Trace: design.sv:15283:5
	input wire instr_gnt_i;
	// Trace: design.sv:15284:5
	input wire instr_rvalid_i;
	// Trace: design.sv:15285:5
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:15286:5
	input wire instr_err_i;
	// Trace: design.sv:15287:5
	input wire instr_err_pmp_i;
	// Trace: design.sv:15290:5
	output reg instr_valid_id_o;
	// Trace: design.sv:15291:5
	output reg [31:0] instr_rdata_id_o;
	// Trace: design.sv:15292:5
	output reg is_compressed_id_o;
	// Trace: design.sv:15293:5
	output reg illegal_c_insn_id_o;
	// Trace: design.sv:15294:5
	output wire [31:0] pc_if_o;
	// Trace: design.sv:15295:5
	output reg [31:0] pc_id_o;
	// Trace: design.sv:15296:5
	output reg is_fetch_failed_o;
	// Trace: design.sv:15299:5
	input wire clear_instr_valid_i;
	// Trace: design.sv:15300:5
	input wire pc_set_i;
	// Trace: design.sv:15301:5
	input wire [31:0] mepc_i;
	// Trace: design.sv:15302:5
	input wire [31:0] uepc_i;
	// Trace: design.sv:15304:5
	input wire [31:0] depc_i;
	// Trace: design.sv:15306:5
	input wire [3:0] pc_mux_i;
	// Trace: design.sv:15307:5
	input wire [2:0] exc_pc_mux_i;
	// Trace: design.sv:15309:5
	input wire [4:0] m_exc_vec_pc_mux_i;
	// Trace: design.sv:15310:5
	input wire [4:0] u_exc_vec_pc_mux_i;
	// Trace: design.sv:15311:5
	output wire csr_mtvec_init_o;
	// Trace: design.sv:15314:5
	input wire [31:0] jump_target_id_i;
	// Trace: design.sv:15315:5
	input wire [31:0] jump_target_ex_i;
	// Trace: design.sv:15318:5
	input wire hwlp_jump_i;
	// Trace: design.sv:15319:5
	input wire [31:0] hwlp_target_i;
	// Trace: design.sv:15322:5
	input wire halt_if_i;
	// Trace: design.sv:15323:5
	input wire id_ready_i;
	// Trace: design.sv:15326:5
	output wire if_busy_o;
	// Trace: design.sv:15327:5
	output wire perf_imiss_o;
	// Trace: design.sv:15330:3
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:15332:3
	wire if_valid;
	wire if_ready;
	// Trace: design.sv:15335:3
	wire prefetch_busy;
	// Trace: design.sv:15336:3
	reg branch_req;
	// Trace: design.sv:15337:3
	reg [31:0] branch_addr_n;
	// Trace: design.sv:15339:3
	wire fetch_valid;
	// Trace: design.sv:15340:3
	reg fetch_ready;
	// Trace: design.sv:15341:3
	wire [31:0] fetch_rdata;
	// Trace: design.sv:15343:3
	reg [31:0] exc_pc;
	// Trace: design.sv:15345:3
	reg [23:0] trap_base_addr;
	// Trace: design.sv:15346:3
	reg [4:0] exc_vec_pc_mux;
	// Trace: design.sv:15347:3
	wire fetch_failed;
	// Trace: design.sv:15349:3
	wire aligner_ready;
	// Trace: design.sv:15350:3
	wire instr_valid;
	// Trace: design.sv:15352:3
	wire illegal_c_insn;
	// Trace: design.sv:15353:3
	wire [31:0] instr_aligned;
	// Trace: design.sv:15354:3
	wire [31:0] instr_decompressed;
	// Trace: design.sv:15355:3
	wire instr_compressed_int;
	// Trace: design.sv:15359:3
	localparam cv32e40p_pkg_EXC_PC_DBD = 3'b010;
	localparam cv32e40p_pkg_EXC_PC_DBE = 3'b011;
	localparam cv32e40p_pkg_EXC_PC_EXCEPTION = 3'b000;
	localparam cv32e40p_pkg_EXC_PC_IRQ = 3'b001;
	localparam cv32e40p_pkg_TRAP_MACHINE = 2'b00;
	localparam cv32e40p_pkg_TRAP_USER = 2'b01;
	always @(*) begin : EXC_PC_MUX
		if (_sv2v_0)
			;
		// Trace: design.sv:15360:5
		(* full_case, parallel_case *)
		case (trap_addr_mux_i)
			cv32e40p_pkg_TRAP_MACHINE:
				// Trace: design.sv:15361:21
				trap_base_addr = m_trap_base_addr_i;
			cv32e40p_pkg_TRAP_USER:
				// Trace: design.sv:15362:21
				trap_base_addr = u_trap_base_addr_i;
			default:
				// Trace: design.sv:15363:21
				trap_base_addr = m_trap_base_addr_i;
		endcase
		(* full_case, parallel_case *)
		case (trap_addr_mux_i)
			cv32e40p_pkg_TRAP_MACHINE:
				// Trace: design.sv:15367:21
				exc_vec_pc_mux = m_exc_vec_pc_mux_i;
			cv32e40p_pkg_TRAP_USER:
				// Trace: design.sv:15368:21
				exc_vec_pc_mux = u_exc_vec_pc_mux_i;
			default:
				// Trace: design.sv:15369:21
				exc_vec_pc_mux = m_exc_vec_pc_mux_i;
		endcase
		(* full_case, parallel_case *)
		case (exc_pc_mux_i)
			cv32e40p_pkg_EXC_PC_EXCEPTION:
				// Trace: design.sv:15374:7
				exc_pc = {trap_base_addr, 8'h00};
			cv32e40p_pkg_EXC_PC_IRQ:
				// Trace: design.sv:15375:19
				exc_pc = {trap_base_addr, 1'b0, exc_vec_pc_mux, 2'b00};
			cv32e40p_pkg_EXC_PC_DBD:
				// Trace: design.sv:15376:19
				exc_pc = {dm_halt_addr_i[31:2], 2'b00};
			cv32e40p_pkg_EXC_PC_DBE:
				// Trace: design.sv:15377:19
				exc_pc = {dm_exception_addr_i[31:2], 2'b00};
			default:
				// Trace: design.sv:15378:16
				exc_pc = {trap_base_addr, 8'h00};
		endcase
	end
	// Trace: design.sv:15383:3
	localparam cv32e40p_pkg_PC_BOOT = 4'b0000;
	localparam cv32e40p_pkg_PC_BRANCH = 4'b0011;
	localparam cv32e40p_pkg_PC_DRET = 4'b0111;
	localparam cv32e40p_pkg_PC_EXCEPTION = 4'b0100;
	localparam cv32e40p_pkg_PC_FENCEI = 4'b0001;
	localparam cv32e40p_pkg_PC_HWLOOP = 4'b1000;
	localparam cv32e40p_pkg_PC_JUMP = 4'b0010;
	localparam cv32e40p_pkg_PC_MRET = 4'b0101;
	localparam cv32e40p_pkg_PC_URET = 4'b0110;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15385:5
		branch_addr_n = {boot_addr_i[31:2], 2'b00};
		// Trace: design.sv:15387:5
		(* full_case, parallel_case *)
		case (pc_mux_i)
			cv32e40p_pkg_PC_BOOT:
				// Trace: design.sv:15388:16
				branch_addr_n = {boot_addr_i[31:2], 2'b00};
			cv32e40p_pkg_PC_JUMP:
				// Trace: design.sv:15389:16
				branch_addr_n = jump_target_id_i;
			cv32e40p_pkg_PC_BRANCH:
				// Trace: design.sv:15390:18
				branch_addr_n = jump_target_ex_i;
			cv32e40p_pkg_PC_EXCEPTION:
				// Trace: design.sv:15391:21
				branch_addr_n = exc_pc;
			cv32e40p_pkg_PC_MRET:
				// Trace: design.sv:15392:16
				branch_addr_n = mepc_i;
			cv32e40p_pkg_PC_URET:
				// Trace: design.sv:15393:16
				branch_addr_n = uepc_i;
			cv32e40p_pkg_PC_DRET:
				// Trace: design.sv:15394:16
				branch_addr_n = depc_i;
			cv32e40p_pkg_PC_FENCEI:
				// Trace: design.sv:15395:18
				branch_addr_n = pc_id_o + 4;
			cv32e40p_pkg_PC_HWLOOP:
				// Trace: design.sv:15396:18
				branch_addr_n = hwlp_target_i;
			default:
				;
		endcase
	end
	// Trace: design.sv:15402:3
	assign csr_mtvec_init_o = (pc_mux_i == cv32e40p_pkg_PC_BOOT) & pc_set_i;
	// Trace: design.sv:15404:3
	assign fetch_failed = 1'b0;
	// Trace: design.sv:15407:3
	cv32e40p_prefetch_buffer #(
		.PULP_OBI(PULP_OBI),
		.PULP_XPULP(PULP_XPULP)
	) prefetch_buffer_i(
		.clk(clk),
		.rst_n(rst_n),
		.req_i(req_i),
		.branch_i(branch_req),
		.branch_addr_i({branch_addr_n[31:1], 1'b0}),
		.hwlp_jump_i(hwlp_jump_i),
		.hwlp_target_i(hwlp_target_i),
		.fetch_ready_i(fetch_ready),
		.fetch_valid_o(fetch_valid),
		.fetch_rdata_o(fetch_rdata),
		.instr_req_o(instr_req_o),
		.instr_addr_o(instr_addr_o),
		.instr_gnt_i(instr_gnt_i),
		.instr_rvalid_i(instr_rvalid_i),
		.instr_err_i(instr_err_i),
		.instr_err_pmp_i(instr_err_pmp_i),
		.instr_rdata_i(instr_rdata_i),
		.busy_o(prefetch_busy)
	);
	// Trace: design.sv:15440:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15442:5
		fetch_ready = 1'b0;
		// Trace: design.sv:15443:5
		branch_req = 1'b0;
		// Trace: design.sv:15445:5
		if (pc_set_i)
			// Trace: design.sv:15446:7
			branch_req = 1'b1;
		else if (fetch_valid) begin
			begin
				// Trace: design.sv:15448:7
				if (req_i && if_valid)
					// Trace: design.sv:15449:9
					fetch_ready = aligner_ready;
			end
		end
	end
	// Trace: design.sv:15454:3
	assign if_busy_o = prefetch_busy;
	// Trace: design.sv:15455:3
	assign perf_imiss_o = !fetch_valid && !branch_req;
	// Trace: design.sv:15458:3
	always @(posedge clk or negedge rst_n) begin : IF_ID_PIPE_REGISTERS
		// Trace: design.sv:15459:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:15460:7
			instr_valid_id_o <= 1'b0;
			// Trace: design.sv:15461:7
			instr_rdata_id_o <= 1'sb0;
			// Trace: design.sv:15462:7
			is_fetch_failed_o <= 1'b0;
			// Trace: design.sv:15463:7
			pc_id_o <= 1'sb0;
			// Trace: design.sv:15464:7
			is_compressed_id_o <= 1'b0;
			// Trace: design.sv:15465:7
			illegal_c_insn_id_o <= 1'b0;
		end
		else
			// Trace: design.sv:15468:7
			if (if_valid && instr_valid) begin
				// Trace: design.sv:15469:9
				instr_valid_id_o <= 1'b1;
				// Trace: design.sv:15470:9
				instr_rdata_id_o <= instr_decompressed;
				// Trace: design.sv:15471:9
				is_compressed_id_o <= instr_compressed_int;
				// Trace: design.sv:15472:9
				illegal_c_insn_id_o <= illegal_c_insn;
				// Trace: design.sv:15473:9
				is_fetch_failed_o <= 1'b0;
				// Trace: design.sv:15474:9
				pc_id_o <= pc_if_o;
			end
			else if (clear_instr_valid_i) begin
				// Trace: design.sv:15476:9
				instr_valid_id_o <= 1'b0;
				// Trace: design.sv:15477:9
				is_fetch_failed_o <= fetch_failed;
			end
	end
	// Trace: design.sv:15482:3
	assign if_ready = fetch_valid & id_ready_i;
	// Trace: design.sv:15483:3
	assign if_valid = ~halt_if_i & if_ready;
	// Trace: design.sv:15485:3
	cv32e40p_aligner aligner_i(
		.clk(clk),
		.rst_n(rst_n),
		.fetch_valid_i(fetch_valid),
		.aligner_ready_o(aligner_ready),
		.if_valid_i(if_valid),
		.fetch_rdata_i(fetch_rdata),
		.instr_aligned_o(instr_aligned),
		.instr_valid_o(instr_valid),
		.branch_addr_i({branch_addr_n[31:1], 1'b0}),
		.branch_i(branch_req),
		.hwlp_addr_i(hwlp_target_i),
		.hwlp_update_pc_i(hwlp_jump_i),
		.pc_o(pc_if_o)
	);
	// Trace: design.sv:15501:3
	cv32e40p_compressed_decoder #(.FPU(FPU)) compressed_decoder_i(
		.instr_i(instr_aligned),
		.instr_o(instr_decompressed),
		.is_compressed_o(instr_compressed_int),
		.illegal_instr_o(illegal_c_insn)
	);
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_load_store_unit (
	clk,
	rst_n,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_err_i,
	data_err_pmp_i,
	data_addr_o,
	data_we_o,
	data_be_o,
	data_wdata_o,
	data_rdata_i,
	data_we_ex_i,
	data_type_ex_i,
	data_wdata_ex_i,
	data_reg_offset_ex_i,
	data_load_event_ex_i,
	data_sign_ext_ex_i,
	data_rdata_ex_o,
	data_req_ex_i,
	operand_a_ex_i,
	operand_b_ex_i,
	addr_useincr_ex_i,
	data_misaligned_ex_i,
	data_misaligned_o,
	data_atop_ex_i,
	data_atop_o,
	p_elw_start_o,
	p_elw_finish_o,
	lsu_ready_ex_o,
	lsu_ready_wb_o,
	busy_o
);
	reg _sv2v_0;
	// Trace: design.sv:15573:15
	parameter PULP_OBI = 0;
	// Trace: design.sv:15575:5
	input wire clk;
	// Trace: design.sv:15576:5
	input wire rst_n;
	// Trace: design.sv:15579:5
	output wire data_req_o;
	// Trace: design.sv:15580:5
	input wire data_gnt_i;
	// Trace: design.sv:15581:5
	input wire data_rvalid_i;
	// Trace: design.sv:15582:5
	input wire data_err_i;
	// Trace: design.sv:15583:5
	input wire data_err_pmp_i;
	// Trace: design.sv:15585:5
	output wire [31:0] data_addr_o;
	// Trace: design.sv:15586:5
	output wire data_we_o;
	// Trace: design.sv:15587:5
	output wire [3:0] data_be_o;
	// Trace: design.sv:15588:5
	output wire [31:0] data_wdata_o;
	// Trace: design.sv:15589:5
	input wire [31:0] data_rdata_i;
	// Trace: design.sv:15592:5
	input wire data_we_ex_i;
	// Trace: design.sv:15593:5
	input wire [1:0] data_type_ex_i;
	// Trace: design.sv:15594:5
	input wire [31:0] data_wdata_ex_i;
	// Trace: design.sv:15595:5
	input wire [1:0] data_reg_offset_ex_i;
	// Trace: design.sv:15596:5
	input wire data_load_event_ex_i;
	// Trace: design.sv:15597:5
	input wire [1:0] data_sign_ext_ex_i;
	// Trace: design.sv:15599:5
	output wire [31:0] data_rdata_ex_o;
	// Trace: design.sv:15600:5
	input wire data_req_ex_i;
	// Trace: design.sv:15601:5
	input wire [31:0] operand_a_ex_i;
	// Trace: design.sv:15602:5
	input wire [31:0] operand_b_ex_i;
	// Trace: design.sv:15603:5
	input wire addr_useincr_ex_i;
	// Trace: design.sv:15605:5
	input wire data_misaligned_ex_i;
	// Trace: design.sv:15606:5
	output reg data_misaligned_o;
	// Trace: design.sv:15608:5
	input wire [5:0] data_atop_ex_i;
	// Trace: design.sv:15609:5
	output wire [5:0] data_atop_o;
	// Trace: design.sv:15611:5
	output wire p_elw_start_o;
	// Trace: design.sv:15612:5
	output wire p_elw_finish_o;
	// Trace: design.sv:15615:5
	output wire lsu_ready_ex_o;
	// Trace: design.sv:15616:5
	output wire lsu_ready_wb_o;
	// Trace: design.sv:15618:5
	output wire busy_o;
	// Trace: design.sv:15621:3
	localparam DEPTH = 2;
	// Trace: design.sv:15624:3
	wire trans_valid;
	// Trace: design.sv:15625:3
	wire trans_ready;
	// Trace: design.sv:15626:3
	wire [31:0] trans_addr;
	// Trace: design.sv:15627:3
	wire trans_we;
	// Trace: design.sv:15628:3
	wire [3:0] trans_be;
	// Trace: design.sv:15629:3
	wire [31:0] trans_wdata;
	// Trace: design.sv:15630:3
	wire [5:0] trans_atop;
	// Trace: design.sv:15633:3
	wire resp_valid;
	// Trace: design.sv:15634:3
	wire [31:0] resp_rdata;
	// Trace: design.sv:15635:3
	wire resp_err;
	// Trace: design.sv:15638:3
	reg [1:0] cnt_q;
	// Trace: design.sv:15639:3
	reg [1:0] next_cnt;
	// Trace: design.sv:15640:3
	wire count_up;
	// Trace: design.sv:15641:3
	wire count_down;
	// Trace: design.sv:15643:3
	wire ctrl_update;
	// Trace: design.sv:15645:3
	wire [31:0] data_addr_int;
	// Trace: design.sv:15648:3
	reg [1:0] data_type_q;
	// Trace: design.sv:15649:3
	reg [1:0] rdata_offset_q;
	// Trace: design.sv:15650:3
	reg [1:0] data_sign_ext_q;
	// Trace: design.sv:15651:3
	reg data_we_q;
	// Trace: design.sv:15652:3
	reg data_load_event_q;
	// Trace: design.sv:15654:3
	wire [1:0] wdata_offset;
	// Trace: design.sv:15656:3
	reg [3:0] data_be;
	// Trace: design.sv:15657:3
	reg [31:0] data_wdata;
	// Trace: design.sv:15659:3
	wire misaligned_st;
	// Trace: design.sv:15660:3
	wire load_err_o;
	wire store_err_o;
	// Trace: design.sv:15662:3
	reg [31:0] rdata_q;
	// Trace: design.sv:15665:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15666:5
		case (data_type_ex_i)
			2'b00:
				// Trace: design.sv:15668:9
				if (misaligned_st == 1'b0)
					// Trace: design.sv:15669:11
					case (data_addr_int[1:0])
						2'b00:
							// Trace: design.sv:15670:20
							data_be = 4'b1111;
						2'b01:
							// Trace: design.sv:15671:20
							data_be = 4'b1110;
						2'b10:
							// Trace: design.sv:15672:20
							data_be = 4'b1100;
						2'b11:
							// Trace: design.sv:15673:20
							data_be = 4'b1000;
					endcase
				else
					// Trace: design.sv:15677:11
					case (data_addr_int[1:0])
						2'b00:
							// Trace: design.sv:15678:20
							data_be = 4'b0000;
						2'b01:
							// Trace: design.sv:15679:20
							data_be = 4'b0001;
						2'b10:
							// Trace: design.sv:15680:20
							data_be = 4'b0011;
						2'b11:
							// Trace: design.sv:15681:20
							data_be = 4'b0111;
					endcase
			2'b01:
				// Trace: design.sv:15688:9
				if (misaligned_st == 1'b0)
					// Trace: design.sv:15689:11
					case (data_addr_int[1:0])
						2'b00:
							// Trace: design.sv:15690:20
							data_be = 4'b0011;
						2'b01:
							// Trace: design.sv:15691:20
							data_be = 4'b0110;
						2'b10:
							// Trace: design.sv:15692:20
							data_be = 4'b1100;
						2'b11:
							// Trace: design.sv:15693:20
							data_be = 4'b1000;
					endcase
				else
					// Trace: design.sv:15697:11
					data_be = 4'b0001;
			2'b10, 2'b11:
				// Trace: design.sv:15702:9
				case (data_addr_int[1:0])
					2'b00:
						// Trace: design.sv:15703:18
						data_be = 4'b0001;
					2'b01:
						// Trace: design.sv:15704:18
						data_be = 4'b0010;
					2'b10:
						// Trace: design.sv:15705:18
						data_be = 4'b0100;
					2'b11:
						// Trace: design.sv:15706:18
						data_be = 4'b1000;
				endcase
		endcase
	end
	// Trace: design.sv:15717:3
	assign wdata_offset = data_addr_int[1:0] - data_reg_offset_ex_i[1:0];
	// Trace: design.sv:15718:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15719:5
		case (wdata_offset)
			2'b00:
				// Trace: design.sv:15720:14
				data_wdata = data_wdata_ex_i[31:0];
			2'b01:
				// Trace: design.sv:15721:14
				data_wdata = {data_wdata_ex_i[23:0], data_wdata_ex_i[31:24]};
			2'b10:
				// Trace: design.sv:15722:14
				data_wdata = {data_wdata_ex_i[15:0], data_wdata_ex_i[31:16]};
			2'b11:
				// Trace: design.sv:15723:14
				data_wdata = {data_wdata_ex_i[7:0], data_wdata_ex_i[31:8]};
		endcase
	end
	// Trace: design.sv:15730:3
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:15731:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:15732:7
			data_type_q <= 1'sb0;
			// Trace: design.sv:15733:7
			rdata_offset_q <= 1'sb0;
			// Trace: design.sv:15734:7
			data_sign_ext_q <= 1'sb0;
			// Trace: design.sv:15735:7
			data_we_q <= 1'b0;
			// Trace: design.sv:15736:7
			data_load_event_q <= 1'b0;
		end
		else if (ctrl_update) begin
			// Trace: design.sv:15740:7
			data_type_q <= data_type_ex_i;
			// Trace: design.sv:15741:7
			rdata_offset_q <= data_addr_int[1:0];
			// Trace: design.sv:15742:7
			data_sign_ext_q <= data_sign_ext_ex_i;
			// Trace: design.sv:15743:7
			data_we_q <= data_we_ex_i;
			// Trace: design.sv:15744:7
			data_load_event_q <= data_load_event_ex_i;
		end
	// Trace: design.sv:15749:3
	assign p_elw_start_o = data_load_event_ex_i && data_req_o;
	// Trace: design.sv:15750:3
	assign p_elw_finish_o = (data_load_event_q && data_rvalid_i) && !data_misaligned_ex_i;
	// Trace: design.sv:15761:3
	reg [31:0] data_rdata_ext;
	// Trace: design.sv:15763:3
	reg [31:0] rdata_w_ext;
	// Trace: design.sv:15764:3
	reg [31:0] rdata_h_ext;
	// Trace: design.sv:15765:3
	reg [31:0] rdata_b_ext;
	// Trace: design.sv:15768:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15769:5
		case (rdata_offset_q)
			2'b00:
				// Trace: design.sv:15770:14
				rdata_w_ext = resp_rdata[31:0];
			2'b01:
				// Trace: design.sv:15771:14
				rdata_w_ext = {resp_rdata[7:0], rdata_q[31:8]};
			2'b10:
				// Trace: design.sv:15772:14
				rdata_w_ext = {resp_rdata[15:0], rdata_q[31:16]};
			2'b11:
				// Trace: design.sv:15773:14
				rdata_w_ext = {resp_rdata[23:0], rdata_q[31:24]};
		endcase
	end
	// Trace: design.sv:15778:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15779:5
		case (rdata_offset_q)
			2'b00:
				// Trace: design.sv:15781:9
				if (data_sign_ext_q == 2'b00)
					// Trace: design.sv:15781:39
					rdata_h_ext = {16'h0000, resp_rdata[15:0]};
				else if (data_sign_ext_q == 2'b10)
					// Trace: design.sv:15782:44
					rdata_h_ext = {16'hffff, resp_rdata[15:0]};
				else
					// Trace: design.sv:15783:14
					rdata_h_ext = {{16 {resp_rdata[15]}}, resp_rdata[15:0]};
			2'b01:
				// Trace: design.sv:15787:9
				if (data_sign_ext_q == 2'b00)
					// Trace: design.sv:15787:39
					rdata_h_ext = {16'h0000, resp_rdata[23:8]};
				else if (data_sign_ext_q == 2'b10)
					// Trace: design.sv:15788:44
					rdata_h_ext = {16'hffff, resp_rdata[23:8]};
				else
					// Trace: design.sv:15789:14
					rdata_h_ext = {{16 {resp_rdata[23]}}, resp_rdata[23:8]};
			2'b10:
				// Trace: design.sv:15793:9
				if (data_sign_ext_q == 2'b00)
					// Trace: design.sv:15793:39
					rdata_h_ext = {16'h0000, resp_rdata[31:16]};
				else if (data_sign_ext_q == 2'b10)
					// Trace: design.sv:15794:44
					rdata_h_ext = {16'hffff, resp_rdata[31:16]};
				else
					// Trace: design.sv:15795:14
					rdata_h_ext = {{16 {resp_rdata[31]}}, resp_rdata[31:16]};
			2'b11:
				// Trace: design.sv:15799:9
				if (data_sign_ext_q == 2'b00)
					// Trace: design.sv:15799:39
					rdata_h_ext = {16'h0000, resp_rdata[7:0], rdata_q[31:24]};
				else if (data_sign_ext_q == 2'b10)
					// Trace: design.sv:15801:11
					rdata_h_ext = {16'hffff, resp_rdata[7:0], rdata_q[31:24]};
				else
					// Trace: design.sv:15802:14
					rdata_h_ext = {{16 {resp_rdata[7]}}, resp_rdata[7:0], rdata_q[31:24]};
		endcase
	end
	// Trace: design.sv:15808:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15809:5
		case (rdata_offset_q)
			2'b00:
				// Trace: design.sv:15811:9
				if (data_sign_ext_q == 2'b00)
					// Trace: design.sv:15811:39
					rdata_b_ext = {24'h000000, resp_rdata[7:0]};
				else if (data_sign_ext_q == 2'b10)
					// Trace: design.sv:15812:44
					rdata_b_ext = {24'hffffff, resp_rdata[7:0]};
				else
					// Trace: design.sv:15813:14
					rdata_b_ext = {{24 {resp_rdata[7]}}, resp_rdata[7:0]};
			2'b01:
				// Trace: design.sv:15817:9
				if (data_sign_ext_q == 2'b00)
					// Trace: design.sv:15817:39
					rdata_b_ext = {24'h000000, resp_rdata[15:8]};
				else if (data_sign_ext_q == 2'b10)
					// Trace: design.sv:15818:44
					rdata_b_ext = {24'hffffff, resp_rdata[15:8]};
				else
					// Trace: design.sv:15819:14
					rdata_b_ext = {{24 {resp_rdata[15]}}, resp_rdata[15:8]};
			2'b10:
				// Trace: design.sv:15823:9
				if (data_sign_ext_q == 2'b00)
					// Trace: design.sv:15823:39
					rdata_b_ext = {24'h000000, resp_rdata[23:16]};
				else if (data_sign_ext_q == 2'b10)
					// Trace: design.sv:15824:44
					rdata_b_ext = {24'hffffff, resp_rdata[23:16]};
				else
					// Trace: design.sv:15825:14
					rdata_b_ext = {{24 {resp_rdata[23]}}, resp_rdata[23:16]};
			2'b11:
				// Trace: design.sv:15829:9
				if (data_sign_ext_q == 2'b00)
					// Trace: design.sv:15829:39
					rdata_b_ext = {24'h000000, resp_rdata[31:24]};
				else if (data_sign_ext_q == 2'b10)
					// Trace: design.sv:15830:44
					rdata_b_ext = {24'hffffff, resp_rdata[31:24]};
				else
					// Trace: design.sv:15831:14
					rdata_b_ext = {{24 {resp_rdata[31]}}, resp_rdata[31:24]};
		endcase
	end
	// Trace: design.sv:15837:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15838:5
		case (data_type_q)
			2'b00:
				// Trace: design.sv:15839:21
				data_rdata_ext = rdata_w_ext;
			2'b01:
				// Trace: design.sv:15840:21
				data_rdata_ext = rdata_h_ext;
			2'b10, 2'b11:
				// Trace: design.sv:15841:21
				data_rdata_ext = rdata_b_ext;
		endcase
	end
	// Trace: design.sv:15845:3
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:15846:5
		if (rst_n == 1'b0)
			// Trace: design.sv:15847:7
			rdata_q <= 1'sb0;
		else
			// Trace: design.sv:15849:7
			if (resp_valid && ~data_we_q) begin
				begin
					// Trace: design.sv:15855:9
					if ((data_misaligned_ex_i == 1'b1) || (data_misaligned_o == 1'b1))
						// Trace: design.sv:15855:76
						rdata_q <= resp_rdata;
					else
						// Trace: design.sv:15856:14
						rdata_q <= data_rdata_ext;
				end
			end
	// Trace: design.sv:15862:3
	assign data_rdata_ex_o = (resp_valid == 1'b1 ? data_rdata_ext : rdata_q);
	// Trace: design.sv:15864:3
	assign misaligned_st = data_misaligned_ex_i;
	// Trace: design.sv:15867:3
	assign load_err_o = (data_gnt_i && data_err_pmp_i) && ~data_we_o;
	// Trace: design.sv:15868:3
	assign store_err_o = (data_gnt_i && data_err_pmp_i) && data_we_o;
	// Trace: design.sv:15874:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15875:5
		data_misaligned_o = 1'b0;
		// Trace: design.sv:15877:5
		if ((data_req_ex_i == 1'b1) && (data_misaligned_ex_i == 1'b0))
			// Trace: design.sv:15878:7
			case (data_type_ex_i)
				2'b00:
					// Trace: design.sv:15881:11
					if (data_addr_int[1:0] != 2'b00)
						// Trace: design.sv:15881:44
						data_misaligned_o = 1'b1;
				2'b01:
					// Trace: design.sv:15885:11
					if (data_addr_int[1:0] == 2'b11)
						// Trace: design.sv:15885:44
						data_misaligned_o = 1'b1;
			endcase
	end
	// Trace: design.sv:15892:3
	assign data_addr_int = (addr_useincr_ex_i ? operand_a_ex_i + operand_b_ex_i : operand_a_ex_i);
	// Trace: design.sv:15895:3
	assign busy_o = (cnt_q != 2'b00) || trans_valid;
	// Trace: design.sv:15907:3
	assign trans_addr = (data_misaligned_ex_i ? {data_addr_int[31:2], 2'b00} : data_addr_int);
	// Trace: design.sv:15908:3
	assign trans_we = data_we_ex_i;
	// Trace: design.sv:15909:3
	assign trans_be = data_be;
	// Trace: design.sv:15910:3
	assign trans_wdata = data_wdata;
	// Trace: design.sv:15911:3
	assign trans_atop = data_atop_ex_i;
	// Trace: design.sv:15914:3
	generate
		if (PULP_OBI == 0) begin : gen_no_pulp_obi
			// Trace: design.sv:15919:7
			assign trans_valid = data_req_ex_i && (cnt_q < DEPTH);
		end
		else begin : gen_pulp_obi
			// Trace: design.sv:15923:7
			assign trans_valid = (cnt_q == 2'b00 ? data_req_ex_i && (cnt_q < DEPTH) : (data_req_ex_i && (cnt_q < DEPTH)) && resp_valid);
		end
	endgenerate
	// Trace: design.sv:15930:3
	assign lsu_ready_wb_o = (cnt_q == 2'b00 ? 1'b1 : resp_valid);
	// Trace: design.sv:15943:3
	assign lsu_ready_ex_o = (data_req_ex_i == 1'b0 ? 1'b1 : (cnt_q == 2'b00 ? trans_valid && trans_ready : (cnt_q == 2'b01 ? (resp_valid && trans_valid) && trans_ready : resp_valid)));
	// Trace: design.sv:15949:3
	assign ctrl_update = lsu_ready_ex_o && data_req_ex_i;
	// Trace: design.sv:15961:3
	assign count_up = trans_valid && trans_ready;
	// Trace: design.sv:15962:3
	assign count_down = resp_valid;
	// Trace: design.sv:15964:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:15965:5
		(* full_case, parallel_case *)
		case ({count_up, count_down})
			2'b00:
				// Trace: design.sv:15969:9
				next_cnt = cnt_q;
			2'b01:
				// Trace: design.sv:15972:9
				next_cnt = cnt_q - 1'b1;
			2'b10:
				// Trace: design.sv:15975:9
				next_cnt = cnt_q + 1'b1;
			2'b11:
				// Trace: design.sv:15978:9
				next_cnt = cnt_q;
		endcase
	end
	// Trace: design.sv:15988:3
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:15989:5
		if (rst_n == 1'b0)
			// Trace: design.sv:15990:7
			cnt_q <= 1'sb0;
		else
			// Trace: design.sv:15992:7
			cnt_q <= next_cnt;
	// Trace: design.sv:16001:3
	cv32e40p_obi_interface #(.TRANS_STABLE(1)) data_obi_i(
		.clk(clk),
		.rst_n(rst_n),
		.trans_valid_i(trans_valid),
		.trans_ready_o(trans_ready),
		.trans_addr_i(trans_addr),
		.trans_we_i(trans_we),
		.trans_be_i(trans_be),
		.trans_wdata_i(trans_wdata),
		.trans_atop_i(trans_atop),
		.resp_valid_o(resp_valid),
		.resp_rdata_o(resp_rdata),
		.resp_err_o(resp_err),
		.obi_req_o(data_req_o),
		.obi_gnt_i(data_gnt_i),
		.obi_addr_o(data_addr_o),
		.obi_we_o(data_we_o),
		.obi_be_o(data_be_o),
		.obi_wdata_o(data_wdata_o),
		.obi_atop_o(data_atop_o),
		.obi_rdata_i(data_rdata_i),
		.obi_rvalid_i(data_rvalid_i),
		.obi_err_i(data_err_i)
	);
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_mult (
	clk,
	rst_n,
	enable_i,
	operator_i,
	short_subword_i,
	short_signed_i,
	op_a_i,
	op_b_i,
	op_c_i,
	imm_i,
	dot_signed_i,
	dot_op_a_i,
	dot_op_b_i,
	dot_op_c_i,
	is_clpx_i,
	clpx_shift_i,
	clpx_img_i,
	result_o,
	multicycle_o,
	ready_o,
	ex_ready_i
);
	reg _sv2v_0;
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:16124:5
	input wire clk;
	// Trace: design.sv:16125:5
	input wire rst_n;
	// Trace: design.sv:16127:5
	input wire enable_i;
	// Trace: design.sv:16128:5
	localparam cv32e40p_pkg_MUL_OP_WIDTH = 3;
	// removed localparam type cv32e40p_pkg_mul_opcode_e
	input wire [2:0] operator_i;
	// Trace: design.sv:16131:5
	input wire short_subword_i;
	// Trace: design.sv:16132:5
	input wire [1:0] short_signed_i;
	// Trace: design.sv:16134:5
	input wire [31:0] op_a_i;
	// Trace: design.sv:16135:5
	input wire [31:0] op_b_i;
	// Trace: design.sv:16136:5
	input wire [31:0] op_c_i;
	// Trace: design.sv:16138:5
	input wire [4:0] imm_i;
	// Trace: design.sv:16142:5
	input wire [1:0] dot_signed_i;
	// Trace: design.sv:16143:5
	input wire [31:0] dot_op_a_i;
	// Trace: design.sv:16144:5
	input wire [31:0] dot_op_b_i;
	// Trace: design.sv:16145:5
	input wire [31:0] dot_op_c_i;
	// Trace: design.sv:16146:5
	input wire is_clpx_i;
	// Trace: design.sv:16147:5
	input wire [1:0] clpx_shift_i;
	// Trace: design.sv:16148:5
	input wire clpx_img_i;
	// Trace: design.sv:16150:5
	output reg [31:0] result_o;
	// Trace: design.sv:16152:5
	output reg multicycle_o;
	// Trace: design.sv:16153:5
	output wire ready_o;
	// Trace: design.sv:16154:5
	input wire ex_ready_i;
	// Trace: design.sv:16165:3
	wire [16:0] short_op_a;
	// Trace: design.sv:16166:3
	wire [16:0] short_op_b;
	// Trace: design.sv:16167:3
	wire [32:0] short_op_c;
	// Trace: design.sv:16168:3
	wire [33:0] short_mul;
	// Trace: design.sv:16169:3
	wire [33:0] short_mac;
	// Trace: design.sv:16170:3
	wire [31:0] short_round;
	wire [31:0] short_round_tmp;
	// Trace: design.sv:16171:3
	wire [33:0] short_result;
	// Trace: design.sv:16173:3
	wire short_mac_msb1;
	// Trace: design.sv:16174:3
	wire short_mac_msb0;
	// Trace: design.sv:16176:3
	wire [4:0] short_imm;
	// Trace: design.sv:16177:3
	wire [1:0] short_subword;
	// Trace: design.sv:16178:3
	wire [1:0] short_signed;
	// Trace: design.sv:16179:3
	wire short_shift_arith;
	// Trace: design.sv:16180:3
	reg [4:0] mulh_imm;
	// Trace: design.sv:16181:3
	reg [1:0] mulh_subword;
	// Trace: design.sv:16182:3
	reg [1:0] mulh_signed;
	// Trace: design.sv:16183:3
	reg mulh_shift_arith;
	// Trace: design.sv:16184:3
	reg mulh_carry_q;
	// Trace: design.sv:16185:3
	reg mulh_active;
	// Trace: design.sv:16186:3
	reg mulh_save;
	// Trace: design.sv:16187:3
	reg mulh_clearcarry;
	// Trace: design.sv:16188:3
	reg mulh_ready;
	// Trace: design.sv:16190:3
	// removed localparam type cv32e40p_pkg_mult_state_e
	reg [2:0] mulh_CS;
	reg [2:0] mulh_NS;
	// Trace: design.sv:16193:3
	assign short_round_tmp = 32'h00000001 << imm_i;
	// Trace: design.sv:16194:3
	function automatic [2:0] sv2v_cast_9F558;
		input reg [2:0] inp;
		sv2v_cast_9F558 = inp;
	endfunction
	assign short_round = (operator_i == sv2v_cast_9F558(3'b011) ? {1'b0, short_round_tmp[31:1]} : {32 {1'sb0}});
	// Trace: design.sv:16197:3
	assign short_op_a[15:0] = (short_subword[0] ? op_a_i[31:16] : op_a_i[15:0]);
	// Trace: design.sv:16198:3
	assign short_op_b[15:0] = (short_subword[1] ? op_b_i[31:16] : op_b_i[15:0]);
	// Trace: design.sv:16200:3
	assign short_op_a[16] = short_signed[0] & short_op_a[15];
	// Trace: design.sv:16201:3
	assign short_op_b[16] = short_signed[1] & short_op_b[15];
	// Trace: design.sv:16203:3
	assign short_op_c = (mulh_active ? $signed({mulh_carry_q, op_c_i}) : $signed(op_c_i));
	// Trace: design.sv:16205:3
	assign short_mul = $signed(short_op_a) * $signed(short_op_b);
	// Trace: design.sv:16206:3
	assign short_mac = ($signed(short_op_c) + $signed(short_mul)) + $signed(short_round);
	// Trace: design.sv:16209:3
	assign short_result = $signed({short_shift_arith & short_mac_msb1, short_shift_arith & short_mac_msb0, short_mac[31:0]}) >>> short_imm;
	// Trace: design.sv:16214:3
	assign short_imm = (mulh_active ? mulh_imm : imm_i);
	// Trace: design.sv:16215:3
	assign short_subword = (mulh_active ? mulh_subword : {2 {short_subword_i}});
	// Trace: design.sv:16216:3
	assign short_signed = (mulh_active ? mulh_signed : short_signed_i);
	// Trace: design.sv:16217:3
	assign short_shift_arith = (mulh_active ? mulh_shift_arith : short_signed_i[0]);
	// Trace: design.sv:16219:3
	assign short_mac_msb1 = (mulh_active ? short_mac[33] : short_mac[31]);
	// Trace: design.sv:16220:3
	assign short_mac_msb0 = (mulh_active ? short_mac[32] : short_mac[31]);
	// Trace: design.sv:16223:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:16224:5
		mulh_NS = mulh_CS;
		// Trace: design.sv:16225:5
		mulh_imm = 5'd0;
		// Trace: design.sv:16226:5
		mulh_subword = 2'b00;
		// Trace: design.sv:16227:5
		mulh_signed = 2'b00;
		// Trace: design.sv:16228:5
		mulh_shift_arith = 1'b0;
		// Trace: design.sv:16229:5
		mulh_ready = 1'b0;
		// Trace: design.sv:16230:5
		mulh_active = 1'b1;
		// Trace: design.sv:16231:5
		mulh_save = 1'b0;
		// Trace: design.sv:16232:5
		mulh_clearcarry = 1'b0;
		// Trace: design.sv:16233:5
		multicycle_o = 1'b0;
		// Trace: design.sv:16235:5
		case (mulh_CS)
			3'd0: begin
				// Trace: design.sv:16237:9
				mulh_active = 1'b0;
				// Trace: design.sv:16238:9
				mulh_ready = 1'b1;
				// Trace: design.sv:16239:9
				mulh_save = 1'b0;
				// Trace: design.sv:16240:9
				if ((operator_i == sv2v_cast_9F558(3'b110)) && enable_i) begin
					// Trace: design.sv:16241:11
					mulh_ready = 1'b0;
					// Trace: design.sv:16242:11
					mulh_NS = 3'd1;
				end
			end
			3'd1: begin
				// Trace: design.sv:16247:9
				multicycle_o = 1'b1;
				// Trace: design.sv:16248:9
				mulh_imm = 5'd16;
				// Trace: design.sv:16249:9
				mulh_active = 1'b1;
				// Trace: design.sv:16251:9
				mulh_save = 1'b0;
				// Trace: design.sv:16252:9
				mulh_NS = 3'd2;
			end
			3'd2: begin
				// Trace: design.sv:16257:9
				multicycle_o = 1'b1;
				// Trace: design.sv:16259:9
				mulh_signed = {short_signed_i[1], 1'b0};
				// Trace: design.sv:16260:9
				mulh_subword = 2'b10;
				// Trace: design.sv:16261:9
				mulh_save = 1'b1;
				// Trace: design.sv:16262:9
				mulh_shift_arith = 1'b1;
				// Trace: design.sv:16263:9
				mulh_NS = 3'd3;
			end
			3'd3: begin
				// Trace: design.sv:16271:9
				multicycle_o = 1'b1;
				// Trace: design.sv:16273:9
				mulh_signed = {1'b0, short_signed_i[0]};
				// Trace: design.sv:16274:9
				mulh_subword = 2'b01;
				// Trace: design.sv:16275:9
				mulh_imm = 5'd16;
				// Trace: design.sv:16276:9
				mulh_save = 1'b1;
				// Trace: design.sv:16277:9
				mulh_clearcarry = 1'b1;
				// Trace: design.sv:16278:9
				mulh_shift_arith = 1'b1;
				// Trace: design.sv:16279:9
				mulh_NS = 3'd4;
			end
			3'd4: begin
				// Trace: design.sv:16286:9
				mulh_signed = short_signed_i;
				// Trace: design.sv:16287:9
				mulh_subword = 2'b11;
				// Trace: design.sv:16288:9
				mulh_ready = 1'b1;
				// Trace: design.sv:16289:9
				if (ex_ready_i)
					// Trace: design.sv:16289:25
					mulh_NS = 3'd0;
			end
		endcase
	end
	// Trace: design.sv:16294:3
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:16295:5
		if (~rst_n) begin
			// Trace: design.sv:16296:7
			mulh_CS <= 3'd0;
			// Trace: design.sv:16297:7
			mulh_carry_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:16299:7
			mulh_CS <= mulh_NS;
			// Trace: design.sv:16301:7
			if (mulh_save)
				// Trace: design.sv:16301:22
				mulh_carry_q <= ~mulh_clearcarry & short_mac[32];
			else if (ex_ready_i)
				// Trace: design.sv:16303:9
				mulh_carry_q <= 1'b0;
		end
	// Trace: design.sv:16308:3
	wire [31:0] int_op_a_msu;
	// Trace: design.sv:16309:3
	wire [31:0] int_op_b_msu;
	// Trace: design.sv:16310:3
	wire [31:0] int_result;
	// Trace: design.sv:16312:3
	wire int_is_msu;
	// Trace: design.sv:16314:3
	assign int_is_msu = operator_i == sv2v_cast_9F558(3'b001);
	// Trace: design.sv:16316:3
	assign int_op_a_msu = op_a_i ^ {32 {int_is_msu}};
	// Trace: design.sv:16317:3
	assign int_op_b_msu = op_b_i & {32 {int_is_msu}};
	// Trace: design.sv:16319:3
	assign int_result = ($signed(op_c_i) + $signed(int_op_b_msu)) + ($signed(int_op_a_msu) * $signed(op_b_i));
	// Trace: design.sv:16337:3
	wire [31:0] dot_char_result;
	// Trace: design.sv:16338:3
	wire [32:0] dot_short_result;
	// Trace: design.sv:16339:3
	wire [31:0] accumulator;
	// Trace: design.sv:16340:3
	wire [15:0] clpx_shift_result;
	// Trace: design.sv:16341:3
	wire [35:0] dot_char_op_a;
	// Trace: design.sv:16342:3
	wire [35:0] dot_char_op_b;
	// Trace: design.sv:16343:3
	wire [71:0] dot_char_mul;
	// Trace: design.sv:16345:3
	wire [33:0] dot_short_op_a;
	// Trace: design.sv:16346:3
	wire [33:0] dot_short_op_b;
	// Trace: design.sv:16347:3
	wire [67:0] dot_short_mul;
	// Trace: design.sv:16348:3
	wire [16:0] dot_short_op_a_1_neg;
	// Trace: design.sv:16349:3
	wire [31:0] dot_short_op_b_ext;
	// Trace: design.sv:16351:3
	assign dot_char_op_a[0+:9] = {dot_signed_i[1] & dot_op_a_i[7], dot_op_a_i[7:0]};
	// Trace: design.sv:16352:3
	assign dot_char_op_a[9+:9] = {dot_signed_i[1] & dot_op_a_i[15], dot_op_a_i[15:8]};
	// Trace: design.sv:16353:3
	assign dot_char_op_a[18+:9] = {dot_signed_i[1] & dot_op_a_i[23], dot_op_a_i[23:16]};
	// Trace: design.sv:16354:3
	assign dot_char_op_a[27+:9] = {dot_signed_i[1] & dot_op_a_i[31], dot_op_a_i[31:24]};
	// Trace: design.sv:16356:3
	assign dot_char_op_b[0+:9] = {dot_signed_i[0] & dot_op_b_i[7], dot_op_b_i[7:0]};
	// Trace: design.sv:16357:3
	assign dot_char_op_b[9+:9] = {dot_signed_i[0] & dot_op_b_i[15], dot_op_b_i[15:8]};
	// Trace: design.sv:16358:3
	assign dot_char_op_b[18+:9] = {dot_signed_i[0] & dot_op_b_i[23], dot_op_b_i[23:16]};
	// Trace: design.sv:16359:3
	assign dot_char_op_b[27+:9] = {dot_signed_i[0] & dot_op_b_i[31], dot_op_b_i[31:24]};
	// Trace: design.sv:16361:3
	assign dot_char_mul[0+:18] = $signed(dot_char_op_a[0+:9]) * $signed(dot_char_op_b[0+:9]);
	// Trace: design.sv:16362:3
	assign dot_char_mul[18+:18] = $signed(dot_char_op_a[9+:9]) * $signed(dot_char_op_b[9+:9]);
	// Trace: design.sv:16363:3
	assign dot_char_mul[36+:18] = $signed(dot_char_op_a[18+:9]) * $signed(dot_char_op_b[18+:9]);
	// Trace: design.sv:16364:3
	assign dot_char_mul[54+:18] = $signed(dot_char_op_a[27+:9]) * $signed(dot_char_op_b[27+:9]);
	// Trace: design.sv:16366:3
	assign dot_char_result = ((($signed(dot_char_mul[0+:18]) + $signed(dot_char_mul[18+:18])) + $signed(dot_char_mul[36+:18])) + $signed(dot_char_mul[54+:18])) + $signed(dot_op_c_i);
	// Trace: design.sv:16379:3
	assign dot_short_op_a[0+:17] = {dot_signed_i[1] & dot_op_a_i[15], dot_op_a_i[15:0]};
	// Trace: design.sv:16380:3
	assign dot_short_op_a[17+:17] = {dot_signed_i[1] & dot_op_a_i[31], dot_op_a_i[31:16]};
	// Trace: design.sv:16381:3
	assign dot_short_op_a_1_neg = dot_short_op_a[17+:17] ^ {17 {is_clpx_i & ~clpx_img_i}};
	// Trace: design.sv:16383:3
	assign dot_short_op_b[0+:17] = (is_clpx_i & clpx_img_i ? {dot_signed_i[0] & dot_op_b_i[31], dot_op_b_i[31:16]} : {dot_signed_i[0] & dot_op_b_i[15], dot_op_b_i[15:0]});
	// Trace: design.sv:16388:3
	assign dot_short_op_b[17+:17] = (is_clpx_i & clpx_img_i ? {dot_signed_i[0] & dot_op_b_i[15], dot_op_b_i[15:0]} : {dot_signed_i[0] & dot_op_b_i[31], dot_op_b_i[31:16]});
	// Trace: design.sv:16394:3
	assign dot_short_mul[0+:34] = $signed(dot_short_op_a[0+:17]) * $signed(dot_short_op_b[0+:17]);
	// Trace: design.sv:16395:3
	assign dot_short_mul[34+:34] = $signed(dot_short_op_a_1_neg) * $signed(dot_short_op_b[17+:17]);
	// Trace: design.sv:16397:3
	assign dot_short_op_b_ext = $signed(dot_short_op_b[17+:17]);
	// Trace: design.sv:16398:3
	assign accumulator = (is_clpx_i ? dot_short_op_b_ext & {32 {~clpx_img_i}} : $signed(dot_op_c_i));
	// Trace: design.sv:16400:3
	assign dot_short_result = ($signed(dot_short_mul[31-:32]) + $signed(dot_short_mul[65-:32])) + $signed(accumulator);
	// Trace: design.sv:16407:3
	assign clpx_shift_result = $signed(dot_short_result[31:15]) >>> clpx_shift_i;
	// Trace: design.sv:16418:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:16419:5
		result_o = 1'sb0;
		// Trace: design.sv:16421:5
		(* full_case, parallel_case *)
		case (operator_i)
			sv2v_cast_9F558(3'b000), sv2v_cast_9F558(3'b001):
				// Trace: design.sv:16422:29
				result_o = int_result[31:0];
			sv2v_cast_9F558(3'b010), sv2v_cast_9F558(3'b011), sv2v_cast_9F558(3'b110):
				// Trace: design.sv:16424:29
				result_o = short_result[31:0];
			sv2v_cast_9F558(3'b100):
				// Trace: design.sv:16426:17
				result_o = dot_char_result[31:0];
			sv2v_cast_9F558(3'b101):
				// Trace: design.sv:16428:9
				if (is_clpx_i) begin
					begin
						// Trace: design.sv:16429:11
						if (clpx_img_i) begin
							// Trace: design.sv:16430:13
							result_o[31:16] = clpx_shift_result;
							// Trace: design.sv:16431:13
							result_o[15:0] = dot_op_c_i[15:0];
						end
						else begin
							// Trace: design.sv:16433:13
							result_o[15:0] = clpx_shift_result;
							// Trace: design.sv:16434:13
							result_o[31:16] = dot_op_c_i[31:16];
						end
					end
				end
				else
					// Trace: design.sv:16437:11
					result_o = dot_short_result[31:0];
			default:
				;
		endcase
	end
	// Trace: design.sv:16445:3
	assign ready_o = mulh_ready;
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_prefetch_buffer (
	clk,
	rst_n,
	req_i,
	branch_i,
	branch_addr_i,
	hwlp_jump_i,
	hwlp_target_i,
	fetch_ready_i,
	fetch_valid_o,
	fetch_rdata_o,
	instr_req_o,
	instr_gnt_i,
	instr_addr_o,
	instr_rdata_i,
	instr_rvalid_i,
	instr_err_i,
	instr_err_pmp_i,
	busy_o
);
	// Trace: design.sv:16510:15
	parameter PULP_OBI = 0;
	// Trace: design.sv:16511:15
	parameter PULP_XPULP = 1;
	// Trace: design.sv:16513:5
	input wire clk;
	// Trace: design.sv:16514:5
	input wire rst_n;
	// Trace: design.sv:16516:5
	input wire req_i;
	// Trace: design.sv:16517:5
	input wire branch_i;
	// Trace: design.sv:16518:5
	input wire [31:0] branch_addr_i;
	// Trace: design.sv:16520:5
	input wire hwlp_jump_i;
	// Trace: design.sv:16521:5
	input wire [31:0] hwlp_target_i;
	// Trace: design.sv:16523:5
	input wire fetch_ready_i;
	// Trace: design.sv:16524:5
	output wire fetch_valid_o;
	// Trace: design.sv:16525:5
	output wire [31:0] fetch_rdata_o;
	// Trace: design.sv:16528:5
	output wire instr_req_o;
	// Trace: design.sv:16529:5
	input wire instr_gnt_i;
	// Trace: design.sv:16530:5
	output wire [31:0] instr_addr_o;
	// Trace: design.sv:16531:5
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:16532:5
	input wire instr_rvalid_i;
	// Trace: design.sv:16533:5
	input wire instr_err_i;
	// Trace: design.sv:16534:5
	input wire instr_err_pmp_i;
	// Trace: design.sv:16537:5
	output wire busy_o;
	// Trace: design.sv:16542:3
	localparam FIFO_DEPTH = 2;
	// Trace: design.sv:16543:3
	localparam [31:0] FIFO_ADDR_DEPTH = 1;
	// Trace: design.sv:16546:3
	wire trans_valid;
	// Trace: design.sv:16547:3
	wire trans_ready;
	// Trace: design.sv:16548:3
	wire [31:0] trans_addr;
	// Trace: design.sv:16550:3
	wire fifo_flush;
	// Trace: design.sv:16551:3
	wire fifo_flush_but_first;
	// Trace: design.sv:16552:3
	wire [FIFO_ADDR_DEPTH:0] fifo_cnt;
	// Trace: design.sv:16554:3
	wire [31:0] fifo_rdata;
	// Trace: design.sv:16555:3
	wire fifo_push;
	// Trace: design.sv:16556:3
	wire fifo_pop;
	// Trace: design.sv:16557:3
	wire fifo_empty;
	// Trace: design.sv:16560:3
	wire resp_valid;
	// Trace: design.sv:16561:3
	wire [31:0] resp_rdata;
	// Trace: design.sv:16562:3
	wire resp_err;
	// Trace: design.sv:16568:3
	cv32e40p_prefetch_controller #(
		.DEPTH(FIFO_DEPTH),
		.PULP_OBI(PULP_OBI),
		.PULP_XPULP(PULP_XPULP)
	) prefetch_controller_i(
		.clk(clk),
		.rst_n(rst_n),
		.req_i(req_i),
		.branch_i(branch_i),
		.branch_addr_i(branch_addr_i),
		.busy_o(busy_o),
		.hwlp_jump_i(hwlp_jump_i),
		.hwlp_target_i(hwlp_target_i),
		.trans_valid_o(trans_valid),
		.trans_ready_i(trans_ready),
		.trans_addr_o(trans_addr),
		.resp_valid_i(resp_valid),
		.fetch_ready_i(fetch_ready_i),
		.fetch_valid_o(fetch_valid_o),
		.fifo_push_o(fifo_push),
		.fifo_pop_o(fifo_pop),
		.fifo_flush_o(fifo_flush),
		.fifo_flush_but_first_o(fifo_flush_but_first),
		.fifo_cnt_i(fifo_cnt),
		.fifo_empty_i(fifo_empty)
	);
	// Trace: design.sv:16605:3
	cv32e40p_fifo #(
		.FALL_THROUGH(1'b0),
		.DATA_WIDTH(32),
		.DEPTH(FIFO_DEPTH)
	) fifo_i(
		.clk_i(clk),
		.rst_ni(rst_n),
		.flush_i(fifo_flush),
		.flush_but_first_i(fifo_flush_but_first),
		.testmode_i(1'b0),
		.full_o(),
		.empty_o(fifo_empty),
		.cnt_o(fifo_cnt),
		.data_i(resp_rdata),
		.push_i(fifo_push),
		.data_o(fifo_rdata),
		.pop_i(fifo_pop)
	);
	// Trace: design.sv:16626:3
	assign fetch_rdata_o = (fifo_empty ? resp_rdata : fifo_rdata);
	// Trace: design.sv:16632:3
	cv32e40p_obi_interface #(.TRANS_STABLE(0)) instruction_obi_i(
		.clk(clk),
		.rst_n(rst_n),
		.trans_valid_i(trans_valid),
		.trans_ready_o(trans_ready),
		.trans_addr_i({trans_addr[31:2], 2'b00}),
		.trans_we_i(1'b0),
		.trans_be_i(4'b1111),
		.trans_wdata_i(32'b00000000000000000000000000000000),
		.trans_atop_i(6'b000000),
		.resp_valid_o(resp_valid),
		.resp_rdata_o(resp_rdata),
		.resp_err_o(resp_err),
		.obi_req_o(instr_req_o),
		.obi_gnt_i(instr_gnt_i),
		.obi_addr_o(instr_addr_o),
		.obi_we_o(),
		.obi_be_o(),
		.obi_wdata_o(),
		.obi_atop_o(),
		.obi_rdata_i(instr_rdata_i),
		.obi_rvalid_i(instr_rvalid_i),
		.obi_err_i(instr_err_i)
	);
endmodule
module cv32e40p_prefetch_controller (
	clk,
	rst_n,
	req_i,
	branch_i,
	branch_addr_i,
	busy_o,
	hwlp_jump_i,
	hwlp_target_i,
	trans_valid_o,
	trans_ready_i,
	trans_addr_o,
	resp_valid_i,
	fetch_ready_i,
	fetch_valid_o,
	fifo_push_o,
	fifo_pop_o,
	fifo_flush_o,
	fifo_flush_but_first_o,
	fifo_cnt_i,
	fifo_empty_i
);
	reg _sv2v_0;
	// Trace: design.sv:16777:15
	parameter PULP_OBI = 0;
	// Trace: design.sv:16778:15
	parameter PULP_XPULP = 1;
	// Trace: design.sv:16779:15
	parameter DEPTH = 4;
	// Trace: design.sv:16780:15
	parameter FIFO_ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:16782:5
	input wire clk;
	// Trace: design.sv:16783:5
	input wire rst_n;
	// Trace: design.sv:16786:5
	input wire req_i;
	// Trace: design.sv:16787:5
	input wire branch_i;
	// Trace: design.sv:16788:5
	input wire [31:0] branch_addr_i;
	// Trace: design.sv:16789:5
	output wire busy_o;
	// Trace: design.sv:16792:5
	input wire hwlp_jump_i;
	// Trace: design.sv:16793:5
	input wire [31:0] hwlp_target_i;
	// Trace: design.sv:16796:5
	output wire trans_valid_o;
	// Trace: design.sv:16797:5
	input wire trans_ready_i;
	// Trace: design.sv:16798:5
	output reg [31:0] trans_addr_o;
	// Trace: design.sv:16801:5
	input wire resp_valid_i;
	// Trace: design.sv:16804:5
	input wire fetch_ready_i;
	// Trace: design.sv:16805:5
	output wire fetch_valid_o;
	// Trace: design.sv:16808:5
	output wire fifo_push_o;
	// Trace: design.sv:16809:5
	output wire fifo_pop_o;
	// Trace: design.sv:16810:5
	output wire fifo_flush_o;
	// Trace: design.sv:16811:5
	output wire fifo_flush_but_first_o;
	// Trace: design.sv:16812:5
	input wire [FIFO_ADDR_DEPTH:0] fifo_cnt_i;
	// Trace: design.sv:16813:5
	input wire fifo_empty_i;
	// Trace: design.sv:16816:3
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:16818:3
	// removed localparam type cv32e40p_pkg_prefetch_state_e
	reg state_q;
	reg next_state;
	// Trace: design.sv:16820:3
	reg [FIFO_ADDR_DEPTH:0] cnt_q;
	// Trace: design.sv:16821:3
	reg [FIFO_ADDR_DEPTH:0] next_cnt;
	// Trace: design.sv:16822:3
	wire count_up;
	// Trace: design.sv:16823:3
	wire count_down;
	// Trace: design.sv:16825:3
	reg [FIFO_ADDR_DEPTH:0] flush_cnt_q;
	// Trace: design.sv:16826:3
	reg [FIFO_ADDR_DEPTH:0] next_flush_cnt;
	// Trace: design.sv:16829:3
	reg [31:0] trans_addr_q;
	wire [31:0] trans_addr_incr;
	// Trace: design.sv:16832:3
	wire [31:0] aligned_branch_addr;
	// Trace: design.sv:16835:3
	wire fifo_valid;
	// Trace: design.sv:16836:3
	wire [FIFO_ADDR_DEPTH:0] fifo_cnt_masked;
	// Trace: design.sv:16839:3
	wire hwlp_wait_resp_flush;
	// Trace: design.sv:16840:3
	reg hwlp_flush_after_resp;
	// Trace: design.sv:16841:3
	reg [FIFO_ADDR_DEPTH:0] hwlp_flush_cnt_delayed_q;
	// Trace: design.sv:16842:3
	wire hwlp_flush_resp_delayed;
	// Trace: design.sv:16843:3
	wire hwlp_flush_resp;
	// Trace: design.sv:16850:3
	assign busy_o = (cnt_q != 3'b000) || trans_valid_o;
	// Trace: design.sv:16859:3
	assign fetch_valid_o = (fifo_valid || resp_valid_i) && !(branch_i || (flush_cnt_q > 0));
	// Trace: design.sv:16871:3
	assign aligned_branch_addr = {branch_addr_i[31:2], 2'b00};
	// Trace: design.sv:16874:3
	assign trans_addr_incr = {trans_addr_q[31:2], 2'b00} + 32'd4;
	// Trace: design.sv:16877:3
	generate
		if (PULP_OBI == 0) begin : gen_no_pulp_obi
			// Trace: design.sv:16882:7
			assign trans_valid_o = req_i && ((fifo_cnt_masked + cnt_q) < DEPTH);
		end
		else begin : gen_pulp_obi
			// Trace: design.sv:16886:7
			assign trans_valid_o = (cnt_q == 3'b000 ? req_i && ((fifo_cnt_masked + cnt_q) < DEPTH) : (req_i && ((fifo_cnt_masked + cnt_q) < DEPTH)) && resp_valid_i);
		end
	endgenerate
	// Trace: design.sv:16897:3
	assign fifo_cnt_masked = (branch_i || hwlp_jump_i ? {(FIFO_ADDR_DEPTH >= 0 ? FIFO_ADDR_DEPTH + 1 : 1 - FIFO_ADDR_DEPTH) {1'sb0}} : fifo_cnt_i);
	// Trace: design.sv:16900:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:16901:5
		next_state = state_q;
		// Trace: design.sv:16902:5
		trans_addr_o = trans_addr_q;
		// Trace: design.sv:16904:5
		case (state_q)
			1'd0: begin
				// Trace: design.sv:16907:9
				// Trace: design.sv:16908:11
				if (branch_i)
					// Trace: design.sv:16911:13
					trans_addr_o = aligned_branch_addr;
				else if (hwlp_jump_i)
					// Trace: design.sv:16913:13
					trans_addr_o = hwlp_target_i;
				else
					// Trace: design.sv:16915:13
					trans_addr_o = trans_addr_incr;
				if ((branch_i || hwlp_jump_i) && !(trans_valid_o && trans_ready_i))
					// Trace: design.sv:16920:11
					next_state = 1'd1;
			end
			1'd1: begin
				// Trace: design.sv:16928:9
				trans_addr_o = (branch_i ? aligned_branch_addr : trans_addr_q);
				// Trace: design.sv:16929:9
				if (trans_valid_o && trans_ready_i)
					// Trace: design.sv:16931:11
					next_state = 1'd0;
			end
		endcase
	end
	// Trace: design.sv:16946:3
	assign fifo_valid = !fifo_empty_i;
	// Trace: design.sv:16947:3
	assign fifo_push_o = (resp_valid_i && (fifo_valid || !fetch_ready_i)) && !(branch_i || (flush_cnt_q > 0));
	// Trace: design.sv:16948:3
	assign fifo_pop_o = fifo_valid && fetch_ready_i;
	// Trace: design.sv:16959:3
	assign count_up = trans_valid_o && trans_ready_i;
	// Trace: design.sv:16960:3
	assign count_down = resp_valid_i;
	// Trace: design.sv:16962:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:16963:5
		case ({count_up, count_down})
			2'b00:
				// Trace: design.sv:16967:9
				next_cnt = cnt_q;
			2'b01:
				// Trace: design.sv:16970:9
				next_cnt = cnt_q - 1'b1;
			2'b10:
				// Trace: design.sv:16973:9
				next_cnt = cnt_q + 1'b1;
			2'b11:
				// Trace: design.sv:16976:9
				next_cnt = cnt_q;
		endcase
	end
	// Trace: design.sv:16981:3
	generate
		if (PULP_XPULP) begin : gen_hwlp
			// Trace: design.sv:16988:7
			assign fifo_flush_o = branch_i || ((hwlp_jump_i && !fifo_empty_i) && fifo_pop_o);
			// Trace: design.sv:16989:7
			assign fifo_flush_but_first_o = (hwlp_jump_i && !fifo_empty_i) && !fifo_pop_o;
			// Trace: design.sv:16997:7
			assign hwlp_flush_resp = hwlp_jump_i && !(fifo_empty_i && !resp_valid_i);
			// Trace: design.sv:17006:7
			assign hwlp_wait_resp_flush = hwlp_jump_i && (fifo_empty_i && !resp_valid_i);
			// Trace: design.sv:17008:7
			always @(posedge clk or negedge rst_n)
				// Trace: design.sv:17009:9
				if (~rst_n) begin
					// Trace: design.sv:17010:11
					hwlp_flush_after_resp <= 1'b0;
					// Trace: design.sv:17011:11
					hwlp_flush_cnt_delayed_q <= 2'b00;
				end
				else
					// Trace: design.sv:17013:11
					if (branch_i) begin
						// Trace: design.sv:17015:13
						hwlp_flush_after_resp <= 1'b0;
						// Trace: design.sv:17016:13
						hwlp_flush_cnt_delayed_q <= 2'b00;
					end
					else
						// Trace: design.sv:17018:13
						if (hwlp_wait_resp_flush) begin
							// Trace: design.sv:17019:15
							hwlp_flush_after_resp <= 1'b1;
							// Trace: design.sv:17021:15
							hwlp_flush_cnt_delayed_q <= cnt_q - 1'b1;
						end
						else
							// Trace: design.sv:17024:15
							if (hwlp_flush_resp_delayed) begin
								// Trace: design.sv:17025:17
								hwlp_flush_after_resp <= 1'b0;
								// Trace: design.sv:17026:17
								hwlp_flush_cnt_delayed_q <= 2'b00;
							end
			// Trace: design.sv:17036:7
			assign hwlp_flush_resp_delayed = hwlp_flush_after_resp && resp_valid_i;
		end
		else begin : gen_no_hwlp
			// Trace: design.sv:17041:7
			assign fifo_flush_o = branch_i;
			// Trace: design.sv:17042:7
			assign fifo_flush_but_first_o = 1'b0;
			// Trace: design.sv:17043:7
			assign hwlp_flush_resp = 1'b0;
			// Trace: design.sv:17044:7
			assign hwlp_wait_resp_flush = 1'b0;
			// Trace: design.sv:17046:7
			wire [1:1] sv2v_tmp_9BC28;
			assign sv2v_tmp_9BC28 = 1'b0;
			always @(*) hwlp_flush_after_resp = sv2v_tmp_9BC28;
			// Trace: design.sv:17047:7
			wire [(FIFO_ADDR_DEPTH >= 0 ? FIFO_ADDR_DEPTH + 1 : 1 - FIFO_ADDR_DEPTH):1] sv2v_tmp_2B514;
			assign sv2v_tmp_2B514 = 2'b00;
			always @(*) hwlp_flush_cnt_delayed_q = sv2v_tmp_2B514;
			// Trace: design.sv:17048:7
			assign hwlp_flush_resp_delayed = 1'b0;
		end
	endgenerate
	// Trace: design.sv:17058:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:17059:5
		next_flush_cnt = flush_cnt_q;
		// Trace: design.sv:17064:5
		if (branch_i || hwlp_flush_resp) begin
			// Trace: design.sv:17065:7
			next_flush_cnt = cnt_q;
			// Trace: design.sv:17066:7
			if (resp_valid_i && (cnt_q > 0))
				// Trace: design.sv:17067:9
				next_flush_cnt = cnt_q - 1'b1;
		end
		else if (hwlp_flush_resp_delayed)
			// Trace: design.sv:17073:7
			next_flush_cnt = hwlp_flush_cnt_delayed_q;
		else if (resp_valid_i && (flush_cnt_q > 0))
			// Trace: design.sv:17075:7
			next_flush_cnt = flush_cnt_q - 1'b1;
	end
	// Trace: design.sv:17083:3
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:17084:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:17085:7
			state_q <= 1'd0;
			// Trace: design.sv:17086:7
			cnt_q <= 1'sb0;
			// Trace: design.sv:17087:7
			flush_cnt_q <= 1'sb0;
			// Trace: design.sv:17088:7
			trans_addr_q <= 1'sb0;
		end
		else begin
			// Trace: design.sv:17090:7
			state_q <= next_state;
			// Trace: design.sv:17091:7
			cnt_q <= next_cnt;
			// Trace: design.sv:17092:7
			flush_cnt_q <= next_flush_cnt;
			// Trace: design.sv:17093:7
			if ((branch_i || hwlp_jump_i) || (trans_valid_o && trans_ready_i))
				// Trace: design.sv:17094:9
				trans_addr_q <= trans_addr_o;
		end
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_obi_interface (
	clk,
	rst_n,
	trans_valid_i,
	trans_ready_o,
	trans_addr_i,
	trans_we_i,
	trans_be_i,
	trans_wdata_i,
	trans_atop_i,
	resp_valid_o,
	resp_rdata_o,
	resp_err_o,
	obi_req_o,
	obi_gnt_i,
	obi_addr_o,
	obi_we_o,
	obi_be_o,
	obi_wdata_o,
	obi_atop_o,
	obi_rdata_i,
	obi_rvalid_i,
	obi_err_i
);
	reg _sv2v_0;
	// Trace: design.sv:17138:15
	parameter TRANS_STABLE = 0;
	// Trace: design.sv:17140:5
	input wire clk;
	// Trace: design.sv:17141:5
	input wire rst_n;
	// Trace: design.sv:17144:5
	input wire trans_valid_i;
	// Trace: design.sv:17145:5
	output wire trans_ready_o;
	// Trace: design.sv:17146:5
	input wire [31:0] trans_addr_i;
	// Trace: design.sv:17147:5
	input wire trans_we_i;
	// Trace: design.sv:17148:5
	input wire [3:0] trans_be_i;
	// Trace: design.sv:17149:5
	input wire [31:0] trans_wdata_i;
	// Trace: design.sv:17150:5
	input wire [5:0] trans_atop_i;
	// Trace: design.sv:17153:5
	output wire resp_valid_o;
	// Trace: design.sv:17154:5
	output wire [31:0] resp_rdata_o;
	// Trace: design.sv:17155:5
	output wire resp_err_o;
	// Trace: design.sv:17158:5
	output reg obi_req_o;
	// Trace: design.sv:17159:5
	input wire obi_gnt_i;
	// Trace: design.sv:17160:5
	output reg [31:0] obi_addr_o;
	// Trace: design.sv:17161:5
	output reg obi_we_o;
	// Trace: design.sv:17162:5
	output reg [3:0] obi_be_o;
	// Trace: design.sv:17163:5
	output reg [31:0] obi_wdata_o;
	// Trace: design.sv:17164:5
	output reg [5:0] obi_atop_o;
	// Trace: design.sv:17165:5
	input wire [31:0] obi_rdata_i;
	// Trace: design.sv:17166:5
	input wire obi_rvalid_i;
	// Trace: design.sv:17167:5
	input wire obi_err_i;
	// Trace: design.sv:17170:3
	reg state_q;
	reg next_state;
	// Trace: design.sv:17184:3
	assign resp_valid_o = obi_rvalid_i;
	// Trace: design.sv:17185:3
	assign resp_rdata_o = obi_rdata_i;
	// Trace: design.sv:17186:3
	assign resp_err_o = obi_err_i;
	// Trace: design.sv:17193:3
	generate
		if (TRANS_STABLE) begin : gen_trans_stable
			// Trace: design.sv:17198:7
			wire [1:1] sv2v_tmp_E8019;
			assign sv2v_tmp_E8019 = trans_valid_i;
			always @(*) obi_req_o = sv2v_tmp_E8019;
			// Trace: design.sv:17199:7
			wire [32:1] sv2v_tmp_2DFD9;
			assign sv2v_tmp_2DFD9 = trans_addr_i;
			always @(*) obi_addr_o = sv2v_tmp_2DFD9;
			// Trace: design.sv:17200:7
			wire [1:1] sv2v_tmp_367C5;
			assign sv2v_tmp_367C5 = trans_we_i;
			always @(*) obi_we_o = sv2v_tmp_367C5;
			// Trace: design.sv:17201:7
			wire [4:1] sv2v_tmp_738B5;
			assign sv2v_tmp_738B5 = trans_be_i;
			always @(*) obi_be_o = sv2v_tmp_738B5;
			// Trace: design.sv:17202:7
			wire [32:1] sv2v_tmp_F8E9B;
			assign sv2v_tmp_F8E9B = trans_wdata_i;
			always @(*) obi_wdata_o = sv2v_tmp_F8E9B;
			// Trace: design.sv:17203:7
			wire [6:1] sv2v_tmp_E7AA9;
			assign sv2v_tmp_E7AA9 = trans_atop_i;
			always @(*) obi_atop_o = sv2v_tmp_E7AA9;
			// Trace: design.sv:17205:7
			assign trans_ready_o = obi_gnt_i;
			// Trace: design.sv:17208:7
			wire [1:1] sv2v_tmp_7058D;
			assign sv2v_tmp_7058D = 1'd0;
			always @(*) state_q = sv2v_tmp_7058D;
			// Trace: design.sv:17209:7
			wire [1:1] sv2v_tmp_B3134;
			assign sv2v_tmp_B3134 = 1'd0;
			always @(*) next_state = sv2v_tmp_B3134;
		end
		else begin : gen_no_trans_stable
			// Trace: design.sv:17213:7
			reg [31:0] obi_addr_q;
			// Trace: design.sv:17214:7
			reg obi_we_q;
			// Trace: design.sv:17215:7
			reg [3:0] obi_be_q;
			// Trace: design.sv:17216:7
			reg [31:0] obi_wdata_q;
			// Trace: design.sv:17217:7
			reg [5:0] obi_atop_q;
			// Trace: design.sv:17228:7
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:17229:9
				next_state = state_q;
				// Trace: design.sv:17231:9
				case (state_q)
					1'd0:
						// Trace: design.sv:17235:13
						if (obi_req_o && !obi_gnt_i)
							// Trace: design.sv:17238:15
							next_state = 1'd1;
					1'd1:
						// Trace: design.sv:17244:13
						if (obi_gnt_i)
							// Trace: design.sv:17246:15
							next_state = 1'd0;
				endcase
			end
			// Trace: design.sv:17253:7
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:17254:9
				if (state_q == 1'd0) begin
					// Trace: design.sv:17255:11
					obi_req_o = trans_valid_i;
					// Trace: design.sv:17256:11
					obi_addr_o = trans_addr_i;
					// Trace: design.sv:17257:11
					obi_we_o = trans_we_i;
					// Trace: design.sv:17258:11
					obi_be_o = trans_be_i;
					// Trace: design.sv:17259:11
					obi_wdata_o = trans_wdata_i;
					// Trace: design.sv:17260:11
					obi_atop_o = trans_atop_i;
				end
				else begin
					// Trace: design.sv:17263:11
					obi_req_o = 1'b1;
					// Trace: design.sv:17264:11
					obi_addr_o = obi_addr_q;
					// Trace: design.sv:17265:11
					obi_we_o = obi_we_q;
					// Trace: design.sv:17266:11
					obi_be_o = obi_be_q;
					// Trace: design.sv:17267:11
					obi_wdata_o = obi_wdata_q;
					// Trace: design.sv:17268:11
					obi_atop_o = obi_atop_q;
				end
			end
			// Trace: design.sv:17276:7
			always @(posedge clk or negedge rst_n)
				// Trace: design.sv:17277:9
				if (rst_n == 1'b0) begin
					// Trace: design.sv:17278:11
					state_q <= 1'd0;
					// Trace: design.sv:17279:11
					obi_addr_q <= 32'b00000000000000000000000000000000;
					// Trace: design.sv:17280:11
					obi_we_q <= 1'b0;
					// Trace: design.sv:17281:11
					obi_be_q <= 4'b0000;
					// Trace: design.sv:17282:11
					obi_wdata_q <= 32'b00000000000000000000000000000000;
					// Trace: design.sv:17283:11
					obi_atop_q <= 6'b000000;
				end
				else begin
					// Trace: design.sv:17285:11
					state_q <= next_state;
					// Trace: design.sv:17286:11
					if ((state_q == 1'd0) && (next_state == 1'd1)) begin
						// Trace: design.sv:17288:13
						obi_addr_q <= obi_addr_o;
						// Trace: design.sv:17289:13
						obi_we_q <= obi_we_o;
						// Trace: design.sv:17290:13
						obi_be_q <= obi_be_o;
						// Trace: design.sv:17291:13
						obi_wdata_q <= obi_wdata_o;
						// Trace: design.sv:17292:13
						obi_atop_q <= obi_atop_o;
					end
				end
			// Trace: design.sv:17300:7
			assign trans_ready_o = state_q == 1'd0;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_aligner (
	clk,
	rst_n,
	fetch_valid_i,
	aligner_ready_o,
	if_valid_i,
	fetch_rdata_i,
	instr_aligned_o,
	instr_valid_o,
	branch_addr_i,
	branch_i,
	hwlp_addr_i,
	hwlp_update_pc_i,
	pc_o
);
	reg _sv2v_0;
	// Trace: design.sv:17329:5
	input wire clk;
	// Trace: design.sv:17330:5
	input wire rst_n;
	// Trace: design.sv:17332:5
	input wire fetch_valid_i;
	// Trace: design.sv:17333:5
	output reg aligner_ready_o;
	// Trace: design.sv:17335:5
	input wire if_valid_i;
	// Trace: design.sv:17337:5
	input wire [31:0] fetch_rdata_i;
	// Trace: design.sv:17338:5
	output reg [31:0] instr_aligned_o;
	// Trace: design.sv:17339:5
	output reg instr_valid_o;
	// Trace: design.sv:17341:5
	input wire [31:0] branch_addr_i;
	// Trace: design.sv:17342:5
	input wire branch_i;
	// Trace: design.sv:17344:5
	input wire [31:0] hwlp_addr_i;
	// Trace: design.sv:17345:5
	input wire hwlp_update_pc_i;
	// Trace: design.sv:17347:5
	output wire [31:0] pc_o;
	// Trace: design.sv:17350:3
	reg [2:0] state;
	reg [2:0] next_state;
	// Trace: design.sv:17359:3
	reg [15:0] r_instr_h;
	// Trace: design.sv:17360:3
	reg [31:0] hwlp_addr_q;
	// Trace: design.sv:17361:3
	reg [31:0] pc_q;
	reg [31:0] pc_n;
	// Trace: design.sv:17362:3
	reg update_state;
	// Trace: design.sv:17363:3
	wire [31:0] pc_plus4;
	wire [31:0] pc_plus2;
	// Trace: design.sv:17364:3
	reg aligner_ready_q;
	reg hwlp_update_pc_q;
	// Trace: design.sv:17366:3
	assign pc_o = pc_q;
	// Trace: design.sv:17368:3
	assign pc_plus2 = pc_q + 2;
	// Trace: design.sv:17369:3
	assign pc_plus4 = pc_q + 4;
	// Trace: design.sv:17371:3
	always @(posedge clk or negedge rst_n) begin : proc_SEQ_FSM
		// Trace: design.sv:17372:5
		if (~rst_n) begin
			// Trace: design.sv:17373:7
			state <= 3'd0;
			// Trace: design.sv:17374:7
			r_instr_h <= 1'sb0;
			// Trace: design.sv:17375:7
			hwlp_addr_q <= 1'sb0;
			// Trace: design.sv:17376:7
			pc_q <= 1'sb0;
			// Trace: design.sv:17377:7
			aligner_ready_q <= 1'b0;
			// Trace: design.sv:17378:7
			hwlp_update_pc_q <= 1'b0;
		end
		else
			// Trace: design.sv:17380:7
			if (update_state) begin
				// Trace: design.sv:17381:9
				pc_q <= pc_n;
				// Trace: design.sv:17382:9
				state <= next_state;
				// Trace: design.sv:17383:9
				r_instr_h <= fetch_rdata_i[31:16];
				// Trace: design.sv:17384:9
				aligner_ready_q <= aligner_ready_o;
				// Trace: design.sv:17385:9
				hwlp_update_pc_q <= 1'b0;
			end
			else
				// Trace: design.sv:17387:9
				if (hwlp_update_pc_i) begin
					// Trace: design.sv:17388:11
					hwlp_addr_q <= hwlp_addr_i;
					// Trace: design.sv:17389:11
					hwlp_update_pc_q <= 1'b1;
				end
	end
	// Trace: design.sv:17396:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:17399:5
		pc_n = pc_q;
		// Trace: design.sv:17400:5
		instr_valid_o = fetch_valid_i;
		// Trace: design.sv:17401:5
		instr_aligned_o = fetch_rdata_i;
		// Trace: design.sv:17402:5
		aligner_ready_o = 1'b1;
		// Trace: design.sv:17403:5
		update_state = 1'b0;
		// Trace: design.sv:17404:5
		next_state = state;
		// Trace: design.sv:17407:5
		case (state)
			3'd0:
				// Trace: design.sv:17409:9
				if (fetch_rdata_i[1:0] == 2'b11) begin
					// Trace: design.sv:17414:11
					next_state = 3'd0;
					// Trace: design.sv:17415:11
					pc_n = pc_plus4;
					// Trace: design.sv:17416:11
					instr_aligned_o = fetch_rdata_i;
					// Trace: design.sv:17418:11
					update_state = fetch_valid_i & if_valid_i;
					// Trace: design.sv:17419:11
					if (hwlp_update_pc_i || hwlp_update_pc_q)
						// Trace: design.sv:17420:13
						pc_n = (hwlp_update_pc_i ? hwlp_addr_i : hwlp_addr_q);
				end
				else begin
					// Trace: design.sv:17426:11
					next_state = 3'd1;
					// Trace: design.sv:17427:11
					pc_n = pc_plus2;
					// Trace: design.sv:17428:11
					instr_aligned_o = fetch_rdata_i;
					// Trace: design.sv:17430:11
					update_state = fetch_valid_i & if_valid_i;
				end
			3'd1:
				// Trace: design.sv:17436:9
				if (r_instr_h[1:0] == 2'b11) begin
					// Trace: design.sv:17442:11
					next_state = 3'd1;
					// Trace: design.sv:17443:11
					pc_n = pc_plus4;
					// Trace: design.sv:17444:11
					instr_aligned_o = {fetch_rdata_i[15:0], r_instr_h[15:0]};
					// Trace: design.sv:17446:11
					update_state = fetch_valid_i & if_valid_i;
				end
				else begin
					// Trace: design.sv:17453:11
					instr_aligned_o = {fetch_rdata_i[31:16], r_instr_h[15:0]};
					// Trace: design.sv:17454:11
					next_state = 3'd2;
					// Trace: design.sv:17455:11
					instr_valid_o = 1'b1;
					// Trace: design.sv:17456:11
					pc_n = pc_plus2;
					// Trace: design.sv:17459:11
					aligner_ready_o = !fetch_valid_i;
					// Trace: design.sv:17461:11
					update_state = if_valid_i;
				end
			3'd2: begin
				// Trace: design.sv:17468:9
				instr_valid_o = !aligner_ready_q || fetch_valid_i;
				// Trace: design.sv:17469:9
				if (fetch_rdata_i[1:0] == 2'b11) begin
					// Trace: design.sv:17475:11
					next_state = 3'd0;
					// Trace: design.sv:17476:11
					pc_n = pc_plus4;
					// Trace: design.sv:17477:11
					instr_aligned_o = fetch_rdata_i;
					// Trace: design.sv:17479:11
					update_state = (!aligner_ready_q | fetch_valid_i) & if_valid_i;
				end
				else begin
					// Trace: design.sv:17486:11
					next_state = 3'd1;
					// Trace: design.sv:17487:11
					pc_n = pc_plus2;
					// Trace: design.sv:17488:11
					instr_aligned_o = fetch_rdata_i;
					// Trace: design.sv:17490:11
					update_state = (!aligner_ready_q | fetch_valid_i) & if_valid_i;
				end
			end
			3'd3:
				// Trace: design.sv:17497:9
				if (fetch_rdata_i[17:16] == 2'b11) begin
					// Trace: design.sv:17501:11
					next_state = 3'd1;
					// Trace: design.sv:17502:11
					instr_valid_o = 1'b0;
					// Trace: design.sv:17503:11
					pc_n = pc_q;
					// Trace: design.sv:17504:11
					instr_aligned_o = fetch_rdata_i;
					// Trace: design.sv:17506:11
					update_state = fetch_valid_i & if_valid_i;
				end
				else begin
					// Trace: design.sv:17511:11
					next_state = 3'd0;
					// Trace: design.sv:17512:11
					pc_n = pc_plus2;
					// Trace: design.sv:17513:11
					instr_aligned_o = {fetch_rdata_i[31:16], fetch_rdata_i[31:16]};
					// Trace: design.sv:17517:11
					update_state = fetch_valid_i & if_valid_i;
				end
		endcase
		if (branch_i) begin
			// Trace: design.sv:17526:7
			update_state = 1'b1;
			// Trace: design.sv:17527:7
			pc_n = branch_addr_i;
			// Trace: design.sv:17528:7
			next_state = (branch_addr_i[1] ? 3'd3 : 3'd0);
		end
	end
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_sleep_unit (
	clk_ungated_i,
	rst_n,
	clk_gated_o,
	scan_cg_en_i,
	core_sleep_o,
	fetch_enable_i,
	fetch_enable_o,
	if_busy_i,
	ctrl_busy_i,
	lsu_busy_i,
	apu_busy_i,
	pulp_clock_en_i,
	p_elw_start_i,
	p_elw_finish_i,
	debug_p_elw_no_sleep_i,
	wake_from_sleep_i
);
	// Trace: design.sv:17614:15
	parameter PULP_CLUSTER = 0;
	// Trace: design.sv:17617:5
	input wire clk_ungated_i;
	// Trace: design.sv:17618:5
	input wire rst_n;
	// Trace: design.sv:17619:5
	output wire clk_gated_o;
	// Trace: design.sv:17620:5
	input wire scan_cg_en_i;
	// Trace: design.sv:17623:5
	output wire core_sleep_o;
	// Trace: design.sv:17626:5
	input wire fetch_enable_i;
	// Trace: design.sv:17627:5
	output wire fetch_enable_o;
	// Trace: design.sv:17630:5
	input wire if_busy_i;
	// Trace: design.sv:17631:5
	input wire ctrl_busy_i;
	// Trace: design.sv:17632:5
	input wire lsu_busy_i;
	// Trace: design.sv:17633:5
	input wire apu_busy_i;
	// Trace: design.sv:17636:5
	input wire pulp_clock_en_i;
	// Trace: design.sv:17637:5
	input wire p_elw_start_i;
	// Trace: design.sv:17638:5
	input wire p_elw_finish_i;
	// Trace: design.sv:17639:5
	input wire debug_p_elw_no_sleep_i;
	// Trace: design.sv:17642:5
	input wire wake_from_sleep_i;
	// Trace: design.sv:17645:3
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:17647:3
	reg fetch_enable_q;
	// Trace: design.sv:17648:3
	wire fetch_enable_d;
	// Trace: design.sv:17649:3
	reg core_busy_q;
	// Trace: design.sv:17650:3
	wire core_busy_d;
	// Trace: design.sv:17651:3
	reg p_elw_busy_q;
	// Trace: design.sv:17652:3
	wire p_elw_busy_d;
	// Trace: design.sv:17653:3
	wire clock_en;
	// Trace: design.sv:17660:3
	assign fetch_enable_d = (fetch_enable_i ? 1'b1 : fetch_enable_q);
	// Trace: design.sv:17662:3
	generate
		if (PULP_CLUSTER) begin : g_pulp_sleep
			// Trace: design.sv:17666:7
			assign core_busy_d = (p_elw_busy_d ? if_busy_i || apu_busy_i : 1'b1);
			// Trace: design.sv:17669:7
			assign clock_en = fetch_enable_q && (pulp_clock_en_i || core_busy_q);
			// Trace: design.sv:17672:7
			assign core_sleep_o = (p_elw_busy_d && !core_busy_q) && !debug_p_elw_no_sleep_i;
			// Trace: design.sv:17675:7
			assign p_elw_busy_d = (p_elw_start_i ? 1'b1 : (p_elw_finish_i ? 1'b0 : p_elw_busy_q));
		end
		else begin : g_no_pulp_sleep
			// Trace: design.sv:17680:7
			assign core_busy_d = ((if_busy_i || ctrl_busy_i) || lsu_busy_i) || apu_busy_i;
			// Trace: design.sv:17683:7
			assign clock_en = fetch_enable_q && (wake_from_sleep_i || core_busy_q);
			// Trace: design.sv:17687:7
			assign core_sleep_o = fetch_enable_q && !clock_en;
			// Trace: design.sv:17690:7
			assign p_elw_busy_d = 1'b0;
		end
	endgenerate
	// Trace: design.sv:17695:3
	always @(posedge clk_ungated_i or negedge rst_n)
		// Trace: design.sv:17696:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:17697:7
			core_busy_q <= 1'b0;
			// Trace: design.sv:17698:7
			p_elw_busy_q <= 1'b0;
			// Trace: design.sv:17699:7
			fetch_enable_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:17701:7
			core_busy_q <= core_busy_d;
			// Trace: design.sv:17702:7
			p_elw_busy_q <= p_elw_busy_d;
			// Trace: design.sv:17703:7
			fetch_enable_q <= fetch_enable_d;
		end
	// Trace: design.sv:17708:3
	assign fetch_enable_o = fetch_enable_q;
	// Trace: design.sv:17711:3
	cv32e40p_clock_gate core_clock_gate_i(
		.clk_i(clk_ungated_i),
		.en_i(clock_en),
		.scan_cg_en_i(scan_cg_en_i),
		.clk_o(clk_gated_o)
	);
endmodule
module cv32e40p_core (
	clk_i,
	rst_ni,
	pulp_clock_en_i,
	scan_cg_en_i,
	boot_addr_i,
	mtvec_addr_i,
	dm_halt_addr_i,
	hart_id_i,
	dm_exception_addr_i,
	instr_req_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_addr_o,
	instr_rdata_i,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_we_o,
	data_be_o,
	data_addr_o,
	data_wdata_o,
	data_rdata_i,
	apu_req_o,
	apu_gnt_i,
	apu_operands_o,
	apu_op_o,
	apu_flags_o,
	apu_rvalid_i,
	apu_result_i,
	apu_flags_i,
	irq_i,
	irq_ack_o,
	irq_id_o,
	debug_req_i,
	debug_havereset_o,
	debug_running_o,
	debug_halted_o,
	fetch_enable_i,
	core_sleep_o
);
	// removed import cv32e40p_apu_core_pkg::*;
	// Trace: design.sv:17883:15
	parameter PULP_XPULP = 0;
	// Trace: design.sv:17884:15
	parameter PULP_CLUSTER = 0;
	// Trace: design.sv:17885:15
	parameter FPU = 0;
	// Trace: design.sv:17886:15
	parameter PULP_ZFINX = 0;
	// Trace: design.sv:17887:15
	parameter NUM_MHPMCOUNTERS = 1;
	// Trace: design.sv:17890:5
	input wire clk_i;
	// Trace: design.sv:17891:5
	input wire rst_ni;
	// Trace: design.sv:17893:5
	input wire pulp_clock_en_i;
	// Trace: design.sv:17894:5
	input wire scan_cg_en_i;
	// Trace: design.sv:17897:5
	input wire [31:0] boot_addr_i;
	// Trace: design.sv:17898:5
	input wire [31:0] mtvec_addr_i;
	// Trace: design.sv:17899:5
	input wire [31:0] dm_halt_addr_i;
	// Trace: design.sv:17900:5
	input wire [31:0] hart_id_i;
	// Trace: design.sv:17901:5
	input wire [31:0] dm_exception_addr_i;
	// Trace: design.sv:17904:5
	output wire instr_req_o;
	// Trace: design.sv:17905:5
	input wire instr_gnt_i;
	// Trace: design.sv:17906:5
	input wire instr_rvalid_i;
	// Trace: design.sv:17907:5
	output wire [31:0] instr_addr_o;
	// Trace: design.sv:17908:5
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:17911:5
	output wire data_req_o;
	// Trace: design.sv:17912:5
	input wire data_gnt_i;
	// Trace: design.sv:17913:5
	input wire data_rvalid_i;
	// Trace: design.sv:17914:5
	output wire data_we_o;
	// Trace: design.sv:17915:5
	output wire [3:0] data_be_o;
	// Trace: design.sv:17916:5
	output wire [31:0] data_addr_o;
	// Trace: design.sv:17917:5
	output wire [31:0] data_wdata_o;
	// Trace: design.sv:17918:5
	input wire [31:0] data_rdata_i;
	// Trace: design.sv:17922:5
	output wire apu_req_o;
	// Trace: design.sv:17923:5
	input wire apu_gnt_i;
	// Trace: design.sv:17925:5
	localparam cv32e40p_apu_core_pkg_APU_NARGS_CPU = 3;
	output wire [95:0] apu_operands_o;
	// Trace: design.sv:17926:5
	localparam cv32e40p_apu_core_pkg_APU_WOP_CPU = 6;
	output wire [5:0] apu_op_o;
	// Trace: design.sv:17927:5
	localparam cv32e40p_apu_core_pkg_APU_NDSFLAGS_CPU = 15;
	output wire [14:0] apu_flags_o;
	// Trace: design.sv:17929:5
	input wire apu_rvalid_i;
	// Trace: design.sv:17930:5
	input wire [31:0] apu_result_i;
	// Trace: design.sv:17931:5
	localparam cv32e40p_apu_core_pkg_APU_NUSFLAGS_CPU = 5;
	input wire [4:0] apu_flags_i;
	// Trace: design.sv:17934:5
	input wire [31:0] irq_i;
	// Trace: design.sv:17935:5
	output wire irq_ack_o;
	// Trace: design.sv:17936:5
	output wire [4:0] irq_id_o;
	// Trace: design.sv:17939:5
	input wire debug_req_i;
	// Trace: design.sv:17940:5
	output wire debug_havereset_o;
	// Trace: design.sv:17941:5
	output wire debug_running_o;
	// Trace: design.sv:17942:5
	output wire debug_halted_o;
	// Trace: design.sv:17945:5
	input wire fetch_enable_i;
	// Trace: design.sv:17946:5
	output wire core_sleep_o;
	// Trace: design.sv:17949:3
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:17952:3
	localparam PULP_SECURE = 0;
	// Trace: design.sv:17953:3
	localparam N_PMP_ENTRIES = 16;
	// Trace: design.sv:17954:3
	localparam USE_PMP = 0;
	// Trace: design.sv:17955:3
	localparam A_EXTENSION = 0;
	// Trace: design.sv:17956:3
	localparam DEBUG_TRIGGER_EN = 1;
	// Trace: design.sv:17962:3
	localparam PULP_OBI = 0;
	// Trace: design.sv:17968:3
	wire [5:0] data_atop_o;
	// Trace: design.sv:17969:3
	wire irq_sec_i;
	// Trace: design.sv:17970:3
	wire sec_lvl_o;
	// Trace: design.sv:17972:3
	localparam N_HWLP = 2;
	// Trace: design.sv:17973:3
	localparam N_HWLP_BITS = 1;
	// Trace: design.sv:17974:3
	localparam APU = (FPU == 1 ? 1 : 0);
	// Trace: design.sv:17978:3
	wire instr_valid_id;
	// Trace: design.sv:17979:3
	wire [31:0] instr_rdata_id;
	// Trace: design.sv:17980:3
	wire is_compressed_id;
	// Trace: design.sv:17981:3
	wire illegal_c_insn_id;
	// Trace: design.sv:17982:3
	wire is_fetch_failed_id;
	// Trace: design.sv:17984:3
	wire clear_instr_valid;
	// Trace: design.sv:17985:3
	wire pc_set;
	// Trace: design.sv:17987:3
	wire [3:0] pc_mux_id;
	// Trace: design.sv:17988:3
	wire [2:0] exc_pc_mux_id;
	// Trace: design.sv:17989:3
	wire [4:0] m_exc_vec_pc_mux_id;
	// Trace: design.sv:17990:3
	wire [4:0] u_exc_vec_pc_mux_id;
	// Trace: design.sv:17991:3
	wire [4:0] exc_cause;
	// Trace: design.sv:17993:3
	wire [1:0] trap_addr_mux;
	// Trace: design.sv:17995:3
	wire [31:0] pc_if;
	// Trace: design.sv:17996:3
	wire [31:0] pc_id;
	// Trace: design.sv:17999:3
	wire is_decoding;
	// Trace: design.sv:18001:3
	wire useincr_addr_ex;
	// Trace: design.sv:18002:3
	wire data_misaligned;
	// Trace: design.sv:18004:3
	wire mult_multicycle;
	// Trace: design.sv:18007:3
	wire [31:0] jump_target_id;
	wire [31:0] jump_target_ex;
	// Trace: design.sv:18008:3
	wire branch_in_ex;
	// Trace: design.sv:18009:3
	wire branch_decision;
	// Trace: design.sv:18011:3
	wire ctrl_busy;
	// Trace: design.sv:18012:3
	wire if_busy;
	// Trace: design.sv:18013:3
	wire lsu_busy;
	// Trace: design.sv:18014:3
	wire apu_busy;
	// Trace: design.sv:18016:3
	wire [31:0] pc_ex;
	// Trace: design.sv:18019:3
	wire alu_en_ex;
	// Trace: design.sv:18020:3
	localparam cv32e40p_pkg_ALU_OP_WIDTH = 7;
	// removed localparam type cv32e40p_pkg_alu_opcode_e
	wire [6:0] alu_operator_ex;
	// Trace: design.sv:18021:3
	wire [31:0] alu_operand_a_ex;
	// Trace: design.sv:18022:3
	wire [31:0] alu_operand_b_ex;
	// Trace: design.sv:18023:3
	wire [31:0] alu_operand_c_ex;
	// Trace: design.sv:18024:3
	wire [4:0] bmask_a_ex;
	// Trace: design.sv:18025:3
	wire [4:0] bmask_b_ex;
	// Trace: design.sv:18026:3
	wire [1:0] imm_vec_ext_ex;
	// Trace: design.sv:18027:3
	wire [1:0] alu_vec_mode_ex;
	// Trace: design.sv:18028:3
	wire alu_is_clpx_ex;
	wire alu_is_subrot_ex;
	// Trace: design.sv:18029:3
	wire [1:0] alu_clpx_shift_ex;
	// Trace: design.sv:18032:3
	localparam cv32e40p_pkg_MUL_OP_WIDTH = 3;
	// removed localparam type cv32e40p_pkg_mul_opcode_e
	wire [2:0] mult_operator_ex;
	// Trace: design.sv:18033:3
	wire [31:0] mult_operand_a_ex;
	// Trace: design.sv:18034:3
	wire [31:0] mult_operand_b_ex;
	// Trace: design.sv:18035:3
	wire [31:0] mult_operand_c_ex;
	// Trace: design.sv:18036:3
	wire mult_en_ex;
	// Trace: design.sv:18037:3
	wire mult_sel_subword_ex;
	// Trace: design.sv:18038:3
	wire [1:0] mult_signed_mode_ex;
	// Trace: design.sv:18039:3
	wire [4:0] mult_imm_ex;
	// Trace: design.sv:18040:3
	wire [31:0] mult_dot_op_a_ex;
	// Trace: design.sv:18041:3
	wire [31:0] mult_dot_op_b_ex;
	// Trace: design.sv:18042:3
	wire [31:0] mult_dot_op_c_ex;
	// Trace: design.sv:18043:3
	wire [1:0] mult_dot_signed_ex;
	// Trace: design.sv:18044:3
	wire mult_is_clpx_ex;
	// Trace: design.sv:18045:3
	wire [1:0] mult_clpx_shift_ex;
	// Trace: design.sv:18046:3
	wire mult_clpx_img_ex;
	// Trace: design.sv:18049:3
	localparam cv32e40p_pkg_C_RM = 3;
	wire [2:0] frm_csr;
	// Trace: design.sv:18050:3
	localparam cv32e40p_pkg_C_FFLAG = 5;
	wire [4:0] fflags_csr;
	// Trace: design.sv:18051:3
	wire fflags_we;
	// Trace: design.sv:18054:3
	wire apu_en_ex;
	// Trace: design.sv:18055:3
	wire [14:0] apu_flags_ex;
	// Trace: design.sv:18056:3
	wire [5:0] apu_op_ex;
	// Trace: design.sv:18057:3
	wire [1:0] apu_lat_ex;
	// Trace: design.sv:18058:3
	wire [95:0] apu_operands_ex;
	// Trace: design.sv:18059:3
	wire [5:0] apu_waddr_ex;
	// Trace: design.sv:18061:3
	wire [17:0] apu_read_regs;
	// Trace: design.sv:18062:3
	wire [2:0] apu_read_regs_valid;
	// Trace: design.sv:18063:3
	wire apu_read_dep;
	// Trace: design.sv:18064:3
	wire [11:0] apu_write_regs;
	// Trace: design.sv:18065:3
	wire [1:0] apu_write_regs_valid;
	// Trace: design.sv:18066:3
	wire apu_write_dep;
	// Trace: design.sv:18068:3
	wire perf_apu_type;
	// Trace: design.sv:18069:3
	wire perf_apu_cont;
	// Trace: design.sv:18070:3
	wire perf_apu_dep;
	// Trace: design.sv:18071:3
	wire perf_apu_wb;
	// Trace: design.sv:18074:3
	wire [5:0] regfile_waddr_ex;
	// Trace: design.sv:18075:3
	wire regfile_we_ex;
	// Trace: design.sv:18076:3
	wire [5:0] regfile_waddr_fw_wb_o;
	// Trace: design.sv:18077:3
	wire regfile_we_wb;
	// Trace: design.sv:18078:3
	wire [31:0] regfile_wdata;
	// Trace: design.sv:18080:3
	wire [5:0] regfile_alu_waddr_ex;
	// Trace: design.sv:18081:3
	wire regfile_alu_we_ex;
	// Trace: design.sv:18083:3
	wire [5:0] regfile_alu_waddr_fw;
	// Trace: design.sv:18084:3
	wire regfile_alu_we_fw;
	// Trace: design.sv:18085:3
	wire [31:0] regfile_alu_wdata_fw;
	// Trace: design.sv:18088:3
	wire csr_access_ex;
	// Trace: design.sv:18089:3
	localparam cv32e40p_pkg_CSR_OP_WIDTH = 2;
	// removed localparam type cv32e40p_pkg_csr_opcode_e
	wire [1:0] csr_op_ex;
	// Trace: design.sv:18090:3
	wire [23:0] mtvec;
	wire [23:0] utvec;
	// Trace: design.sv:18091:3
	wire [1:0] mtvec_mode;
	// Trace: design.sv:18092:3
	wire [1:0] utvec_mode;
	// Trace: design.sv:18094:3
	wire [1:0] csr_op;
	// Trace: design.sv:18095:3
	// removed localparam type cv32e40p_pkg_csr_num_e
	wire [11:0] csr_addr;
	// Trace: design.sv:18096:3
	wire [11:0] csr_addr_int;
	// Trace: design.sv:18097:3
	wire [31:0] csr_rdata;
	// Trace: design.sv:18098:3
	wire [31:0] csr_wdata;
	// Trace: design.sv:18099:3
	// removed localparam type cv32e40p_pkg_PrivLvl_t
	wire [1:0] current_priv_lvl;
	// Trace: design.sv:18102:3
	wire data_we_ex;
	// Trace: design.sv:18103:3
	wire [5:0] data_atop_ex;
	// Trace: design.sv:18104:3
	wire [1:0] data_type_ex;
	// Trace: design.sv:18105:3
	wire [1:0] data_sign_ext_ex;
	// Trace: design.sv:18106:3
	wire [1:0] data_reg_offset_ex;
	// Trace: design.sv:18107:3
	wire data_req_ex;
	// Trace: design.sv:18108:3
	wire data_load_event_ex;
	// Trace: design.sv:18109:3
	wire data_misaligned_ex;
	// Trace: design.sv:18111:3
	wire p_elw_start;
	// Trace: design.sv:18112:3
	wire p_elw_finish;
	// Trace: design.sv:18114:3
	wire [31:0] lsu_rdata;
	// Trace: design.sv:18117:3
	wire halt_if;
	// Trace: design.sv:18118:3
	wire id_ready;
	// Trace: design.sv:18119:3
	wire ex_ready;
	// Trace: design.sv:18121:3
	wire id_valid;
	// Trace: design.sv:18122:3
	wire ex_valid;
	// Trace: design.sv:18123:3
	wire wb_valid;
	// Trace: design.sv:18125:3
	wire lsu_ready_ex;
	// Trace: design.sv:18126:3
	wire lsu_ready_wb;
	// Trace: design.sv:18128:3
	wire apu_ready_wb;
	// Trace: design.sv:18131:3
	wire instr_req_int;
	// Trace: design.sv:18134:3
	wire m_irq_enable;
	wire u_irq_enable;
	// Trace: design.sv:18135:3
	wire csr_irq_sec;
	// Trace: design.sv:18136:3
	wire [31:0] mepc;
	wire [31:0] uepc;
	wire [31:0] depc;
	// Trace: design.sv:18137:3
	wire [31:0] mie_bypass;
	// Trace: design.sv:18138:3
	wire [31:0] mip;
	// Trace: design.sv:18140:3
	wire csr_save_cause;
	// Trace: design.sv:18141:3
	wire csr_save_if;
	// Trace: design.sv:18142:3
	wire csr_save_id;
	// Trace: design.sv:18143:3
	wire csr_save_ex;
	// Trace: design.sv:18144:3
	wire [5:0] csr_cause;
	// Trace: design.sv:18145:3
	wire csr_restore_mret_id;
	// Trace: design.sv:18146:3
	wire csr_restore_uret_id;
	// Trace: design.sv:18147:3
	wire csr_restore_dret_id;
	// Trace: design.sv:18148:3
	wire csr_mtvec_init;
	// Trace: design.sv:18151:3
	wire [31:0] mcounteren;
	// Trace: design.sv:18154:3
	wire debug_mode;
	// Trace: design.sv:18155:3
	wire [2:0] debug_cause;
	// Trace: design.sv:18156:3
	wire debug_csr_save;
	// Trace: design.sv:18157:3
	wire debug_single_step;
	// Trace: design.sv:18158:3
	wire debug_ebreakm;
	// Trace: design.sv:18159:3
	wire debug_ebreaku;
	// Trace: design.sv:18160:3
	wire trigger_match;
	// Trace: design.sv:18161:3
	wire debug_p_elw_no_sleep;
	// Trace: design.sv:18164:3
	wire [63:0] hwlp_start;
	// Trace: design.sv:18165:3
	wire [63:0] hwlp_end;
	// Trace: design.sv:18166:3
	wire [63:0] hwlp_cnt;
	// Trace: design.sv:18168:3
	wire [31:0] hwlp_target;
	// Trace: design.sv:18169:3
	wire hwlp_jump;
	// Trace: design.sv:18172:3
	wire [0:0] csr_hwlp_regid;
	// Trace: design.sv:18173:3
	wire [2:0] csr_hwlp_we;
	// Trace: design.sv:18174:3
	wire [31:0] csr_hwlp_data;
	// Trace: design.sv:18177:3
	wire mhpmevent_minstret;
	// Trace: design.sv:18178:3
	wire mhpmevent_load;
	// Trace: design.sv:18179:3
	wire mhpmevent_store;
	// Trace: design.sv:18180:3
	wire mhpmevent_jump;
	// Trace: design.sv:18181:3
	wire mhpmevent_branch;
	// Trace: design.sv:18182:3
	wire mhpmevent_branch_taken;
	// Trace: design.sv:18183:3
	wire mhpmevent_compressed;
	// Trace: design.sv:18184:3
	wire mhpmevent_jr_stall;
	// Trace: design.sv:18185:3
	wire mhpmevent_imiss;
	// Trace: design.sv:18186:3
	wire mhpmevent_ld_stall;
	// Trace: design.sv:18187:3
	wire mhpmevent_pipe_stall;
	// Trace: design.sv:18189:3
	wire perf_imiss;
	// Trace: design.sv:18192:3
	wire wake_from_sleep;
	// Trace: design.sv:18195:3
	wire [511:0] pmp_addr;
	// Trace: design.sv:18196:3
	wire [127:0] pmp_cfg;
	// Trace: design.sv:18198:3
	wire data_req_pmp;
	// Trace: design.sv:18199:3
	wire [31:0] data_addr_pmp;
	// Trace: design.sv:18200:3
	wire data_gnt_pmp;
	// Trace: design.sv:18201:3
	wire data_err_pmp;
	// Trace: design.sv:18202:3
	wire data_err_ack;
	// Trace: design.sv:18203:3
	wire instr_req_pmp;
	// Trace: design.sv:18204:3
	wire instr_gnt_pmp;
	// Trace: design.sv:18205:3
	wire [31:0] instr_addr_pmp;
	// Trace: design.sv:18206:3
	wire instr_err_pmp;
	// Trace: design.sv:18209:3
	assign m_exc_vec_pc_mux_id = (mtvec_mode == 2'b00 ? 5'h00 : exc_cause);
	// Trace: design.sv:18210:3
	assign u_exc_vec_pc_mux_id = (utvec_mode == 2'b00 ? 5'h00 : exc_cause);
	// Trace: design.sv:18213:3
	assign irq_sec_i = 1'b0;
	// Trace: design.sv:18216:3
	assign apu_flags_o = apu_flags_ex;
	// Trace: design.sv:18217:3
	assign fflags_csr = apu_flags_i;
	// Trace: design.sv:18228:3
	wire clk;
	// Trace: design.sv:18229:3
	wire fetch_enable;
	// Trace: design.sv:18231:3
	cv32e40p_sleep_unit #(.PULP_CLUSTER(PULP_CLUSTER)) sleep_unit_i(
		.clk_ungated_i(clk_i),
		.rst_n(rst_ni),
		.clk_gated_o(clk),
		.scan_cg_en_i(scan_cg_en_i),
		.core_sleep_o(core_sleep_o),
		.fetch_enable_i(fetch_enable_i),
		.fetch_enable_o(fetch_enable),
		.if_busy_i(if_busy),
		.ctrl_busy_i(ctrl_busy),
		.lsu_busy_i(lsu_busy),
		.apu_busy_i(apu_busy),
		.pulp_clock_en_i(pulp_clock_en_i),
		.p_elw_start_i(p_elw_start),
		.p_elw_finish_i(p_elw_finish),
		.debug_p_elw_no_sleep_i(debug_p_elw_no_sleep),
		.wake_from_sleep_i(wake_from_sleep)
	);
	// Trace: design.sv:18272:3
	cv32e40p_if_stage #(
		.PULP_XPULP(PULP_XPULP),
		.PULP_OBI(PULP_OBI),
		.PULP_SECURE(PULP_SECURE),
		.FPU(FPU)
	) if_stage_i(
		.clk(clk),
		.rst_n(rst_ni),
		.boot_addr_i(boot_addr_i[31:0]),
		.dm_exception_addr_i(dm_exception_addr_i[31:0]),
		.dm_halt_addr_i(dm_halt_addr_i[31:0]),
		.m_trap_base_addr_i(mtvec),
		.u_trap_base_addr_i(utvec),
		.trap_addr_mux_i(trap_addr_mux),
		.req_i(instr_req_int),
		.instr_req_o(instr_req_pmp),
		.instr_addr_o(instr_addr_pmp),
		.instr_gnt_i(instr_gnt_pmp),
		.instr_rvalid_i(instr_rvalid_i),
		.instr_rdata_i(instr_rdata_i),
		.instr_err_i(1'b0),
		.instr_err_pmp_i(instr_err_pmp),
		.instr_valid_id_o(instr_valid_id),
		.instr_rdata_id_o(instr_rdata_id),
		.is_fetch_failed_o(is_fetch_failed_id),
		.clear_instr_valid_i(clear_instr_valid),
		.pc_set_i(pc_set),
		.mepc_i(mepc),
		.uepc_i(uepc),
		.depc_i(depc),
		.pc_mux_i(pc_mux_id),
		.exc_pc_mux_i(exc_pc_mux_id),
		.pc_id_o(pc_id),
		.pc_if_o(pc_if),
		.is_compressed_id_o(is_compressed_id),
		.illegal_c_insn_id_o(illegal_c_insn_id),
		.m_exc_vec_pc_mux_i(m_exc_vec_pc_mux_id),
		.u_exc_vec_pc_mux_i(u_exc_vec_pc_mux_id),
		.csr_mtvec_init_o(csr_mtvec_init),
		.hwlp_jump_i(hwlp_jump),
		.hwlp_target_i(hwlp_target),
		.jump_target_id_i(jump_target_id),
		.jump_target_ex_i(jump_target_ex),
		.halt_if_i(halt_if),
		.id_ready_i(id_ready),
		.if_busy_o(if_busy),
		.perf_imiss_o(perf_imiss)
	);
	// Trace: design.sv:18360:3
	cv32e40p_id_stage #(
		.PULP_XPULP(PULP_XPULP),
		.PULP_CLUSTER(PULP_CLUSTER),
		.N_HWLP(N_HWLP),
		.PULP_SECURE(PULP_SECURE),
		.USE_PMP(USE_PMP),
		.A_EXTENSION(A_EXTENSION),
		.APU(APU),
		.FPU(FPU),
		.PULP_ZFINX(PULP_ZFINX),
		.APU_NARGS_CPU(cv32e40p_apu_core_pkg_APU_NARGS_CPU),
		.APU_WOP_CPU(cv32e40p_apu_core_pkg_APU_WOP_CPU),
		.APU_NDSFLAGS_CPU(cv32e40p_apu_core_pkg_APU_NDSFLAGS_CPU),
		.APU_NUSFLAGS_CPU(cv32e40p_apu_core_pkg_APU_NUSFLAGS_CPU),
		.DEBUG_TRIGGER_EN(DEBUG_TRIGGER_EN)
	) id_stage_i(
		.clk(clk),
		.clk_ungated_i(clk_i),
		.rst_n(rst_ni),
		.scan_cg_en_i(scan_cg_en_i),
		.fetch_enable_i(fetch_enable),
		.ctrl_busy_o(ctrl_busy),
		.is_decoding_o(is_decoding),
		.instr_valid_i(instr_valid_id),
		.instr_rdata_i(instr_rdata_id),
		.instr_req_o(instr_req_int),
		.branch_in_ex_o(branch_in_ex),
		.branch_decision_i(branch_decision),
		.jump_target_o(jump_target_id),
		.clear_instr_valid_o(clear_instr_valid),
		.pc_set_o(pc_set),
		.pc_mux_o(pc_mux_id),
		.exc_pc_mux_o(exc_pc_mux_id),
		.exc_cause_o(exc_cause),
		.trap_addr_mux_o(trap_addr_mux),
		.is_fetch_failed_i(is_fetch_failed_id),
		.pc_id_i(pc_id),
		.is_compressed_i(is_compressed_id),
		.illegal_c_insn_i(illegal_c_insn_id),
		.halt_if_o(halt_if),
		.id_ready_o(id_ready),
		.ex_ready_i(ex_ready),
		.wb_ready_i(lsu_ready_wb),
		.id_valid_o(id_valid),
		.ex_valid_i(ex_valid),
		.pc_ex_o(pc_ex),
		.alu_en_ex_o(alu_en_ex),
		.alu_operator_ex_o(alu_operator_ex),
		.alu_operand_a_ex_o(alu_operand_a_ex),
		.alu_operand_b_ex_o(alu_operand_b_ex),
		.alu_operand_c_ex_o(alu_operand_c_ex),
		.bmask_a_ex_o(bmask_a_ex),
		.bmask_b_ex_o(bmask_b_ex),
		.imm_vec_ext_ex_o(imm_vec_ext_ex),
		.alu_vec_mode_ex_o(alu_vec_mode_ex),
		.alu_is_clpx_ex_o(alu_is_clpx_ex),
		.alu_is_subrot_ex_o(alu_is_subrot_ex),
		.alu_clpx_shift_ex_o(alu_clpx_shift_ex),
		.regfile_waddr_ex_o(regfile_waddr_ex),
		.regfile_we_ex_o(regfile_we_ex),
		.regfile_alu_we_ex_o(regfile_alu_we_ex),
		.regfile_alu_waddr_ex_o(regfile_alu_waddr_ex),
		.mult_operator_ex_o(mult_operator_ex),
		.mult_en_ex_o(mult_en_ex),
		.mult_sel_subword_ex_o(mult_sel_subword_ex),
		.mult_signed_mode_ex_o(mult_signed_mode_ex),
		.mult_operand_a_ex_o(mult_operand_a_ex),
		.mult_operand_b_ex_o(mult_operand_b_ex),
		.mult_operand_c_ex_o(mult_operand_c_ex),
		.mult_imm_ex_o(mult_imm_ex),
		.mult_dot_op_a_ex_o(mult_dot_op_a_ex),
		.mult_dot_op_b_ex_o(mult_dot_op_b_ex),
		.mult_dot_op_c_ex_o(mult_dot_op_c_ex),
		.mult_dot_signed_ex_o(mult_dot_signed_ex),
		.mult_is_clpx_ex_o(mult_is_clpx_ex),
		.mult_clpx_shift_ex_o(mult_clpx_shift_ex),
		.mult_clpx_img_ex_o(mult_clpx_img_ex),
		.frm_i(frm_csr),
		.apu_en_ex_o(apu_en_ex),
		.apu_op_ex_o(apu_op_ex),
		.apu_lat_ex_o(apu_lat_ex),
		.apu_operands_ex_o(apu_operands_ex),
		.apu_flags_ex_o(apu_flags_ex),
		.apu_waddr_ex_o(apu_waddr_ex),
		.apu_read_regs_o(apu_read_regs),
		.apu_read_regs_valid_o(apu_read_regs_valid),
		.apu_read_dep_i(apu_read_dep),
		.apu_write_regs_o(apu_write_regs),
		.apu_write_regs_valid_o(apu_write_regs_valid),
		.apu_write_dep_i(apu_write_dep),
		.apu_perf_dep_o(perf_apu_dep),
		.apu_busy_i(apu_busy),
		.csr_access_ex_o(csr_access_ex),
		.csr_op_ex_o(csr_op_ex),
		.current_priv_lvl_i(current_priv_lvl),
		.csr_irq_sec_o(csr_irq_sec),
		.csr_cause_o(csr_cause),
		.csr_save_if_o(csr_save_if),
		.csr_save_id_o(csr_save_id),
		.csr_save_ex_o(csr_save_ex),
		.csr_restore_mret_id_o(csr_restore_mret_id),
		.csr_restore_uret_id_o(csr_restore_uret_id),
		.csr_restore_dret_id_o(csr_restore_dret_id),
		.csr_save_cause_o(csr_save_cause),
		.hwlp_start_o(hwlp_start),
		.hwlp_end_o(hwlp_end),
		.hwlp_cnt_o(hwlp_cnt),
		.hwlp_jump_o(hwlp_jump),
		.hwlp_target_o(hwlp_target),
		.csr_hwlp_regid_i(csr_hwlp_regid),
		.csr_hwlp_we_i(csr_hwlp_we),
		.csr_hwlp_data_i(csr_hwlp_data),
		.data_req_ex_o(data_req_ex),
		.data_we_ex_o(data_we_ex),
		.atop_ex_o(data_atop_ex),
		.data_type_ex_o(data_type_ex),
		.data_sign_ext_ex_o(data_sign_ext_ex),
		.data_reg_offset_ex_o(data_reg_offset_ex),
		.data_load_event_ex_o(data_load_event_ex),
		.data_misaligned_ex_o(data_misaligned_ex),
		.prepost_useincr_ex_o(useincr_addr_ex),
		.data_misaligned_i(data_misaligned),
		.data_err_i(data_err_pmp),
		.data_err_ack_o(data_err_ack),
		.irq_i(irq_i),
		.irq_sec_i((PULP_SECURE ? irq_sec_i : 1'b0)),
		.mie_bypass_i(mie_bypass),
		.mip_o(mip),
		.m_irq_enable_i(m_irq_enable),
		.u_irq_enable_i(u_irq_enable),
		.irq_ack_o(irq_ack_o),
		.irq_id_o(irq_id_o),
		.debug_mode_o(debug_mode),
		.debug_cause_o(debug_cause),
		.debug_csr_save_o(debug_csr_save),
		.debug_req_i(debug_req_i),
		.debug_havereset_o(debug_havereset_o),
		.debug_running_o(debug_running_o),
		.debug_halted_o(debug_halted_o),
		.debug_single_step_i(debug_single_step),
		.debug_ebreakm_i(debug_ebreakm),
		.debug_ebreaku_i(debug_ebreaku),
		.trigger_match_i(trigger_match),
		.debug_p_elw_no_sleep_o(debug_p_elw_no_sleep),
		.wake_from_sleep_o(wake_from_sleep),
		.regfile_waddr_wb_i(regfile_waddr_fw_wb_o),
		.regfile_we_wb_i(regfile_we_wb),
		.regfile_wdata_wb_i(regfile_wdata),
		.regfile_alu_waddr_fw_i(regfile_alu_waddr_fw),
		.regfile_alu_we_fw_i(regfile_alu_we_fw),
		.regfile_alu_wdata_fw_i(regfile_alu_wdata_fw),
		.mult_multicycle_i(mult_multicycle),
		.mhpmevent_minstret_o(mhpmevent_minstret),
		.mhpmevent_load_o(mhpmevent_load),
		.mhpmevent_store_o(mhpmevent_store),
		.mhpmevent_jump_o(mhpmevent_jump),
		.mhpmevent_branch_o(mhpmevent_branch),
		.mhpmevent_branch_taken_o(mhpmevent_branch_taken),
		.mhpmevent_compressed_o(mhpmevent_compressed),
		.mhpmevent_jr_stall_o(mhpmevent_jr_stall),
		.mhpmevent_imiss_o(mhpmevent_imiss),
		.mhpmevent_ld_stall_o(mhpmevent_ld_stall),
		.mhpmevent_pipe_stall_o(mhpmevent_pipe_stall),
		.perf_imiss_i(perf_imiss),
		.mcounteren_i(mcounteren)
	);
	// Trace: design.sv:18592:3
	cv32e40p_ex_stage #(
		.FPU(FPU),
		.APU_NARGS_CPU(cv32e40p_apu_core_pkg_APU_NARGS_CPU),
		.APU_WOP_CPU(cv32e40p_apu_core_pkg_APU_WOP_CPU),
		.APU_NDSFLAGS_CPU(cv32e40p_apu_core_pkg_APU_NDSFLAGS_CPU),
		.APU_NUSFLAGS_CPU(cv32e40p_apu_core_pkg_APU_NUSFLAGS_CPU)
	) ex_stage_i(
		.clk(clk),
		.rst_n(rst_ni),
		.alu_en_i(alu_en_ex),
		.alu_operator_i(alu_operator_ex),
		.alu_operand_a_i(alu_operand_a_ex),
		.alu_operand_b_i(alu_operand_b_ex),
		.alu_operand_c_i(alu_operand_c_ex),
		.bmask_a_i(bmask_a_ex),
		.bmask_b_i(bmask_b_ex),
		.imm_vec_ext_i(imm_vec_ext_ex),
		.alu_vec_mode_i(alu_vec_mode_ex),
		.alu_is_clpx_i(alu_is_clpx_ex),
		.alu_is_subrot_i(alu_is_subrot_ex),
		.alu_clpx_shift_i(alu_clpx_shift_ex),
		.mult_operator_i(mult_operator_ex),
		.mult_operand_a_i(mult_operand_a_ex),
		.mult_operand_b_i(mult_operand_b_ex),
		.mult_operand_c_i(mult_operand_c_ex),
		.mult_en_i(mult_en_ex),
		.mult_sel_subword_i(mult_sel_subword_ex),
		.mult_signed_mode_i(mult_signed_mode_ex),
		.mult_imm_i(mult_imm_ex),
		.mult_dot_op_a_i(mult_dot_op_a_ex),
		.mult_dot_op_b_i(mult_dot_op_b_ex),
		.mult_dot_op_c_i(mult_dot_op_c_ex),
		.mult_dot_signed_i(mult_dot_signed_ex),
		.mult_is_clpx_i(mult_is_clpx_ex),
		.mult_clpx_shift_i(mult_clpx_shift_ex),
		.mult_clpx_img_i(mult_clpx_img_ex),
		.mult_multicycle_o(mult_multicycle),
		.fpu_fflags_we_o(fflags_we),
		.apu_en_i(apu_en_ex),
		.apu_op_i(apu_op_ex),
		.apu_lat_i(apu_lat_ex),
		.apu_operands_i(apu_operands_ex),
		.apu_waddr_i(apu_waddr_ex),
		.apu_flags_i(apu_flags_ex),
		.apu_read_regs_i(apu_read_regs),
		.apu_read_regs_valid_i(apu_read_regs_valid),
		.apu_read_dep_o(apu_read_dep),
		.apu_write_regs_i(apu_write_regs),
		.apu_write_regs_valid_i(apu_write_regs_valid),
		.apu_write_dep_o(apu_write_dep),
		.apu_perf_type_o(perf_apu_type),
		.apu_perf_cont_o(perf_apu_cont),
		.apu_perf_wb_o(perf_apu_wb),
		.apu_ready_wb_o(apu_ready_wb),
		.apu_busy_o(apu_busy),
		.apu_req_o(apu_req_o),
		.apu_gnt_i(apu_gnt_i),
		.apu_operands_o(apu_operands_o),
		.apu_op_o(apu_op_o),
		.apu_rvalid_i(apu_rvalid_i),
		.apu_result_i(apu_result_i),
		.lsu_en_i(data_req_ex),
		.lsu_rdata_i(lsu_rdata),
		.csr_access_i(csr_access_ex),
		.csr_rdata_i(csr_rdata),
		.branch_in_ex_i(branch_in_ex),
		.regfile_alu_waddr_i(regfile_alu_waddr_ex),
		.regfile_alu_we_i(regfile_alu_we_ex),
		.regfile_waddr_i(regfile_waddr_ex),
		.regfile_we_i(regfile_we_ex),
		.regfile_waddr_wb_o(regfile_waddr_fw_wb_o),
		.regfile_we_wb_o(regfile_we_wb),
		.regfile_wdata_wb_o(regfile_wdata),
		.jump_target_o(jump_target_ex),
		.branch_decision_o(branch_decision),
		.regfile_alu_waddr_fw_o(regfile_alu_waddr_fw),
		.regfile_alu_we_fw_o(regfile_alu_we_fw),
		.regfile_alu_wdata_fw_o(regfile_alu_wdata_fw),
		.is_decoding_i(is_decoding),
		.lsu_ready_ex_i(lsu_ready_ex),
		.lsu_err_i(data_err_pmp),
		.ex_ready_o(ex_ready),
		.ex_valid_o(ex_valid),
		.wb_ready_i(lsu_ready_wb)
	);
	// Trace: design.sv:18720:3
	cv32e40p_load_store_unit #(.PULP_OBI(PULP_OBI)) load_store_unit_i(
		.clk(clk),
		.rst_n(rst_ni),
		.data_req_o(data_req_pmp),
		.data_gnt_i(data_gnt_pmp),
		.data_rvalid_i(data_rvalid_i),
		.data_err_i(1'b0),
		.data_err_pmp_i(data_err_pmp),
		.data_addr_o(data_addr_pmp),
		.data_we_o(data_we_o),
		.data_atop_o(data_atop_o),
		.data_be_o(data_be_o),
		.data_wdata_o(data_wdata_o),
		.data_rdata_i(data_rdata_i),
		.data_we_ex_i(data_we_ex),
		.data_atop_ex_i(data_atop_ex),
		.data_type_ex_i(data_type_ex),
		.data_wdata_ex_i(alu_operand_c_ex),
		.data_reg_offset_ex_i(data_reg_offset_ex),
		.data_load_event_ex_i(data_load_event_ex),
		.data_sign_ext_ex_i(data_sign_ext_ex),
		.data_rdata_ex_o(lsu_rdata),
		.data_req_ex_i(data_req_ex),
		.operand_a_ex_i(alu_operand_a_ex),
		.operand_b_ex_i(alu_operand_b_ex),
		.addr_useincr_ex_i(useincr_addr_ex),
		.data_misaligned_ex_i(data_misaligned_ex),
		.data_misaligned_o(data_misaligned),
		.p_elw_start_o(p_elw_start),
		.p_elw_finish_o(p_elw_finish),
		.lsu_ready_ex_o(lsu_ready_ex),
		.lsu_ready_wb_o(lsu_ready_wb),
		.busy_o(lsu_busy)
	);
	// Trace: design.sv:18769:3
	assign wb_valid = lsu_ready_wb;
	// Trace: design.sv:18782:3
	cv32e40p_cs_registers #(
		.A_EXTENSION(A_EXTENSION),
		.FPU(FPU),
		.APU(APU),
		.PULP_SECURE(PULP_SECURE),
		.USE_PMP(USE_PMP),
		.N_PMP_ENTRIES(N_PMP_ENTRIES),
		.NUM_MHPMCOUNTERS(NUM_MHPMCOUNTERS),
		.PULP_XPULP(PULP_XPULP),
		.PULP_CLUSTER(PULP_CLUSTER),
		.DEBUG_TRIGGER_EN(DEBUG_TRIGGER_EN)
	) cs_registers_i(
		.clk(clk),
		.rst_n(rst_ni),
		.hart_id_i(hart_id_i),
		.mtvec_o(mtvec),
		.utvec_o(utvec),
		.mtvec_mode_o(mtvec_mode),
		.utvec_mode_o(utvec_mode),
		.mtvec_addr_i(mtvec_addr_i[31:0]),
		.csr_mtvec_init_i(csr_mtvec_init),
		.csr_addr_i(csr_addr),
		.csr_wdata_i(csr_wdata),
		.csr_op_i(csr_op),
		.csr_rdata_o(csr_rdata),
		.frm_o(frm_csr),
		.fflags_i(fflags_csr),
		.fflags_we_i(fflags_we),
		.mie_bypass_o(mie_bypass),
		.mip_i(mip),
		.m_irq_enable_o(m_irq_enable),
		.u_irq_enable_o(u_irq_enable),
		.csr_irq_sec_i(csr_irq_sec),
		.sec_lvl_o(sec_lvl_o),
		.mepc_o(mepc),
		.uepc_o(uepc),
		.mcounteren_o(mcounteren),
		.debug_mode_i(debug_mode),
		.debug_cause_i(debug_cause),
		.debug_csr_save_i(debug_csr_save),
		.depc_o(depc),
		.debug_single_step_o(debug_single_step),
		.debug_ebreakm_o(debug_ebreakm),
		.debug_ebreaku_o(debug_ebreaku),
		.trigger_match_o(trigger_match),
		.priv_lvl_o(current_priv_lvl),
		.pmp_addr_o(pmp_addr),
		.pmp_cfg_o(pmp_cfg),
		.pc_if_i(pc_if),
		.pc_id_i(pc_id),
		.pc_ex_i(pc_ex),
		.csr_save_if_i(csr_save_if),
		.csr_save_id_i(csr_save_id),
		.csr_save_ex_i(csr_save_ex),
		.csr_restore_mret_i(csr_restore_mret_id),
		.csr_restore_uret_i(csr_restore_uret_id),
		.csr_restore_dret_i(csr_restore_dret_id),
		.csr_cause_i(csr_cause),
		.csr_save_cause_i(csr_save_cause),
		.hwlp_start_i(hwlp_start),
		.hwlp_end_i(hwlp_end),
		.hwlp_cnt_i(hwlp_cnt),
		.hwlp_regid_o(csr_hwlp_regid),
		.hwlp_we_o(csr_hwlp_we),
		.hwlp_data_o(csr_hwlp_data),
		.mhpmevent_minstret_i(mhpmevent_minstret),
		.mhpmevent_load_i(mhpmevent_load),
		.mhpmevent_store_i(mhpmevent_store),
		.mhpmevent_jump_i(mhpmevent_jump),
		.mhpmevent_branch_i(mhpmevent_branch),
		.mhpmevent_branch_taken_i(mhpmevent_branch_taken),
		.mhpmevent_compressed_i(mhpmevent_compressed),
		.mhpmevent_jr_stall_i(mhpmevent_jr_stall),
		.mhpmevent_imiss_i(mhpmevent_imiss),
		.mhpmevent_ld_stall_i(mhpmevent_ld_stall),
		.mhpmevent_pipe_stall_i(mhpmevent_pipe_stall),
		.apu_typeconflict_i(perf_apu_type),
		.apu_contention_i(perf_apu_cont),
		.apu_dep_i(perf_apu_dep),
		.apu_wb_i(perf_apu_wb)
	);
	// Trace: design.sv:18887:3
	assign csr_addr = csr_addr_int;
	// Trace: design.sv:18888:3
	assign csr_wdata = alu_operand_a_ex;
	// Trace: design.sv:18889:3
	assign csr_op = csr_op_ex;
	// Trace: design.sv:18891:3
	function automatic [11:0] sv2v_cast_12;
		input reg [11:0] inp;
		sv2v_cast_12 = inp;
	endfunction
	assign csr_addr_int = sv2v_cast_12((csr_access_ex ? alu_operand_b_ex[11:0] : {12 {1'sb0}}));
	// Trace: design.sv:18904:3
	generate
		if (1) begin : gen_no_pmp
			// Trace: design.sv:18939:7
			assign instr_req_o = instr_req_pmp;
			// Trace: design.sv:18940:7
			assign instr_addr_o = instr_addr_pmp;
			// Trace: design.sv:18941:7
			assign instr_gnt_pmp = instr_gnt_i;
			// Trace: design.sv:18942:7
			assign instr_err_pmp = 1'b0;
			// Trace: design.sv:18944:7
			assign data_req_o = data_req_pmp;
			// Trace: design.sv:18945:7
			assign data_addr_o = data_addr_pmp;
			// Trace: design.sv:18946:7
			assign data_gnt_pmp = data_gnt_i;
			// Trace: design.sv:18947:7
			assign data_err_pmp = 1'b0;
		end
	endgenerate
endmodule
module cv32e40p_apu_disp (
	clk_i,
	rst_ni,
	enable_i,
	apu_lat_i,
	apu_waddr_i,
	apu_waddr_o,
	apu_multicycle_o,
	apu_singlecycle_o,
	active_o,
	stall_o,
	is_decoding_i,
	read_regs_i,
	read_regs_valid_i,
	read_dep_o,
	write_regs_i,
	write_regs_valid_i,
	write_dep_o,
	perf_type_o,
	perf_cont_o,
	apu_req_o,
	apu_gnt_i,
	apu_rvalid_i
);
	reg _sv2v_0;
	// Trace: design.sv:19166:5
	input wire clk_i;
	// Trace: design.sv:19167:5
	input wire rst_ni;
	// Trace: design.sv:19170:5
	input wire enable_i;
	// Trace: design.sv:19171:5
	input wire [1:0] apu_lat_i;
	// Trace: design.sv:19172:5
	input wire [5:0] apu_waddr_i;
	// Trace: design.sv:19175:5
	output reg [5:0] apu_waddr_o;
	// Trace: design.sv:19176:5
	output wire apu_multicycle_o;
	// Trace: design.sv:19177:5
	output wire apu_singlecycle_o;
	// Trace: design.sv:19180:5
	output wire active_o;
	// Trace: design.sv:19183:5
	output wire stall_o;
	// Trace: design.sv:19186:5
	input wire is_decoding_i;
	// Trace: design.sv:19187:5
	input wire [17:0] read_regs_i;
	// Trace: design.sv:19188:5
	input wire [2:0] read_regs_valid_i;
	// Trace: design.sv:19189:5
	output wire read_dep_o;
	// Trace: design.sv:19191:5
	input wire [11:0] write_regs_i;
	// Trace: design.sv:19192:5
	input wire [1:0] write_regs_valid_i;
	// Trace: design.sv:19193:5
	output wire write_dep_o;
	// Trace: design.sv:19196:5
	output wire perf_type_o;
	// Trace: design.sv:19197:5
	output wire perf_cont_o;
	// Trace: design.sv:19201:5
	output wire apu_req_o;
	// Trace: design.sv:19202:5
	input wire apu_gnt_i;
	// Trace: design.sv:19204:5
	input wire apu_rvalid_i;
	// Trace: design.sv:19208:3
	wire [5:0] addr_req;
	reg [5:0] addr_inflight;
	reg [5:0] addr_waiting;
	// Trace: design.sv:19209:3
	reg [5:0] addr_inflight_dn;
	reg [5:0] addr_waiting_dn;
	// Trace: design.sv:19210:3
	wire valid_req;
	reg valid_inflight;
	reg valid_waiting;
	// Trace: design.sv:19211:3
	reg valid_inflight_dn;
	reg valid_waiting_dn;
	// Trace: design.sv:19212:3
	wire returned_req;
	wire returned_inflight;
	wire returned_waiting;
	// Trace: design.sv:19214:3
	wire req_accepted;
	// Trace: design.sv:19215:3
	wire active;
	// Trace: design.sv:19216:3
	reg [1:0] apu_lat;
	// Trace: design.sv:19219:3
	wire [2:0] read_deps_req;
	wire [2:0] read_deps_inflight;
	wire [2:0] read_deps_waiting;
	// Trace: design.sv:19220:3
	wire [1:0] write_deps_req;
	wire [1:0] write_deps_inflight;
	wire [1:0] write_deps_waiting;
	// Trace: design.sv:19221:3
	wire read_dep_req;
	wire read_dep_inflight;
	wire read_dep_waiting;
	// Trace: design.sv:19222:3
	wire write_dep_req;
	wire write_dep_inflight;
	wire write_dep_waiting;
	// Trace: design.sv:19224:3
	wire stall_full;
	wire stall_type;
	wire stall_nack;
	// Trace: design.sv:19227:3
	assign valid_req = enable_i & !(stall_full | stall_type);
	// Trace: design.sv:19228:3
	assign addr_req = apu_waddr_i;
	// Trace: design.sv:19230:3
	assign req_accepted = valid_req & apu_gnt_i;
	// Trace: design.sv:19236:3
	assign returned_req = ((valid_req & apu_rvalid_i) & !valid_inflight) & !valid_waiting;
	// Trace: design.sv:19237:3
	assign returned_inflight = (valid_inflight & apu_rvalid_i) & !valid_waiting;
	// Trace: design.sv:19238:3
	assign returned_waiting = valid_waiting & apu_rvalid_i;
	// Trace: design.sv:19241:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:19242:5
		if (~rst_ni) begin
			// Trace: design.sv:19243:7
			valid_inflight <= 1'b0;
			// Trace: design.sv:19244:7
			valid_waiting <= 1'b0;
			// Trace: design.sv:19245:7
			addr_inflight <= 1'sb0;
			// Trace: design.sv:19246:7
			addr_waiting <= 1'sb0;
		end
		else begin
			// Trace: design.sv:19248:7
			valid_inflight <= valid_inflight_dn;
			// Trace: design.sv:19249:7
			valid_waiting <= valid_waiting_dn;
			// Trace: design.sv:19250:7
			addr_inflight <= addr_inflight_dn;
			// Trace: design.sv:19251:7
			addr_waiting <= addr_waiting_dn;
		end
	// Trace: design.sv:19255:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:19256:5
		valid_inflight_dn = valid_inflight;
		// Trace: design.sv:19257:5
		valid_waiting_dn = valid_waiting;
		// Trace: design.sv:19258:5
		addr_inflight_dn = addr_inflight;
		// Trace: design.sv:19259:5
		addr_waiting_dn = addr_waiting;
		// Trace: design.sv:19261:5
		if (req_accepted & !returned_req) begin
			// Trace: design.sv:19262:7
			valid_inflight_dn = 1'b1;
			// Trace: design.sv:19263:7
			addr_inflight_dn = addr_req;
			// Trace: design.sv:19264:7
			if (valid_inflight & !returned_inflight) begin
				// Trace: design.sv:19265:9
				valid_waiting_dn = 1'b1;
				// Trace: design.sv:19266:9
				addr_waiting_dn = addr_inflight;
			end
			if (returned_waiting) begin
				// Trace: design.sv:19269:9
				valid_waiting_dn = 1'b1;
				// Trace: design.sv:19270:9
				addr_waiting_dn = addr_inflight;
			end
		end
		else if (returned_inflight) begin
			// Trace: design.sv:19274:7
			valid_inflight_dn = 1'sb0;
			// Trace: design.sv:19275:7
			valid_waiting_dn = 1'sb0;
			// Trace: design.sv:19276:7
			addr_inflight_dn = 1'sb0;
			// Trace: design.sv:19277:7
			addr_waiting_dn = 1'sb0;
		end
		else if (returned_waiting) begin
			// Trace: design.sv:19279:7
			valid_waiting_dn = 1'sb0;
			// Trace: design.sv:19280:7
			addr_waiting_dn = 1'sb0;
		end
	end
	// Trace: design.sv:19288:3
	assign active = valid_inflight | valid_waiting;
	// Trace: design.sv:19291:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:19292:5
		if (~rst_ni)
			// Trace: design.sv:19293:7
			apu_lat <= 1'sb0;
		else
			// Trace: design.sv:19295:7
			if (valid_req)
				// Trace: design.sv:19296:9
				apu_lat <= apu_lat_i;
	// Trace: design.sv:19305:3
	genvar _gv_i_3;
	generate
		for (_gv_i_3 = 0; _gv_i_3 < 3; _gv_i_3 = _gv_i_3 + 1) begin : gen_read_deps
			localparam i = _gv_i_3;
			// Trace: design.sv:19307:7
			assign read_deps_req[i] = (read_regs_i[i * 6+:6] == addr_req) & read_regs_valid_i[i];
			// Trace: design.sv:19308:7
			assign read_deps_inflight[i] = (read_regs_i[i * 6+:6] == addr_inflight) & read_regs_valid_i[i];
			// Trace: design.sv:19309:7
			assign read_deps_waiting[i] = (read_regs_i[i * 6+:6] == addr_waiting) & read_regs_valid_i[i];
		end
	endgenerate
	// Trace: design.sv:19313:3
	genvar _gv_i_4;
	generate
		for (_gv_i_4 = 0; _gv_i_4 < 2; _gv_i_4 = _gv_i_4 + 1) begin : gen_write_deps
			localparam i = _gv_i_4;
			// Trace: design.sv:19315:7
			assign write_deps_req[i] = (write_regs_i[i * 6+:6] == addr_req) & write_regs_valid_i[i];
			// Trace: design.sv:19316:7
			assign write_deps_inflight[i] = (write_regs_i[i * 6+:6] == addr_inflight) & write_regs_valid_i[i];
			// Trace: design.sv:19317:7
			assign write_deps_waiting[i] = (write_regs_i[i * 6+:6] == addr_waiting) & write_regs_valid_i[i];
		end
	endgenerate
	// Trace: design.sv:19322:3
	assign read_dep_req = (|read_deps_req & valid_req) & !returned_req;
	// Trace: design.sv:19323:3
	assign read_dep_inflight = (|read_deps_inflight & valid_inflight) & !returned_inflight;
	// Trace: design.sv:19324:3
	assign read_dep_waiting = (|read_deps_waiting & valid_waiting) & !returned_waiting;
	// Trace: design.sv:19325:3
	assign write_dep_req = (|write_deps_req & valid_req) & !returned_req;
	// Trace: design.sv:19326:3
	assign write_dep_inflight = (|write_deps_inflight & valid_inflight) & !returned_inflight;
	// Trace: design.sv:19327:3
	assign write_dep_waiting = (|write_deps_waiting & valid_waiting) & !returned_waiting;
	// Trace: design.sv:19329:3
	assign read_dep_o = ((read_dep_req | read_dep_inflight) | read_dep_waiting) & is_decoding_i;
	// Trace: design.sv:19330:3
	assign write_dep_o = ((write_dep_req | write_dep_inflight) | write_dep_waiting) & is_decoding_i;
	// Trace: design.sv:19336:3
	assign stall_full = valid_inflight & valid_waiting;
	// Trace: design.sv:19340:3
	assign stall_type = (enable_i & active) & (((apu_lat_i == 2'h1) | ((apu_lat_i == 2'h2) & (apu_lat == 2'h3))) | (apu_lat_i == 2'h3));
	// Trace: design.sv:19341:3
	assign stall_nack = valid_req & !apu_gnt_i;
	// Trace: design.sv:19342:3
	assign stall_o = (stall_full | stall_type) | stall_nack;
	// Trace: design.sv:19347:3
	assign apu_req_o = valid_req;
	// Trace: design.sv:19351:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:19352:5
		apu_waddr_o = 1'sb0;
		// Trace: design.sv:19353:5
		if (returned_req)
			// Trace: design.sv:19353:23
			apu_waddr_o = addr_req;
		if (returned_inflight)
			// Trace: design.sv:19354:28
			apu_waddr_o = addr_inflight;
		if (returned_waiting)
			// Trace: design.sv:19355:27
			apu_waddr_o = addr_waiting;
	end
	// Trace: design.sv:19359:3
	assign active_o = active;
	// Trace: design.sv:19362:3
	assign perf_type_o = stall_type;
	// Trace: design.sv:19363:3
	assign perf_cont_o = stall_nack;
	// Trace: design.sv:19365:3
	assign apu_multicycle_o = apu_lat == 2'h3;
	// Trace: design.sv:19366:3
	assign apu_singlecycle_o = ~(valid_inflight | valid_waiting);
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_fifo (
	clk_i,
	rst_ni,
	flush_i,
	flush_but_first_i,
	testmode_i,
	full_o,
	empty_o,
	cnt_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	reg _sv2v_0;
	// Trace: design.sv:19393:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:19394:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:19395:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:19397:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:19399:5
	input wire clk_i;
	// Trace: design.sv:19400:5
	input wire rst_ni;
	// Trace: design.sv:19401:5
	input wire flush_i;
	// Trace: design.sv:19402:5
	input wire flush_but_first_i;
	// Trace: design.sv:19403:5
	input wire testmode_i;
	// Trace: design.sv:19405:5
	output wire full_o;
	// Trace: design.sv:19406:5
	output wire empty_o;
	// Trace: design.sv:19407:5
	output wire [ADDR_DEPTH:0] cnt_o;
	// Trace: design.sv:19409:5
	input wire [DATA_WIDTH - 1:0] data_i;
	// Trace: design.sv:19410:5
	input wire push_i;
	// Trace: design.sv:19412:5
	output reg [DATA_WIDTH - 1:0] data_o;
	// Trace: design.sv:19413:5
	input wire pop_i;
	// Trace: design.sv:19417:3
	localparam [31:0] FIFO_DEPTH = (DEPTH > 0 ? DEPTH : 1);
	// Trace: design.sv:19419:3
	reg gate_clock;
	// Trace: design.sv:19421:3
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	// Trace: design.sv:19423:3
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	// Trace: design.sv:19426:3
	reg [(FIFO_DEPTH * DATA_WIDTH) - 1:0] mem_n;
	reg [(FIFO_DEPTH * DATA_WIDTH) - 1:0] mem_q;
	// Trace: design.sv:19428:3
	assign cnt_o = status_cnt_q;
	// Trace: design.sv:19431:3
	generate
		if (DEPTH == 0) begin : gen_zero_depth
			// Trace: design.sv:19433:7
			assign empty_o = ~push_i;
			// Trace: design.sv:19434:7
			assign full_o = ~pop_i;
		end
		else begin : gen_non_zero_depth
			// Trace: design.sv:19436:7
			assign full_o = status_cnt_q == FIFO_DEPTH[ADDR_DEPTH:0];
			// Trace: design.sv:19437:7
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	// Trace: design.sv:19442:3
	always @(*) begin : read_write_comb
		if (_sv2v_0)
			;
		// Trace: design.sv:19444:5
		read_pointer_n = read_pointer_q;
		// Trace: design.sv:19445:5
		write_pointer_n = write_pointer_q;
		// Trace: design.sv:19446:5
		status_cnt_n = status_cnt_q;
		// Trace: design.sv:19447:5
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q * DATA_WIDTH+:DATA_WIDTH]);
		// Trace: design.sv:19448:5
		mem_n = mem_q;
		// Trace: design.sv:19449:5
		gate_clock = 1'b1;
		// Trace: design.sv:19452:5
		if (push_i && ~full_o) begin
			// Trace: design.sv:19454:7
			mem_n[write_pointer_q * DATA_WIDTH+:DATA_WIDTH] = data_i;
			// Trace: design.sv:19456:7
			gate_clock = 1'b0;
			// Trace: design.sv:19458:7
			if (write_pointer_q == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:19458:62
				write_pointer_n = 1'sb0;
			else
				// Trace: design.sv:19459:12
				write_pointer_n = write_pointer_q + 1;
			// Trace: design.sv:19461:7
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			// Trace: design.sv:19467:7
			if (read_pointer_n == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:19467:61
				read_pointer_n = 1'sb0;
			else
				// Trace: design.sv:19468:12
				read_pointer_n = read_pointer_q + 1;
			// Trace: design.sv:19470:7
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			// Trace: design.sv:19474:49
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			// Trace: design.sv:19478:7
			data_o = data_i;
			// Trace: design.sv:19479:7
			if (pop_i) begin
				// Trace: design.sv:19480:9
				status_cnt_n = status_cnt_q;
				// Trace: design.sv:19481:9
				read_pointer_n = read_pointer_q;
				// Trace: design.sv:19482:9
				write_pointer_n = write_pointer_q;
			end
		end
	end
	// Trace: design.sv:19488:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:19489:5
		if (~rst_ni) begin
			// Trace: design.sv:19490:7
			read_pointer_q <= 1'sb0;
			// Trace: design.sv:19491:7
			write_pointer_q <= 1'sb0;
			// Trace: design.sv:19492:7
			status_cnt_q <= 1'sb0;
		end
		else
			// Trace: design.sv:19494:7
			(* full_case, parallel_case *)
			case (1'b1)
				flush_i: begin
					// Trace: design.sv:19497:11
					read_pointer_q <= 1'sb0;
					// Trace: design.sv:19498:11
					write_pointer_q <= 1'sb0;
					// Trace: design.sv:19499:11
					status_cnt_q <= 1'sb0;
				end
				flush_but_first_i: begin
					// Trace: design.sv:19503:11
					read_pointer_q <= (status_cnt_q > 0 ? read_pointer_q : {ADDR_DEPTH {1'sb0}});
					// Trace: design.sv:19504:11
					write_pointer_q <= (status_cnt_q > 0 ? read_pointer_q + 1 : {ADDR_DEPTH {1'sb0}});
					// Trace: design.sv:19505:11
					status_cnt_q <= (status_cnt_q > 0 ? 1'b1 : {(ADDR_DEPTH >= 0 ? ADDR_DEPTH + 1 : 1 - ADDR_DEPTH) {1'sb0}});
				end
				default: begin
					// Trace: design.sv:19509:11
					read_pointer_q <= read_pointer_n;
					// Trace: design.sv:19510:11
					write_pointer_q <= write_pointer_n;
					// Trace: design.sv:19511:11
					status_cnt_q <= status_cnt_n;
				end
			endcase
	// Trace: design.sv:19517:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:19518:5
		if (~rst_ni)
			// Trace: design.sv:19519:7
			mem_q <= 1'sb0;
		else if (!gate_clock)
			// Trace: design.sv:19521:7
			mem_q <= mem_n;
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_wrapper (
	clk_i,
	rst_ni,
	pulp_clock_en_i,
	scan_cg_en_i,
	boot_addr_i,
	mtvec_addr_i,
	dm_halt_addr_i,
	hart_id_i,
	dm_exception_addr_i,
	instr_req_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_addr_o,
	instr_rdata_i,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_we_o,
	data_be_o,
	data_addr_o,
	data_wdata_o,
	data_rdata_i,
	irq_i,
	irq_ack_o,
	irq_id_o,
	debug_req_i,
	debug_havereset_o,
	debug_running_o,
	debug_halted_o,
	fetch_enable_i,
	core_sleep_o
);
	// Trace: design.sv:19560:15
	parameter PULP_XPULP = 0;
	// Trace: design.sv:19561:15
	parameter PULP_CLUSTER = 0;
	// Trace: design.sv:19562:15
	parameter FPU = 0;
	// Trace: design.sv:19563:15
	parameter PULP_ZFINX = 0;
	// Trace: design.sv:19564:15
	parameter NUM_MHPMCOUNTERS = 1;
	// Trace: design.sv:19567:5
	input wire clk_i;
	// Trace: design.sv:19568:5
	input wire rst_ni;
	// Trace: design.sv:19570:5
	input wire pulp_clock_en_i;
	// Trace: design.sv:19571:5
	input wire scan_cg_en_i;
	// Trace: design.sv:19574:5
	input wire [31:0] boot_addr_i;
	// Trace: design.sv:19575:5
	input wire [31:0] mtvec_addr_i;
	// Trace: design.sv:19576:5
	input wire [31:0] dm_halt_addr_i;
	// Trace: design.sv:19577:5
	input wire [31:0] hart_id_i;
	// Trace: design.sv:19578:5
	input wire [31:0] dm_exception_addr_i;
	// Trace: design.sv:19581:5
	output wire instr_req_o;
	// Trace: design.sv:19582:5
	input wire instr_gnt_i;
	// Trace: design.sv:19583:5
	input wire instr_rvalid_i;
	// Trace: design.sv:19584:5
	output wire [31:0] instr_addr_o;
	// Trace: design.sv:19585:5
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:19588:5
	output wire data_req_o;
	// Trace: design.sv:19589:5
	input wire data_gnt_i;
	// Trace: design.sv:19590:5
	input wire data_rvalid_i;
	// Trace: design.sv:19591:5
	output wire data_we_o;
	// Trace: design.sv:19592:5
	output wire [3:0] data_be_o;
	// Trace: design.sv:19593:5
	output wire [31:0] data_addr_o;
	// Trace: design.sv:19594:5
	output wire [31:0] data_wdata_o;
	// Trace: design.sv:19595:5
	input wire [31:0] data_rdata_i;
	// Trace: design.sv:19598:5
	input wire [31:0] irq_i;
	// Trace: design.sv:19599:5
	output wire irq_ack_o;
	// Trace: design.sv:19600:5
	output wire [4:0] irq_id_o;
	// Trace: design.sv:19603:5
	input wire debug_req_i;
	// Trace: design.sv:19604:5
	output wire debug_havereset_o;
	// Trace: design.sv:19605:5
	output wire debug_running_o;
	// Trace: design.sv:19606:5
	output wire debug_halted_o;
	// Trace: design.sv:19609:5
	input wire fetch_enable_i;
	// Trace: design.sv:19610:5
	output wire core_sleep_o;
	// Trace: design.sv:19613:3
	// removed import cv32e40p_apu_core_pkg::*;
	// Trace: design.sv:19616:3
	wire apu_req;
	// Trace: design.sv:19617:3
	localparam cv32e40p_apu_core_pkg_APU_NARGS_CPU = 3;
	wire [95:0] apu_operands;
	// Trace: design.sv:19618:3
	localparam cv32e40p_apu_core_pkg_APU_WOP_CPU = 6;
	wire [5:0] apu_op;
	// Trace: design.sv:19619:3
	localparam cv32e40p_apu_core_pkg_APU_NDSFLAGS_CPU = 15;
	wire [14:0] apu_flags;
	// Trace: design.sv:19622:3
	wire apu_gnt;
	// Trace: design.sv:19623:3
	wire apu_rvalid;
	// Trace: design.sv:19624:3
	wire [31:0] apu_rdata;
	// Trace: design.sv:19625:3
	localparam cv32e40p_apu_core_pkg_APU_NUSFLAGS_CPU = 5;
	wire [4:0] apu_rflags;
	// Trace: design.sv:19628:3
	cv32e40p_core #(
		.PULP_XPULP(PULP_XPULP),
		.PULP_CLUSTER(PULP_CLUSTER),
		.FPU(FPU),
		.PULP_ZFINX(PULP_ZFINX),
		.NUM_MHPMCOUNTERS(NUM_MHPMCOUNTERS)
	) core_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.pulp_clock_en_i(pulp_clock_en_i),
		.scan_cg_en_i(scan_cg_en_i),
		.boot_addr_i(boot_addr_i),
		.mtvec_addr_i(mtvec_addr_i),
		.dm_halt_addr_i(dm_halt_addr_i),
		.hart_id_i(hart_id_i),
		.dm_exception_addr_i(dm_exception_addr_i),
		.instr_req_o(instr_req_o),
		.instr_gnt_i(instr_gnt_i),
		.instr_rvalid_i(instr_rvalid_i),
		.instr_addr_o(instr_addr_o),
		.instr_rdata_i(instr_rdata_i),
		.data_req_o(data_req_o),
		.data_gnt_i(data_gnt_i),
		.data_rvalid_i(data_rvalid_i),
		.data_we_o(data_we_o),
		.data_be_o(data_be_o),
		.data_addr_o(data_addr_o),
		.data_wdata_o(data_wdata_o),
		.data_rdata_i(data_rdata_i),
		.apu_req_o(apu_req),
		.apu_gnt_i(apu_gnt),
		.apu_operands_o(apu_operands),
		.apu_op_o(apu_op),
		.apu_flags_o(apu_flags),
		.apu_rvalid_i(apu_rvalid),
		.apu_result_i(apu_rdata),
		.apu_flags_i(apu_rflags),
		.irq_i(irq_i),
		.irq_ack_o(irq_ack_o),
		.irq_id_o(irq_id_o),
		.debug_req_i(debug_req_i),
		.debug_havereset_o(debug_havereset_o),
		.debug_running_o(debug_running_o),
		.debug_halted_o(debug_halted_o),
		.fetch_enable_i(fetch_enable_i),
		.core_sleep_o(core_sleep_o)
	);
	// Trace: design.sv:19684:3
	generate
		if (FPU) begin : fpu_gen
			// Trace: design.sv:19687:7
			cv32e40p_fp_wrapper fp_wrapper_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.apu_req_i(apu_req),
				.apu_gnt_o(apu_gnt),
				.apu_operands_i(apu_operands),
				.apu_op_i(apu_op),
				.apu_flags_i(apu_flags),
				.apu_rvalid_o(apu_rvalid),
				.apu_rdata_o(apu_rdata),
				.apu_rflags_o(apu_rflags)
			);
		end
		else begin : no_fpu_gen
			// Trace: design.sv:19701:7
			assign apu_gnt = 1'sb0;
			// Trace: design.sv:19702:7
			assign apu_rvalid = 1'sb0;
			// Trace: design.sv:19703:7
			assign apu_rdata = 1'sb0;
			// Trace: design.sv:19704:7
			assign apu_rflags = 1'sb0;
		end
	endgenerate
endmodule
module cv32e40p_tb_wrapper (
	clk_i,
	rst_ni,
	pulp_clock_en_i,
	scan_cg_en_i,
	boot_addr_i,
	mtvec_addr_i,
	dm_halt_addr_i,
	hart_id_i,
	dm_exception_addr_i,
	instr_req_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_addr_o,
	instr_rdata_i,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_we_o,
	data_be_o,
	data_addr_o,
	data_wdata_o,
	data_rdata_i,
	irq_i,
	irq_ack_o,
	irq_id_o,
	debug_req_i,
	debug_havereset_o,
	debug_running_o,
	debug_halted_o,
	fetch_enable_i,
	core_sleep_o
);
	// removed import cv32e40p_pkg::*;
	// Trace: design.sv:19746:15
	parameter PULP_XPULP = 0;
	// Trace: design.sv:19747:15
	parameter PULP_CLUSTER = 0;
	// Trace: design.sv:19748:15
	parameter FPU = 0;
	// Trace: design.sv:19749:15
	parameter PULP_ZFINX = 0;
	// Trace: design.sv:19750:15
	parameter NUM_MHPMCOUNTERS = 1;
	// Trace: design.sv:19753:5
	input wire clk_i;
	// Trace: design.sv:19754:5
	input wire rst_ni;
	// Trace: design.sv:19756:5
	input wire pulp_clock_en_i;
	// Trace: design.sv:19757:5
	input wire scan_cg_en_i;
	// Trace: design.sv:19760:5
	input wire [31:0] boot_addr_i;
	// Trace: design.sv:19761:5
	input wire [31:0] mtvec_addr_i;
	// Trace: design.sv:19762:5
	input wire [31:0] dm_halt_addr_i;
	// Trace: design.sv:19763:5
	input wire [31:0] hart_id_i;
	// Trace: design.sv:19764:5
	input wire [31:0] dm_exception_addr_i;
	// Trace: design.sv:19767:5
	output wire instr_req_o;
	// Trace: design.sv:19768:5
	input wire instr_gnt_i;
	// Trace: design.sv:19769:5
	input wire instr_rvalid_i;
	// Trace: design.sv:19770:5
	output wire [31:0] instr_addr_o;
	// Trace: design.sv:19771:5
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:19774:5
	output wire data_req_o;
	// Trace: design.sv:19775:5
	input wire data_gnt_i;
	// Trace: design.sv:19776:5
	input wire data_rvalid_i;
	// Trace: design.sv:19777:5
	output wire data_we_o;
	// Trace: design.sv:19778:5
	output wire [3:0] data_be_o;
	// Trace: design.sv:19779:5
	output wire [31:0] data_addr_o;
	// Trace: design.sv:19780:5
	output wire [31:0] data_wdata_o;
	// Trace: design.sv:19781:5
	input wire [31:0] data_rdata_i;
	// Trace: design.sv:19784:5
	input wire [31:0] irq_i;
	// Trace: design.sv:19785:5
	output wire irq_ack_o;
	// Trace: design.sv:19786:5
	output wire [4:0] irq_id_o;
	// Trace: design.sv:19789:5
	input wire debug_req_i;
	// Trace: design.sv:19790:5
	output wire debug_havereset_o;
	// Trace: design.sv:19791:5
	output wire debug_running_o;
	// Trace: design.sv:19792:5
	output wire debug_halted_o;
	// Trace: design.sv:19795:5
	input wire fetch_enable_i;
	// Trace: design.sv:19796:5
	output wire core_sleep_o;
	// Trace: design.sv:20067:3
	cv32e40p_wrapper #(
		.PULP_XPULP(PULP_XPULP),
		.PULP_CLUSTER(PULP_CLUSTER),
		.FPU(FPU),
		.PULP_ZFINX(PULP_ZFINX),
		.NUM_MHPMCOUNTERS(NUM_MHPMCOUNTERS)
	) cv32e40p_wrapper_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.pulp_clock_en_i(pulp_clock_en_i),
		.scan_cg_en_i(scan_cg_en_i),
		.boot_addr_i(boot_addr_i),
		.mtvec_addr_i(mtvec_addr_i),
		.dm_halt_addr_i(dm_halt_addr_i),
		.hart_id_i(hart_id_i),
		.dm_exception_addr_i(dm_exception_addr_i),
		.instr_req_o(instr_req_o),
		.instr_gnt_i(instr_gnt_i),
		.instr_rvalid_i(instr_rvalid_i),
		.instr_addr_o(instr_addr_o),
		.instr_rdata_i(instr_rdata_i),
		.data_req_o(data_req_o),
		.data_gnt_i(data_gnt_i),
		.data_rvalid_i(data_rvalid_i),
		.data_we_o(data_we_o),
		.data_be_o(data_be_o),
		.data_addr_o(data_addr_o),
		.data_wdata_o(data_wdata_o),
		.data_rdata_i(data_rdata_i),
		.irq_i(irq_i),
		.irq_ack_o(irq_ack_o),
		.irq_id_o(irq_id_o),
		.debug_req_i(debug_req_i),
		.debug_havereset_o(debug_havereset_o),
		.debug_running_o(debug_running_o),
		.debug_halted_o(debug_halted_o),
		.fetch_enable_i(fetch_enable_i),
		.core_sleep_o(core_sleep_o)
	);
endmodule
module cv32e40p_register_file (
	clk,
	rst_n,
	scan_cg_en_i,
	raddr_a_i,
	rdata_a_o,
	raddr_b_i,
	rdata_b_o,
	raddr_c_i,
	rdata_c_o,
	waddr_a_i,
	wdata_a_i,
	we_a_i,
	waddr_b_i,
	wdata_b_i,
	we_b_i
);
	// Trace: design.sv:20145:15
	parameter ADDR_WIDTH = 5;
	// Trace: design.sv:20146:15
	parameter DATA_WIDTH = 32;
	// Trace: design.sv:20147:15
	parameter FPU = 0;
	// Trace: design.sv:20148:15
	parameter PULP_ZFINX = 0;
	// Trace: design.sv:20151:5
	input wire clk;
	// Trace: design.sv:20152:5
	input wire rst_n;
	// Trace: design.sv:20154:5
	input wire scan_cg_en_i;
	// Trace: design.sv:20157:5
	input wire [ADDR_WIDTH - 1:0] raddr_a_i;
	// Trace: design.sv:20158:5
	output wire [DATA_WIDTH - 1:0] rdata_a_o;
	// Trace: design.sv:20161:5
	input wire [ADDR_WIDTH - 1:0] raddr_b_i;
	// Trace: design.sv:20162:5
	output wire [DATA_WIDTH - 1:0] rdata_b_o;
	// Trace: design.sv:20165:5
	input wire [ADDR_WIDTH - 1:0] raddr_c_i;
	// Trace: design.sv:20166:5
	output wire [DATA_WIDTH - 1:0] rdata_c_o;
	// Trace: design.sv:20169:5
	input wire [ADDR_WIDTH - 1:0] waddr_a_i;
	// Trace: design.sv:20170:5
	input wire [DATA_WIDTH - 1:0] wdata_a_i;
	// Trace: design.sv:20171:5
	input wire we_a_i;
	// Trace: design.sv:20174:5
	input wire [ADDR_WIDTH - 1:0] waddr_b_i;
	// Trace: design.sv:20175:5
	input wire [DATA_WIDTH - 1:0] wdata_b_i;
	// Trace: design.sv:20176:5
	input wire we_b_i;
	// Trace: design.sv:20180:3
	localparam NUM_WORDS = 2 ** (ADDR_WIDTH - 1);
	// Trace: design.sv:20182:3
	localparam NUM_FP_WORDS = 2 ** (ADDR_WIDTH - 1);
	// Trace: design.sv:20183:3
	localparam NUM_TOT_WORDS = (FPU ? (PULP_ZFINX ? NUM_WORDS : NUM_WORDS + NUM_FP_WORDS) : NUM_WORDS);
	// Trace: design.sv:20186:3
	reg [(NUM_WORDS * DATA_WIDTH) - 1:0] mem;
	// Trace: design.sv:20189:3
	reg [(NUM_FP_WORDS * DATA_WIDTH) - 1:0] mem_fp;
	// Trace: design.sv:20192:3
	wire [ADDR_WIDTH - 1:0] waddr_a;
	// Trace: design.sv:20193:3
	wire [ADDR_WIDTH - 1:0] waddr_b;
	// Trace: design.sv:20196:3
	wire [NUM_TOT_WORDS - 1:0] we_a_dec;
	// Trace: design.sv:20197:3
	wire [NUM_TOT_WORDS - 1:0] we_b_dec;
	// Trace: design.sv:20203:3
	assign rdata_a_o = (raddr_a_i[5] ? mem_fp[raddr_a_i[4:0] * DATA_WIDTH+:DATA_WIDTH] : mem[raddr_a_i[4:0] * DATA_WIDTH+:DATA_WIDTH]);
	// Trace: design.sv:20204:3
	assign rdata_b_o = (raddr_b_i[5] ? mem_fp[raddr_b_i[4:0] * DATA_WIDTH+:DATA_WIDTH] : mem[raddr_b_i[4:0] * DATA_WIDTH+:DATA_WIDTH]);
	// Trace: design.sv:20205:3
	assign rdata_c_o = (raddr_c_i[5] ? mem_fp[raddr_c_i[4:0] * DATA_WIDTH+:DATA_WIDTH] : mem[raddr_c_i[4:0] * DATA_WIDTH+:DATA_WIDTH]);
	// Trace: design.sv:20212:3
	assign waddr_a = waddr_a_i;
	// Trace: design.sv:20213:3
	assign waddr_b = waddr_b_i;
	// Trace: design.sv:20215:3
	genvar _gv_gidx_1;
	// Trace: design.sv:20216:3
	generate
		for (_gv_gidx_1 = 0; _gv_gidx_1 < NUM_TOT_WORDS; _gv_gidx_1 = _gv_gidx_1 + 1) begin : gen_we_decoder
			localparam gidx = _gv_gidx_1;
			// Trace: design.sv:20218:7
			assign we_a_dec[gidx] = (waddr_a == gidx ? we_a_i : 1'b0);
			// Trace: design.sv:20219:7
			assign we_b_dec[gidx] = (waddr_b == gidx ? we_b_i : 1'b0);
		end
	endgenerate
	// Trace: design.sv:20223:3
	genvar _gv_i_5;
	genvar _gv_l_3;
	// Trace: design.sv:20224:3
	// Trace: design.sv:20230:5
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:20231:7
		if (~rst_n)
			// Trace: design.sv:20233:9
			mem[0+:DATA_WIDTH] <= 32'b00000000000000000000000000000000;
		else
			// Trace: design.sv:20236:9
			mem[0+:DATA_WIDTH] <= 32'b00000000000000000000000000000000;
	generate
		for (_gv_i_5 = 1; _gv_i_5 < NUM_WORDS; _gv_i_5 = _gv_i_5 + 1) begin : gen_rf
			localparam i = _gv_i_5;
			// Trace: design.sv:20243:7
			always @(posedge clk or negedge rst_n) begin : register_write_behavioral
				// Trace: design.sv:20244:9
				if (rst_n == 1'b0)
					// Trace: design.sv:20245:11
					mem[i * DATA_WIDTH+:DATA_WIDTH] <= 32'b00000000000000000000000000000000;
				else
					// Trace: design.sv:20247:11
					if (we_b_dec[i] == 1'b1)
						// Trace: design.sv:20247:36
						mem[i * DATA_WIDTH+:DATA_WIDTH] <= wdata_b_i;
					else if (we_a_dec[i] == 1'b1)
						// Trace: design.sv:20248:41
						mem[i * DATA_WIDTH+:DATA_WIDTH] <= wdata_a_i;
			end
		end
		if ((FPU == 1) && (PULP_ZFINX == 0)) begin : gen_mem_fp_write
			for (_gv_l_3 = 0; _gv_l_3 < NUM_FP_WORDS; _gv_l_3 = _gv_l_3 + 1) begin : genblk1
				localparam l = _gv_l_3;
				// Trace: design.sv:20257:9
				always @(posedge clk or negedge rst_n) begin : fp_regs
					// Trace: design.sv:20258:11
					if (rst_n == 1'b0)
						// Trace: design.sv:20258:30
						mem_fp[l * DATA_WIDTH+:DATA_WIDTH] <= 1'sb0;
					else if (we_b_dec[l + NUM_WORDS] == 1'b1)
						// Trace: design.sv:20259:51
						mem_fp[l * DATA_WIDTH+:DATA_WIDTH] <= wdata_b_i;
					else if (we_a_dec[l + NUM_WORDS] == 1'b1)
						// Trace: design.sv:20260:51
						mem_fp[l * DATA_WIDTH+:DATA_WIDTH] <= wdata_a_i;
				end
			end
		end
		else begin : gen_no_mem_fp_write
			// Trace: design.sv:20264:7
			wire [NUM_FP_WORDS * DATA_WIDTH:1] sv2v_tmp_E9FFD;
			assign sv2v_tmp_E9FFD = 'b0;
			always @(*) mem_fp = sv2v_tmp_E9FFD;
		end
	endgenerate
endmodule
module xbar_varlat (
	clk_i,
	rst_ni,
	rr_i,
	req_i,
	add_i,
	wdata_i,
	gnt_o,
	vld_o,
	rdata_o,
	gnt_i,
	req_o,
	vld_i,
	wdata_o,
	rdata_i
);
	// Trace: design.sv:20286:13
	parameter [31:0] AggregateGnt = 1;
	// Trace: design.sv:20287:13
	parameter [31:0] NumIn = 4;
	// Trace: design.sv:20288:13
	parameter [31:0] NumOut = 4;
	// Trace: design.sv:20289:13
	parameter [31:0] ReqDataWidth = 32;
	// Trace: design.sv:20290:13
	parameter [31:0] RespDataWidth = 32;
	// Trace: design.sv:20291:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: design.sv:20292:13
	parameter [31:0] LogNumOut = (NumOut > 1 ? $clog2(NumOut) : 1);
	// Trace: design.sv:20293:13
	parameter [31:0] LogNumIn = (NumIn > 1 ? $clog2(NumIn) : 1);
	// Trace: design.sv:20295:3
	input wire clk_i;
	// Trace: design.sv:20296:3
	input wire rst_ni;
	// Trace: design.sv:20298:3
	input wire [(NumOut * LogNumIn) - 1:0] rr_i;
	// Trace: design.sv:20300:3
	input wire [NumIn - 1:0] req_i;
	// Trace: design.sv:20301:3
	input wire [(NumIn * LogNumOut) - 1:0] add_i;
	// Trace: design.sv:20302:3
	input wire [(NumIn * ReqDataWidth) - 1:0] wdata_i;
	// Trace: design.sv:20303:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: design.sv:20304:3
	output wire [NumIn - 1:0] vld_o;
	// Trace: design.sv:20305:3
	output wire [(NumIn * RespDataWidth) - 1:0] rdata_o;
	// Trace: design.sv:20307:3
	input wire [NumOut - 1:0] gnt_i;
	// Trace: design.sv:20308:3
	output wire [NumOut - 1:0] req_o;
	// Trace: design.sv:20309:3
	input wire [NumOut - 1:0] vld_i;
	// Trace: design.sv:20311:3
	output wire [(NumOut * ReqDataWidth) - 1:0] wdata_o;
	// Trace: design.sv:20313:3
	input wire [(NumOut * RespDataWidth) - 1:0] rdata_i;
	// Trace: design.sv:20334:1
	wire [((NumOut * NumIn) * ReqDataWidth) - 1:0] sl_data;
	// Trace: design.sv:20335:1
	wire [((NumIn * NumOut) * ReqDataWidth) - 1:0] ma_data;
	// Trace: design.sv:20336:1
	wire [(NumOut * NumIn) - 1:0] sl_gnt;
	wire [(NumOut * NumIn) - 1:0] sl_req;
	// Trace: design.sv:20337:1
	wire [(NumIn * NumOut) - 1:0] ma_gnt;
	wire [(NumIn * NumOut) - 1:0] ma_req;
	// Trace: design.sv:20342:1
	genvar _gv_j_4;
	generate
		for (_gv_j_4 = 0; $unsigned(_gv_j_4) < NumIn; _gv_j_4 = _gv_j_4 + 1) begin : gen_inputs
			localparam j = _gv_j_4;
			// Trace: design.sv:20343:3
			addr_dec_resp_mux_varlat #(
				.AggregateGnt(AggregateGnt),
				.NumOut(NumOut),
				.ReqDataWidth(ReqDataWidth),
				.RespDataWidth(RespDataWidth)
			) i_addr_dec_resp_mux(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(req_i[j]),
				.add_i(add_i[j * LogNumOut+:LogNumOut]),
				.data_i(wdata_i[j * ReqDataWidth+:ReqDataWidth]),
				.gnt_o(gnt_o[j]),
				.vld_o(vld_o[j]),
				.rdata_o(rdata_o[j * RespDataWidth+:RespDataWidth]),
				.req_o(ma_req[j * NumOut+:NumOut]),
				.gnt_i(ma_gnt[j * NumOut+:NumOut]),
				.vld_i(vld_i),
				.data_o(ma_data[ReqDataWidth * (j * NumOut)+:ReqDataWidth * NumOut]),
				.rdata_i(rdata_i)
			);
			genvar _gv_k_4;
			for (_gv_k_4 = 0; $unsigned(_gv_k_4) < NumOut; _gv_k_4 = _gv_k_4 + 1) begin : gen_reshape
				localparam k = _gv_k_4;
				// Trace: design.sv:20366:5
				assign sl_req[(k * NumIn) + j] = ma_req[(j * NumOut) + k];
				// Trace: design.sv:20367:5
				assign ma_gnt[(j * NumOut) + k] = sl_gnt[(k * NumIn) + j];
				// Trace: design.sv:20368:5
				assign sl_data[((k * NumIn) + j) * ReqDataWidth+:ReqDataWidth] = ma_data[((j * NumOut) + k) * ReqDataWidth+:ReqDataWidth];
			end
		end
	endgenerate
	// Trace: design.sv:20375:1
	genvar _gv_k_5;
	generate
		for (_gv_k_5 = 0; $unsigned(_gv_k_5) < NumOut; _gv_k_5 = _gv_k_5 + 1) begin : gen_outputs
			localparam k = _gv_k_5;
			if (NumIn == $unsigned(1)) begin : genblk1
				// Trace: design.sv:20377:5
				assign req_o[k] = sl_req[k * NumIn];
				// Trace: design.sv:20378:5
				assign sl_gnt[k * NumIn] = gnt_i[k];
				// Trace: design.sv:20379:5
				assign wdata_o[k * ReqDataWidth+:ReqDataWidth] = sl_data[(k * NumIn) * ReqDataWidth+:ReqDataWidth];
			end
			else begin : gen_rr_arb_tree
				// Trace: design.sv:20381:5
				rr_arb_tree #(
					.NumIn(NumIn),
					.DataWidth(ReqDataWidth),
					.ExtPrio(ExtPrio)
				) i_rr_arb_tree(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.flush_i(1'b0),
					.rr_i(rr_i[k * LogNumIn+:LogNumIn]),
					.req_i(sl_req[k * NumIn+:NumIn]),
					.gnt_o(sl_gnt[k * NumIn+:NumIn]),
					.data_i(sl_data[ReqDataWidth * (k * NumIn)+:ReqDataWidth * NumIn]),
					.gnt_i(gnt_i[k]),
					.req_o(req_o[k]),
					.data_o(wdata_o[k * ReqDataWidth+:ReqDataWidth]),
					.idx_o()
				);
			end
		end
	endgenerate
endmodule
module addr_dec_resp_mux_varlat (
	clk_i,
	rst_ni,
	req_i,
	add_i,
	data_i,
	gnt_o,
	vld_o,
	rdata_o,
	req_o,
	gnt_i,
	vld_i,
	data_o,
	rdata_i
);
	reg _sv2v_0;
	// Trace: design.sv:20432:15
	parameter [31:0] AggregateGnt = 1;
	// Trace: design.sv:20433:15
	parameter [31:0] NumOut = 32;
	// Trace: design.sv:20434:15
	parameter [31:0] ReqDataWidth = 32;
	// Trace: design.sv:20435:15
	parameter [31:0] RespDataWidth = 32;
	// Trace: design.sv:20436:15
	parameter [31:0] LogNumOut = (NumOut > 1 ? $clog2(NumOut) : 1);
	// Trace: design.sv:20438:3
	input wire clk_i;
	// Trace: design.sv:20439:3
	input wire rst_ni;
	// Trace: design.sv:20441:3
	input wire req_i;
	// Trace: design.sv:20442:3
	input wire [LogNumOut - 1:0] add_i;
	// Trace: design.sv:20443:3
	input wire [ReqDataWidth - 1:0] data_i;
	// Trace: design.sv:20444:3
	output wire gnt_o;
	// Trace: design.sv:20445:3
	output wire vld_o;
	// Trace: design.sv:20446:3
	output wire [RespDataWidth - 1:0] rdata_o;
	// Trace: design.sv:20449:3
	output reg [NumOut - 1:0] req_o;
	// Trace: design.sv:20451:3
	input wire [NumOut - 1:0] gnt_i;
	// Trace: design.sv:20452:3
	input wire [NumOut - 1:0] vld_i;
	// Trace: design.sv:20453:3
	output wire [(NumOut * ReqDataWidth) - 1:0] data_o;
	// Trace: design.sv:20454:3
	input wire [(NumOut * RespDataWidth) - 1:0] rdata_i;
	// Trace: design.sv:20457:1
	reg valid_inflight_d;
	reg valid_inflight_q;
	// Trace: design.sv:20462:1
	generate
		if (NumOut == $unsigned(1)) begin : gen_one_output
			// Trace: design.sv:20464:3
			assign data_o[0+:ReqDataWidth] = data_i;
			// Trace: design.sv:20465:3
			assign gnt_o = gnt_i[0];
			// Trace: design.sv:20466:3
			assign rdata_o = rdata_i[0+:RespDataWidth];
			// Trace: design.sv:20467:3
			assign vld_o = vld_i[0] & valid_inflight_q;
			// Trace: design.sv:20470:3
			always @(*) begin : p_addr_dec
				if (_sv2v_0)
					;
				// Trace: design.sv:20471:5
				valid_inflight_d = valid_inflight_q;
				// Trace: design.sv:20472:5
				req_o[0] = 1'sb0;
				// Trace: design.sv:20473:5
				if (~valid_inflight_q) begin
					// Trace: design.sv:20474:7
					req_o[0] = req_i;
					// Trace: design.sv:20475:7
					valid_inflight_d = req_i & gnt_o;
				end
				else begin
					// Trace: design.sv:20478:7
					req_o[0] = 1'sb0;
					// Trace: design.sv:20479:7
					if (vld_o) begin
						// Trace: design.sv:20480:9
						valid_inflight_d = 1'b0;
						// Trace: design.sv:20481:9
						if (req_i) begin
							// Trace: design.sv:20482:11
							req_o[0] = req_i;
							// Trace: design.sv:20483:11
							valid_inflight_d = req_i & gnt_o;
						end
					end
				end
			end
			// Trace: design.sv:20489:3
			always @(posedge clk_i or negedge rst_ni) begin : p_valid_inflight
				// Trace: design.sv:20490:5
				if (!rst_ni)
					// Trace: design.sv:20491:7
					valid_inflight_q <= 1'sb0;
				else
					// Trace: design.sv:20493:7
					valid_inflight_q <= valid_inflight_d;
			end
		end
		else begin : gen_several_outputs
			// Trace: design.sv:20503:3
			always @(*) begin : p_addr_dec
				if (_sv2v_0)
					;
				// Trace: design.sv:20504:5
				req_o = 1'sb0;
				// Trace: design.sv:20505:5
				valid_inflight_d = valid_inflight_q;
				// Trace: design.sv:20506:5
				if (~valid_inflight_q) begin
					// Trace: design.sv:20507:7
					req_o[add_i] = req_i;
					// Trace: design.sv:20508:7
					valid_inflight_d = req_i & gnt_o;
				end
				else begin
					// Trace: design.sv:20511:7
					req_o = 1'sb0;
					// Trace: design.sv:20512:7
					if (vld_o) begin
						// Trace: design.sv:20513:9
						valid_inflight_d = 1'b0;
						// Trace: design.sv:20514:9
						if (req_i) begin
							// Trace: design.sv:20515:11
							req_o[add_i] = req_i;
							// Trace: design.sv:20516:11
							valid_inflight_d = req_i & gnt_o;
						end
					end
				end
			end
			// Trace: design.sv:20523:3
			assign data_o = {NumOut {data_i}};
			// Trace: design.sv:20525:3
			assign gnt_o = (AggregateGnt == 1 ? |gnt_i : gnt_i[add_i]);
			// Trace: design.sv:20527:3
			wire [$clog2(NumOut) - 1:0] bank_sel_d;
			reg [$clog2(NumOut) - 1:0] bank_sel_q;
			// Trace: design.sv:20529:3
			assign rdata_o = rdata_i[bank_sel_q * RespDataWidth+:RespDataWidth];
			// Trace: design.sv:20530:3
			assign vld_o = vld_i[bank_sel_q] & valid_inflight_q;
			// Trace: design.sv:20531:3
			assign bank_sel_d = add_i;
			// Trace: design.sv:20533:3
			always @(posedge clk_i or negedge rst_ni) begin : p_valid_inflight
				// Trace: design.sv:20534:5
				if (!rst_ni) begin
					// Trace: design.sv:20535:7
					valid_inflight_q <= 1'sb0;
					// Trace: design.sv:20536:7
					bank_sel_q <= 1'sb0;
				end
				else begin
					// Trace: design.sv:20538:7
					valid_inflight_q <= valid_inflight_d;
					// Trace: design.sv:20539:7
					if (req_i & gnt_o)
						// Trace: design.sv:20540:9
						bank_sel_q <= bank_sel_d;
				end
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module binary_to_gray (
	A,
	Z
);
	// Trace: design.sv:20576:15
	parameter signed [31:0] N = -1;
	// Trace: design.sv:20578:5
	input wire [N - 1:0] A;
	// Trace: design.sv:20579:5
	output wire [N - 1:0] Z;
	// Trace: design.sv:20581:5
	assign Z = A ^ (A >> 1);
endmodule
// removed package "cb_filter_pkg"
module cc_onehot (
	d_i,
	is_onehot_o
);
	// Trace: design.sv:20627:13
	parameter [31:0] Width = 4;
	// Trace: design.sv:20629:3
	input wire [Width - 1:0] d_i;
	// Trace: design.sv:20630:3
	output wire is_onehot_o;
	// Trace: design.sv:20633:3
	generate
		if (Width == 1) begin : gen_degenerated_onehot
			// Trace: design.sv:20634:5
			assign is_onehot_o = d_i;
		end
		else begin : gen_onehot
			// Trace: design.sv:20636:5
			localparam signed [31:0] LVLS = $clog2(Width) + 1;
			// Trace: design.sv:20638:5
			wire [(LVLS * (2 ** (LVLS - 1))) - 1:0] sum;
			wire [(LVLS * (2 ** (LVLS - 1))) - 1:0] carry;
			// Trace: design.sv:20639:5
			wire [LVLS - 2:0] carry_array;
			// Trace: design.sv:20642:5
			assign sum[0+:2 ** (LVLS - 1)] = $unsigned(d_i);
			genvar _gv_i_6;
			for (_gv_i_6 = 1; _gv_i_6 < LVLS; _gv_i_6 = _gv_i_6 + 1) begin : gen_lvl
				localparam i = _gv_i_6;
				// Trace: design.sv:20647:7
				localparam [31:0] LVLWidth = (2 ** LVLS) / (2 ** i);
				genvar _gv_j_5;
				for (_gv_j_5 = 0; _gv_j_5 < LVLWidth; _gv_j_5 = _gv_j_5 + 2) begin : gen_width
					localparam j = _gv_j_5;
					// Trace: design.sv:20649:9
					assign sum[(i * (2 ** (LVLS - 1))) + (j / 2)] = sum[((i - 1) * (2 ** (LVLS - 1))) + j] ^ sum[((i - 1) * (2 ** (LVLS - 1))) + (j + 1)];
					// Trace: design.sv:20650:9
					assign carry[(i * (2 ** (LVLS - 1))) + (j / 2)] = sum[((i - 1) * (2 ** (LVLS - 1))) + j] & sum[((i - 1) * (2 ** (LVLS - 1))) + (j + 1)];
				end
				// Trace: design.sv:20653:7
				assign carry_array[i - 1] = |carry[(i * (2 ** (LVLS - 1))) + ((LVLWidth / 2) - 1)-:LVLWidth / 2];
			end
			// Trace: design.sv:20655:5
			assign is_onehot_o = sum[(LVLS - 1) * (2 ** (LVLS - 1))] & ~|carry_array;
		end
	endgenerate
endmodule
// removed package "cf_math_pkg"
module clk_int_div (
	clk_i,
	rst_ni,
	en_i,
	test_mode_en_i,
	div_i,
	div_valid_i,
	div_ready_o,
	clk_o,
	cycl_count_o
);
	reg _sv2v_0;
	// Trace: design.sv:20777:13
	parameter [31:0] DIV_VALUE_WIDTH = 4;
	// Trace: design.sv:20779:13
	parameter [31:0] DEFAULT_DIV_VALUE = 0;
	// Trace: design.sv:20781:13
	parameter [0:0] ENABLE_CLOCK_IN_RESET = 1'b0;
	// Trace: design.sv:20783:3
	input wire clk_i;
	// Trace: design.sv:20784:3
	input wire rst_ni;
	// Trace: design.sv:20788:3
	input wire en_i;
	// Trace: design.sv:20791:3
	input wire test_mode_en_i;
	// Trace: design.sv:20795:3
	input wire [DIV_VALUE_WIDTH - 1:0] div_i;
	// Trace: design.sv:20799:3
	input wire div_valid_i;
	// Trace: design.sv:20800:3
	output reg div_ready_o;
	// Trace: design.sv:20807:3
	output wire clk_o;
	// Trace: design.sv:20810:3
	output wire [DIV_VALUE_WIDTH - 1:0] cycl_count_o;
	// Trace: design.sv:20813:3
	generate
		if ($clog2(DEFAULT_DIV_VALUE + 1) > DIV_VALUE_WIDTH) begin : gen_elab_error
			// Trace: design.sv:20814:5
			$error("Default divider value %0d is not representable with the configured", "div value width of %0d bits.", DEFAULT_DIV_VALUE, DIV_VALUE_WIDTH);
		end
	endgenerate
	// Trace: design.sv:20819:3
	reg [DIV_VALUE_WIDTH - 1:0] div_d;
	reg [DIV_VALUE_WIDTH - 1:0] div_q;
	// Trace: design.sv:20820:3
	reg toggle_ffs_en;
	// Trace: design.sv:20821:3
	reg t_ff1_d;
	reg t_ff1_q;
	// Trace: design.sv:20822:3
	reg t_ff1_en;
	// Trace: design.sv:20824:3
	reg t_ff2_d;
	reg t_ff2_q;
	// Trace: design.sv:20825:3
	reg t_ff2_en;
	// Trace: design.sv:20827:3
	reg [DIV_VALUE_WIDTH - 1:0] cycle_cntr_d;
	reg [DIV_VALUE_WIDTH - 1:0] cycle_cntr_q;
	// Trace: design.sv:20828:3
	reg cycle_counter_en;
	// Trace: design.sv:20829:3
	reg clk_div_bypass_en_d;
	reg clk_div_bypass_en_q;
	// Trace: design.sv:20830:3
	wire odd_clk;
	// Trace: design.sv:20831:3
	wire even_clk;
	// Trace: design.sv:20832:3
	wire generated_clock;
	// Trace: design.sv:20833:3
	wire ungated_output_clock;
	// Trace: design.sv:20835:3
	reg use_odd_division_d;
	reg use_odd_division_q;
	// Trace: design.sv:20836:3
	reg gate_en_d;
	reg gate_en_q;
	// Trace: design.sv:20837:3
	reg clear_cycle_counter;
	// Trace: design.sv:20838:3
	reg clear_toggle_flops;
	// Trace: design.sv:20840:3
	// removed localparam type clk_gate_state_e
	// Trace: design.sv:20841:3
	reg [1:0] clk_gate_state_d;
	reg [1:0] clk_gate_state_q;
	// Trace: design.sv:20844:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:20845:5
		div_d = div_q;
		// Trace: design.sv:20846:5
		div_ready_o = 1'b0;
		// Trace: design.sv:20847:5
		clk_div_bypass_en_d = clk_div_bypass_en_q;
		// Trace: design.sv:20848:5
		use_odd_division_d = use_odd_division_q;
		// Trace: design.sv:20849:5
		clk_gate_state_d = clk_gate_state_q;
		// Trace: design.sv:20850:5
		cycle_counter_en = 1'b1;
		// Trace: design.sv:20851:5
		clear_cycle_counter = 1'b0;
		// Trace: design.sv:20852:5
		clear_toggle_flops = 1'b0;
		// Trace: design.sv:20853:5
		toggle_ffs_en = 1'b1;
		// Trace: design.sv:20855:5
		gate_en_d = 1'b0;
		// Trace: design.sv:20856:5
		clk_gate_state_d = clk_gate_state_q;
		// Trace: design.sv:20857:5
		case (clk_gate_state_q)
			2'd0: begin
				// Trace: design.sv:20859:9
				gate_en_d = 1'b1;
				// Trace: design.sv:20860:9
				toggle_ffs_en = 1'b1;
				// Trace: design.sv:20861:9
				if (div_valid_i) begin
					begin
						// Trace: design.sv:20862:11
						if (div_i == div_q)
							// Trace: design.sv:20863:13
							div_ready_o = 1'b1;
						else begin
							// Trace: design.sv:20865:13
							clk_gate_state_d = 2'd1;
							// Trace: design.sv:20866:13
							gate_en_d = 1'b0;
						end
					end
				end
				else if (!en_i && (ungated_output_clock == 1'b0)) begin
					// Trace: design.sv:20871:13
					cycle_counter_en = 1'b0;
					// Trace: design.sv:20872:13
					toggle_ffs_en = 1'b0;
				end
			end
			2'd1: begin
				// Trace: design.sv:20877:9
				gate_en_d = 1'b0;
				// Trace: design.sv:20878:9
				toggle_ffs_en = 1'b1;
				// Trace: design.sv:20883:9
				if ((ungated_output_clock == 1'b0) || clk_div_bypass_en_q) begin
					// Trace: design.sv:20888:11
					toggle_ffs_en = 1'b0;
					// Trace: design.sv:20889:11
					div_d = div_i;
					// Trace: design.sv:20890:11
					div_ready_o = 1'b1;
					// Trace: design.sv:20891:11
					clear_cycle_counter = 1'b1;
					// Trace: design.sv:20892:11
					clear_toggle_flops = 1'b1;
					// Trace: design.sv:20893:11
					use_odd_division_d = div_i[0];
					// Trace: design.sv:20894:11
					clk_div_bypass_en_d = (div_i == 0) || (div_i == 1);
					// Trace: design.sv:20895:11
					clk_gate_state_d = 2'd2;
				end
			end
			2'd2: begin
				// Trace: design.sv:20900:9
				gate_en_d = 1'b0;
				// Trace: design.sv:20905:9
				toggle_ffs_en = 1'b0;
				// Trace: design.sv:20906:9
				if (cycle_cntr_q == (div_q - 1))
					// Trace: design.sv:20907:11
					clk_gate_state_d = 2'd0;
			end
			default:
				// Trace: design.sv:20912:9
				clk_gate_state_d = 2'd0;
		endcase
	end
	// Trace: design.sv:20917:3
	localparam [0:0] UseOddDivisionResetValue = DEFAULT_DIV_VALUE[0];
	// Trace: design.sv:20918:3
	localparam [0:0] ClkDivBypassEnResetValue = (DEFAULT_DIV_VALUE < 2 ? 1'b1 : 1'b0);
	// Trace: design.sv:20920:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:20921:5
		if (!rst_ni) begin
			// Trace: design.sv:20922:7
			use_odd_division_q <= UseOddDivisionResetValue;
			// Trace: design.sv:20923:7
			clk_div_bypass_en_q <= ClkDivBypassEnResetValue;
			// Trace: design.sv:20924:7
			div_q <= DEFAULT_DIV_VALUE;
			// Trace: design.sv:20925:7
			clk_gate_state_q <= 2'd0;
			// Trace: design.sv:20926:7
			gate_en_q <= ENABLE_CLOCK_IN_RESET;
		end
		else begin
			// Trace: design.sv:20928:7
			use_odd_division_q <= use_odd_division_d;
			// Trace: design.sv:20929:7
			clk_div_bypass_en_q <= clk_div_bypass_en_d;
			// Trace: design.sv:20930:7
			div_q <= div_d;
			// Trace: design.sv:20931:7
			clk_gate_state_q <= clk_gate_state_d;
			// Trace: design.sv:20932:7
			gate_en_q <= gate_en_d;
		end
	// Trace: design.sv:20939:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:20940:5
		cycle_cntr_d = cycle_cntr_q;
		// Trace: design.sv:20942:5
		if (clear_cycle_counter)
			// Trace: design.sv:20943:7
			cycle_cntr_d = 1'sb0;
		else
			// Trace: design.sv:20945:7
			if (cycle_counter_en) begin
				begin
					// Trace: design.sv:20949:9
					if (clk_div_bypass_en_q || (cycle_cntr_q == (div_q - 1)))
						// Trace: design.sv:20950:11
						cycle_cntr_d = 1'sb0;
					else
						// Trace: design.sv:20952:11
						cycle_cntr_d = cycle_cntr_q + 1;
				end
			end
	end
	// Trace: design.sv:20958:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:20959:5
		if (!rst_ni)
			// Trace: design.sv:20960:7
			cycle_cntr_q <= 1'sb0;
		else
			// Trace: design.sv:20962:7
			cycle_cntr_q <= cycle_cntr_d;
	// Trace: design.sv:20966:3
	assign cycl_count_o = cycle_cntr_q;
	// Trace: design.sv:20979:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:20980:5
		if (!rst_ni)
			// Trace: design.sv:20981:7
			t_ff1_q = 1'sb0;
		else
			// Trace: design.sv:20983:7
			if (t_ff1_en)
				// Trace: design.sv:20984:9
				t_ff1_q = t_ff1_d;
	// Trace: design.sv:20991:3
	always @(negedge clk_i or negedge rst_ni)
		// Trace: design.sv:20992:5
		if (!rst_ni)
			// Trace: design.sv:20993:7
			t_ff2_q = 1'sb0;
		else
			// Trace: design.sv:20995:7
			if (t_ff2_en)
				// Trace: design.sv:20996:9
				t_ff2_q = t_ff2_d;
	// Trace: design.sv:21001:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:21002:5
		if (clear_toggle_flops) begin
			// Trace: design.sv:21003:7
			t_ff1_d = 1'sb0;
			// Trace: design.sv:21004:7
			t_ff2_d = 1'sb0;
		end
		else begin
			// Trace: design.sv:21006:7
			t_ff1_d = (t_ff1_en ? !t_ff1_q : t_ff1_q);
			// Trace: design.sv:21007:7
			t_ff2_d = (t_ff2_en ? !t_ff2_q : t_ff2_q);
		end
	end
	// Trace: design.sv:21014:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:21015:5
		t_ff1_en = 1'b0;
		// Trace: design.sv:21016:5
		t_ff2_en = 1'b0;
		// Trace: design.sv:21017:5
		if (!clk_div_bypass_en_q && toggle_ffs_en) begin
			begin
				// Trace: design.sv:21018:7
				if (use_odd_division_q) begin
					// Trace: design.sv:21019:9
					t_ff1_en = (cycle_cntr_q == 0 ? 1'b1 : 1'b0);
					// Trace: design.sv:21020:9
					t_ff2_en = (cycle_cntr_q == ((div_q + 1) / 2) ? 1'b1 : 1'b0);
				end
				else
					// Trace: design.sv:21022:9
					t_ff1_en = ((cycle_cntr_q == 0) || (cycle_cntr_q == (div_q / 2)) ? 1'b1 : 1'b0);
			end
		end
	end
	// Trace: design.sv:21027:3
	assign even_clk = t_ff1_q;
	// Trace: design.sv:21030:3
	tc_clk_xor2 i_odd_clk_xor(
		.clk0_i(t_ff1_q),
		.clk1_i(t_ff2_q),
		.clk_o(odd_clk)
	);
	// Trace: design.sv:21037:3
	tc_clk_mux2 i_clk_mux(
		.clk0_i(even_clk),
		.clk1_i(odd_clk),
		.clk_sel_i(use_odd_division_q),
		.clk_o(generated_clock)
	);
	// Trace: design.sv:21045:3
	tc_clk_mux2 i_clk_bypass_mux(
		.clk0_i(generated_clock),
		.clk1_i(clk_i),
		.clk_sel_i(clk_div_bypass_en_q || test_mode_en_i),
		.clk_o(ungated_output_clock)
	);
	// Trace: design.sv:21055:3
	tc_clk_gating #(.IS_FUNCTIONAL(1)) i_clk_gate(
		.clk_i(ungated_output_clock),
		.en_i(gate_en_q & en_i),
		.test_en_i(test_mode_en_i),
		.clk_o(clk_o)
	);
	initial _sv2v_0 = 0;
endmodule
module delta_counter (
	clk_i,
	rst_ni,
	clear_i,
	en_i,
	load_i,
	down_i,
	delta_i,
	d_i,
	q_o,
	overflow_o
);
	reg _sv2v_0;
	// Trace: design.sv:21081:15
	parameter [31:0] WIDTH = 4;
	// Trace: design.sv:21082:15
	parameter [0:0] STICKY_OVERFLOW = 1'b0;
	// Trace: design.sv:21084:5
	input wire clk_i;
	// Trace: design.sv:21085:5
	input wire rst_ni;
	// Trace: design.sv:21086:5
	input wire clear_i;
	// Trace: design.sv:21087:5
	input wire en_i;
	// Trace: design.sv:21088:5
	input wire load_i;
	// Trace: design.sv:21089:5
	input wire down_i;
	// Trace: design.sv:21090:5
	input wire [WIDTH - 1:0] delta_i;
	// Trace: design.sv:21091:5
	input wire [WIDTH - 1:0] d_i;
	// Trace: design.sv:21092:5
	output wire [WIDTH - 1:0] q_o;
	// Trace: design.sv:21093:5
	output wire overflow_o;
	// Trace: design.sv:21095:5
	reg [WIDTH:0] counter_q;
	reg [WIDTH:0] counter_d;
	// Trace: design.sv:21096:5
	generate
		if (STICKY_OVERFLOW) begin : gen_sticky_overflow
			// Trace: design.sv:21097:9
			reg overflow_d;
			reg overflow_q;
			// Trace: design.sv:21098:9
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:21098:54
				overflow_q <= (~rst_ni ? 1'b0 : overflow_d);
			// Trace: design.sv:21099:9
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:21100:13
				overflow_d = overflow_q;
				// Trace: design.sv:21101:13
				if (clear_i || load_i)
					// Trace: design.sv:21102:17
					overflow_d = 1'b0;
				else if (!overflow_q && en_i) begin
					begin
						// Trace: design.sv:21104:17
						if (down_i)
							// Trace: design.sv:21105:21
							overflow_d = delta_i > counter_q[WIDTH - 1:0];
						else
							// Trace: design.sv:21107:21
							overflow_d = counter_q[WIDTH - 1:0] > ({WIDTH {1'b1}} - delta_i);
					end
				end
			end
			// Trace: design.sv:21111:9
			assign overflow_o = overflow_q;
		end
		else begin : gen_transient_overflow
			// Trace: design.sv:21114:9
			assign overflow_o = counter_q[WIDTH];
		end
	endgenerate
	// Trace: design.sv:21116:5
	assign q_o = counter_q[WIDTH - 1:0];
	// Trace: design.sv:21118:5
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:21119:9
		counter_d = counter_q;
		// Trace: design.sv:21121:9
		if (clear_i)
			// Trace: design.sv:21122:13
			counter_d = 1'sb0;
		else if (load_i)
			// Trace: design.sv:21124:13
			counter_d = {1'b0, d_i};
		else if (en_i) begin
			begin
				// Trace: design.sv:21126:13
				if (down_i)
					// Trace: design.sv:21127:17
					counter_d = counter_q - delta_i;
				else
					// Trace: design.sv:21129:17
					counter_d = counter_q + delta_i;
			end
		end
	end
	// Trace: design.sv:21134:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21135:9
		if (!rst_ni)
			// Trace: design.sv:21136:12
			counter_q <= 1'sb0;
		else
			// Trace: design.sv:21138:12
			counter_q <= counter_d;
	initial _sv2v_0 = 0;
endmodule
// removed package "ecc_pkg"
module edge_propagator_tx (
	clk_i,
	rstn_i,
	valid_i,
	ack_i,
	valid_o
);
	// Trace: design.sv:21186:5
	input wire clk_i;
	// Trace: design.sv:21187:5
	input wire rstn_i;
	// Trace: design.sv:21188:5
	input wire valid_i;
	// Trace: design.sv:21189:5
	input wire ack_i;
	// Trace: design.sv:21190:5
	output wire valid_o;
	// Trace: design.sv:21193:5
	reg [1:0] sync_a;
	// Trace: design.sv:21195:5
	reg r_input_reg;
	// Trace: design.sv:21196:5
	wire s_input_reg_next;
	// Trace: design.sv:21198:5
	assign s_input_reg_next = valid_i | (r_input_reg & ~sync_a[0]);
	// Trace: design.sv:21200:5
	always @(negedge rstn_i or posedge clk_i)
		// Trace: design.sv:21201:9
		if (~rstn_i) begin
			// Trace: design.sv:21202:13
			r_input_reg <= 1'b0;
			// Trace: design.sv:21203:13
			sync_a <= 2'b00;
		end
		else begin
			// Trace: design.sv:21205:13
			r_input_reg <= s_input_reg_next;
			// Trace: design.sv:21206:13
			sync_a <= {ack_i, sync_a[1]};
		end
	// Trace: design.sv:21210:5
	assign valid_o = r_input_reg;
endmodule
module exp_backoff (
	clk_i,
	rst_ni,
	set_i,
	clr_i,
	is_zero_o
);
	// Trace: design.sv:21237:13
	parameter [31:0] Seed = 'hffff;
	// Trace: design.sv:21239:13
	parameter [31:0] MaxExp = 16;
	// Trace: design.sv:21241:3
	input wire clk_i;
	// Trace: design.sv:21242:3
	input wire rst_ni;
	// Trace: design.sv:21244:3
	input wire set_i;
	// Trace: design.sv:21246:3
	input wire clr_i;
	// Trace: design.sv:21248:3
	output wire is_zero_o;
	// Trace: design.sv:21252:3
	localparam [31:0] WIDTH = 16;
	// Trace: design.sv:21254:3
	wire [15:0] lfsr_d;
	reg [15:0] lfsr_q;
	wire [15:0] cnt_d;
	reg [15:0] cnt_q;
	wire [15:0] mask_d;
	reg [15:0] mask_q;
	// Trace: design.sv:21255:3
	wire lfsr;
	// Trace: design.sv:21261:3
	assign lfsr = ((lfsr_q[0] ^ lfsr_q[2]) ^ lfsr_q[3]) ^ lfsr_q[5];
	// Trace: design.sv:21266:3
	assign lfsr_d = (set_i ? {lfsr, lfsr_q[15:1]} : lfsr_q);
	// Trace: design.sv:21270:3
	assign mask_d = (clr_i ? {16 {1'sb0}} : (set_i ? {{WIDTH - MaxExp {1'b0}}, mask_q[MaxExp - 2:0], 1'b1} : mask_q));
	// Trace: design.sv:21274:3
	assign cnt_d = (clr_i ? {16 {1'sb0}} : (set_i ? mask_q & lfsr_q : (!is_zero_o ? cnt_q - 1'b1 : {16 {1'sb0}})));
	// Trace: design.sv:21278:3
	assign is_zero_o = cnt_q == {16 {1'sb0}};
	// Trace: design.sv:21280:3
	function automatic [15:0] sv2v_cast_9432F;
		input reg [15:0] inp;
		sv2v_cast_9432F = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:21281:5
		if (!rst_ni) begin
			// Trace: design.sv:21282:7
			lfsr_q <= sv2v_cast_9432F(Seed);
			// Trace: design.sv:21283:7
			mask_q <= 1'sb0;
			// Trace: design.sv:21284:7
			cnt_q <= 1'sb0;
		end
		else begin
			// Trace: design.sv:21286:7
			lfsr_q <= lfsr_d;
			// Trace: design.sv:21287:7
			mask_q <= mask_d;
			// Trace: design.sv:21288:7
			cnt_q <= cnt_d;
		end
	end
endmodule
module fifo_v3 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	reg _sv2v_0;
	// Trace: design.sv:21324:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:21325:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:21326:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:21327:20
	// removed localparam type dtype
	// Trace: design.sv:21329:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:21331:5
	input wire clk_i;
	// Trace: design.sv:21332:5
	input wire rst_ni;
	// Trace: design.sv:21333:5
	input wire flush_i;
	// Trace: design.sv:21334:5
	input wire testmode_i;
	// Trace: design.sv:21336:5
	output wire full_o;
	// Trace: design.sv:21337:5
	output wire empty_o;
	// Trace: design.sv:21338:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:21340:5
	input wire [DATA_WIDTH - 1:0] data_i;
	// Trace: design.sv:21341:5
	input wire push_i;
	// Trace: design.sv:21343:5
	output reg [DATA_WIDTH - 1:0] data_o;
	// Trace: design.sv:21344:5
	input wire pop_i;
	// Trace: design.sv:21348:5
	localparam [31:0] FifoDepth = (DEPTH > 0 ? DEPTH : 1);
	// Trace: design.sv:21350:5
	reg gate_clock;
	// Trace: design.sv:21352:5
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	// Trace: design.sv:21355:5
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	// Trace: design.sv:21357:5
	reg [(FifoDepth * DATA_WIDTH) - 1:0] mem_n;
	reg [(FifoDepth * DATA_WIDTH) - 1:0] mem_q;
	// Trace: design.sv:21359:5
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	// Trace: design.sv:21361:5
	generate
		if (DEPTH == 0) begin : gen_pass_through
			// Trace: design.sv:21362:9
			assign empty_o = ~push_i;
			// Trace: design.sv:21363:9
			assign full_o = ~pop_i;
		end
		else begin : gen_fifo
			// Trace: design.sv:21365:9
			assign full_o = status_cnt_q == FifoDepth[ADDR_DEPTH:0];
			// Trace: design.sv:21366:9
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	// Trace: design.sv:21371:5
	always @(*) begin : read_write_comb
		if (_sv2v_0)
			;
		// Trace: design.sv:21373:9
		read_pointer_n = read_pointer_q;
		// Trace: design.sv:21374:9
		write_pointer_n = write_pointer_q;
		// Trace: design.sv:21375:9
		status_cnt_n = status_cnt_q;
		// Trace: design.sv:21376:9
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q * DATA_WIDTH+:DATA_WIDTH]);
		// Trace: design.sv:21377:9
		mem_n = mem_q;
		// Trace: design.sv:21378:9
		gate_clock = 1'b1;
		// Trace: design.sv:21381:9
		if (push_i && ~full_o) begin
			// Trace: design.sv:21383:13
			mem_n[write_pointer_q * DATA_WIDTH+:DATA_WIDTH] = data_i;
			// Trace: design.sv:21385:13
			gate_clock = 1'b0;
			// Trace: design.sv:21387:13
			if (write_pointer_q == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21388:17
				write_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21390:17
				write_pointer_n = write_pointer_q + 1;
			// Trace: design.sv:21392:13
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			// Trace: design.sv:21398:13
			if (read_pointer_n == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21399:17
				read_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21401:17
				read_pointer_n = read_pointer_q + 1;
			// Trace: design.sv:21403:13
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			// Trace: design.sv:21408:13
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			// Trace: design.sv:21412:13
			data_o = data_i;
			// Trace: design.sv:21413:13
			if (pop_i) begin
				// Trace: design.sv:21414:17
				status_cnt_n = status_cnt_q;
				// Trace: design.sv:21415:17
				read_pointer_n = read_pointer_q;
				// Trace: design.sv:21416:17
				write_pointer_n = write_pointer_q;
			end
		end
	end
	// Trace: design.sv:21422:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21423:9
		if (~rst_ni) begin
			// Trace: design.sv:21424:13
			read_pointer_q <= 1'sb0;
			// Trace: design.sv:21425:13
			write_pointer_q <= 1'sb0;
			// Trace: design.sv:21426:13
			status_cnt_q <= 1'sb0;
		end
		else
			// Trace: design.sv:21428:13
			if (flush_i) begin
				// Trace: design.sv:21429:17
				read_pointer_q <= 1'sb0;
				// Trace: design.sv:21430:17
				write_pointer_q <= 1'sb0;
				// Trace: design.sv:21431:17
				status_cnt_q <= 1'sb0;
			end
			else begin
				// Trace: design.sv:21433:17
				read_pointer_q <= read_pointer_n;
				// Trace: design.sv:21434:17
				write_pointer_q <= write_pointer_n;
				// Trace: design.sv:21435:17
				status_cnt_q <= status_cnt_n;
			end
	// Trace: design.sv:21440:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21441:9
		if (~rst_ni)
			// Trace: design.sv:21442:13
			mem_q <= 1'sb0;
		else if (!gate_clock)
			// Trace: design.sv:21444:13
			mem_q <= mem_n;
	initial _sv2v_0 = 0;
endmodule
module fifo_v3_19420_E888C (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	// removed localparam type dtype_dtype_DATA_WIDTH_type
	parameter [31:0] dtype_dtype_DATA_WIDTH = 0;
	reg _sv2v_0;
	// Trace: design.sv:21324:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:21325:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:21326:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:21327:20
	// removed localparam type dtype
	// Trace: design.sv:21329:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:21331:5
	input wire clk_i;
	// Trace: design.sv:21332:5
	input wire rst_ni;
	// Trace: design.sv:21333:5
	input wire flush_i;
	// Trace: design.sv:21334:5
	input wire testmode_i;
	// Trace: design.sv:21336:5
	output wire full_o;
	// Trace: design.sv:21337:5
	output wire empty_o;
	// Trace: design.sv:21338:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:21340:5
	input wire [dtype_dtype_DATA_WIDTH - 1:0] data_i;
	// Trace: design.sv:21341:5
	input wire push_i;
	// Trace: design.sv:21343:5
	output reg [dtype_dtype_DATA_WIDTH - 1:0] data_o;
	// Trace: design.sv:21344:5
	input wire pop_i;
	// Trace: design.sv:21348:5
	localparam [31:0] FifoDepth = (DEPTH > 0 ? DEPTH : 1);
	// Trace: design.sv:21350:5
	reg gate_clock;
	// Trace: design.sv:21352:5
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	// Trace: design.sv:21355:5
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	// Trace: design.sv:21357:5
	reg [(FifoDepth * dtype_dtype_DATA_WIDTH) - 1:0] mem_n;
	reg [(FifoDepth * dtype_dtype_DATA_WIDTH) - 1:0] mem_q;
	// Trace: design.sv:21359:5
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	// Trace: design.sv:21361:5
	generate
		if (DEPTH == 0) begin : gen_pass_through
			// Trace: design.sv:21362:9
			assign empty_o = ~push_i;
			// Trace: design.sv:21363:9
			assign full_o = ~pop_i;
		end
		else begin : gen_fifo
			// Trace: design.sv:21365:9
			assign full_o = status_cnt_q == FifoDepth[ADDR_DEPTH:0];
			// Trace: design.sv:21366:9
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	// Trace: design.sv:21371:5
	always @(*) begin : read_write_comb
		if (_sv2v_0)
			;
		// Trace: design.sv:21373:9
		read_pointer_n = read_pointer_q;
		// Trace: design.sv:21374:9
		write_pointer_n = write_pointer_q;
		// Trace: design.sv:21375:9
		status_cnt_n = status_cnt_q;
		// Trace: design.sv:21376:9
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q * dtype_dtype_DATA_WIDTH+:dtype_dtype_DATA_WIDTH]);
		// Trace: design.sv:21377:9
		mem_n = mem_q;
		// Trace: design.sv:21378:9
		gate_clock = 1'b1;
		// Trace: design.sv:21381:9
		if (push_i && ~full_o) begin
			// Trace: design.sv:21383:13
			mem_n[write_pointer_q * dtype_dtype_DATA_WIDTH+:dtype_dtype_DATA_WIDTH] = data_i;
			// Trace: design.sv:21385:13
			gate_clock = 1'b0;
			// Trace: design.sv:21387:13
			if (write_pointer_q == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21388:17
				write_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21390:17
				write_pointer_n = write_pointer_q + 1;
			// Trace: design.sv:21392:13
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			// Trace: design.sv:21398:13
			if (read_pointer_n == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21399:17
				read_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21401:17
				read_pointer_n = read_pointer_q + 1;
			// Trace: design.sv:21403:13
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			// Trace: design.sv:21408:13
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			// Trace: design.sv:21412:13
			data_o = data_i;
			// Trace: design.sv:21413:13
			if (pop_i) begin
				// Trace: design.sv:21414:17
				status_cnt_n = status_cnt_q;
				// Trace: design.sv:21415:17
				read_pointer_n = read_pointer_q;
				// Trace: design.sv:21416:17
				write_pointer_n = write_pointer_q;
			end
		end
	end
	// Trace: design.sv:21422:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21423:9
		if (~rst_ni) begin
			// Trace: design.sv:21424:13
			read_pointer_q <= 1'sb0;
			// Trace: design.sv:21425:13
			write_pointer_q <= 1'sb0;
			// Trace: design.sv:21426:13
			status_cnt_q <= 1'sb0;
		end
		else
			// Trace: design.sv:21428:13
			if (flush_i) begin
				// Trace: design.sv:21429:17
				read_pointer_q <= 1'sb0;
				// Trace: design.sv:21430:17
				write_pointer_q <= 1'sb0;
				// Trace: design.sv:21431:17
				status_cnt_q <= 1'sb0;
			end
			else begin
				// Trace: design.sv:21433:17
				read_pointer_q <= read_pointer_n;
				// Trace: design.sv:21434:17
				write_pointer_q <= write_pointer_n;
				// Trace: design.sv:21435:17
				status_cnt_q <= status_cnt_n;
			end
	// Trace: design.sv:21440:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21441:9
		if (~rst_ni)
			// Trace: design.sv:21442:13
			mem_q <= 1'sb0;
		else if (!gate_clock)
			// Trace: design.sv:21444:13
			mem_q <= mem_n;
	initial _sv2v_0 = 0;
endmodule
module fifo_v3_463D7_52D08 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	// removed localparam type dtype_T_AddrWidth_type
	// removed localparam type dtype_T_AtopWidth_type
	// removed localparam type dtype_T_DataWidth_type
	// removed localparam type dtype_T_NumBanks_type
	parameter [31:0] dtype_T_AddrWidth = 0;
	parameter [31:0] dtype_T_AtopWidth = 0;
	parameter [31:0] dtype_T_DataWidth = 0;
	parameter [31:0] dtype_T_NumBanks = 0;
	reg _sv2v_0;
	// Trace: design.sv:21324:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:21325:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:21326:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:21327:20
	// removed localparam type dtype
	// Trace: design.sv:21329:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:21331:5
	input wire clk_i;
	// Trace: design.sv:21332:5
	input wire rst_ni;
	// Trace: design.sv:21333:5
	input wire flush_i;
	// Trace: design.sv:21334:5
	input wire testmode_i;
	// Trace: design.sv:21336:5
	output wire full_o;
	// Trace: design.sv:21337:5
	output wire empty_o;
	// Trace: design.sv:21338:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:21340:5
	input wire [(((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0:0] data_i;
	// Trace: design.sv:21341:5
	input wire push_i;
	// Trace: design.sv:21343:5
	output reg [(((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0:0] data_o;
	// Trace: design.sv:21344:5
	input wire pop_i;
	// Trace: design.sv:21348:5
	localparam [31:0] FifoDepth = (DEPTH > 0 ? DEPTH : 1);
	// Trace: design.sv:21350:5
	reg gate_clock;
	// Trace: design.sv:21352:5
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	// Trace: design.sv:21355:5
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	// Trace: design.sv:21357:5
	reg [(((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? (FifoDepth * ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 1)) - 1 : (FifoDepth * (1 - ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0))) + ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) - 1)):(((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? 0 : (((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0)] mem_n;
	reg [(((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? (FifoDepth * ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 1)) - 1 : (FifoDepth * (1 - ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0))) + ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) - 1)):(((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? 0 : (((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0)] mem_q;
	// Trace: design.sv:21359:5
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	// Trace: design.sv:21361:5
	generate
		if (DEPTH == 0) begin : gen_pass_through
			// Trace: design.sv:21362:9
			assign empty_o = ~push_i;
			// Trace: design.sv:21363:9
			assign full_o = ~pop_i;
		end
		else begin : gen_fifo
			// Trace: design.sv:21365:9
			assign full_o = status_cnt_q == FifoDepth[ADDR_DEPTH:0];
			// Trace: design.sv:21366:9
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	// Trace: design.sv:21371:5
	always @(*) begin : read_write_comb
		if (_sv2v_0)
			;
		// Trace: design.sv:21373:9
		read_pointer_n = read_pointer_q;
		// Trace: design.sv:21374:9
		write_pointer_n = write_pointer_q;
		// Trace: design.sv:21375:9
		status_cnt_n = status_cnt_q;
		// Trace: design.sv:21376:9
		data_o = (DEPTH == 0 ? data_i : mem_q[(((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? 0 : (((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) + (read_pointer_q * (((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? (((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 1 : 1 - ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0)))+:(((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? (((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 1 : 1 - ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0))]);
		// Trace: design.sv:21377:9
		mem_n = mem_q;
		// Trace: design.sv:21378:9
		gate_clock = 1'b1;
		// Trace: design.sv:21381:9
		if (push_i && ~full_o) begin
			// Trace: design.sv:21383:13
			mem_n[(((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? 0 : (((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) + (write_pointer_q * (((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? (((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 1 : 1 - ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0)))+:(((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0) >= 0 ? (((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 1 : 1 - ((((dtype_T_AddrWidth + (dtype_T_DataWidth / dtype_T_NumBanks)) + ((dtype_T_DataWidth / dtype_T_NumBanks) / 8)) + dtype_T_AtopWidth) + 0))] = data_i;
			// Trace: design.sv:21385:13
			gate_clock = 1'b0;
			// Trace: design.sv:21387:13
			if (write_pointer_q == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21388:17
				write_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21390:17
				write_pointer_n = write_pointer_q + 1;
			// Trace: design.sv:21392:13
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			// Trace: design.sv:21398:13
			if (read_pointer_n == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21399:17
				read_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21401:17
				read_pointer_n = read_pointer_q + 1;
			// Trace: design.sv:21403:13
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			// Trace: design.sv:21408:13
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			// Trace: design.sv:21412:13
			data_o = data_i;
			// Trace: design.sv:21413:13
			if (pop_i) begin
				// Trace: design.sv:21414:17
				status_cnt_n = status_cnt_q;
				// Trace: design.sv:21415:17
				read_pointer_n = read_pointer_q;
				// Trace: design.sv:21416:17
				write_pointer_n = write_pointer_q;
			end
		end
	end
	// Trace: design.sv:21422:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21423:9
		if (~rst_ni) begin
			// Trace: design.sv:21424:13
			read_pointer_q <= 1'sb0;
			// Trace: design.sv:21425:13
			write_pointer_q <= 1'sb0;
			// Trace: design.sv:21426:13
			status_cnt_q <= 1'sb0;
		end
		else
			// Trace: design.sv:21428:13
			if (flush_i) begin
				// Trace: design.sv:21429:17
				read_pointer_q <= 1'sb0;
				// Trace: design.sv:21430:17
				write_pointer_q <= 1'sb0;
				// Trace: design.sv:21431:17
				status_cnt_q <= 1'sb0;
			end
			else begin
				// Trace: design.sv:21433:17
				read_pointer_q <= read_pointer_n;
				// Trace: design.sv:21434:17
				write_pointer_q <= write_pointer_n;
				// Trace: design.sv:21435:17
				status_cnt_q <= status_cnt_n;
			end
	// Trace: design.sv:21440:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21441:9
		if (~rst_ni)
			// Trace: design.sv:21442:13
			mem_q <= 1'sb0;
		else if (!gate_clock)
			// Trace: design.sv:21444:13
			mem_q <= mem_n;
	initial _sv2v_0 = 0;
endmodule
module fifo_v3_4D453 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	reg _sv2v_0;
	// Trace: design.sv:21324:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:21325:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:21326:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:21327:20
	// removed localparam type dtype
	// Trace: design.sv:21329:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:21331:5
	input wire clk_i;
	// Trace: design.sv:21332:5
	input wire rst_ni;
	// Trace: design.sv:21333:5
	input wire flush_i;
	// Trace: design.sv:21334:5
	input wire testmode_i;
	// Trace: design.sv:21336:5
	output wire full_o;
	// Trace: design.sv:21337:5
	output wire empty_o;
	// Trace: design.sv:21338:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:21340:5
	input wire [31:0] data_i;
	// Trace: design.sv:21341:5
	input wire push_i;
	// Trace: design.sv:21343:5
	output reg [31:0] data_o;
	// Trace: design.sv:21344:5
	input wire pop_i;
	// Trace: design.sv:21348:5
	localparam [31:0] FifoDepth = (DEPTH > 0 ? DEPTH : 1);
	// Trace: design.sv:21350:5
	reg gate_clock;
	// Trace: design.sv:21352:5
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	// Trace: design.sv:21355:5
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	// Trace: design.sv:21357:5
	reg [(FifoDepth * 32) - 1:0] mem_n;
	reg [(FifoDepth * 32) - 1:0] mem_q;
	// Trace: design.sv:21359:5
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	// Trace: design.sv:21361:5
	generate
		if (DEPTH == 0) begin : gen_pass_through
			// Trace: design.sv:21362:9
			assign empty_o = ~push_i;
			// Trace: design.sv:21363:9
			assign full_o = ~pop_i;
		end
		else begin : gen_fifo
			// Trace: design.sv:21365:9
			assign full_o = status_cnt_q == FifoDepth[ADDR_DEPTH:0];
			// Trace: design.sv:21366:9
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	// Trace: design.sv:21371:5
	always @(*) begin : read_write_comb
		if (_sv2v_0)
			;
		// Trace: design.sv:21373:9
		read_pointer_n = read_pointer_q;
		// Trace: design.sv:21374:9
		write_pointer_n = write_pointer_q;
		// Trace: design.sv:21375:9
		status_cnt_n = status_cnt_q;
		// Trace: design.sv:21376:9
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q * 32+:32]);
		// Trace: design.sv:21377:9
		mem_n = mem_q;
		// Trace: design.sv:21378:9
		gate_clock = 1'b1;
		// Trace: design.sv:21381:9
		if (push_i && ~full_o) begin
			// Trace: design.sv:21383:13
			mem_n[write_pointer_q * 32+:32] = data_i;
			// Trace: design.sv:21385:13
			gate_clock = 1'b0;
			// Trace: design.sv:21387:13
			if (write_pointer_q == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21388:17
				write_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21390:17
				write_pointer_n = write_pointer_q + 1;
			// Trace: design.sv:21392:13
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			// Trace: design.sv:21398:13
			if (read_pointer_n == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21399:17
				read_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21401:17
				read_pointer_n = read_pointer_q + 1;
			// Trace: design.sv:21403:13
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			// Trace: design.sv:21408:13
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			// Trace: design.sv:21412:13
			data_o = data_i;
			// Trace: design.sv:21413:13
			if (pop_i) begin
				// Trace: design.sv:21414:17
				status_cnt_n = status_cnt_q;
				// Trace: design.sv:21415:17
				read_pointer_n = read_pointer_q;
				// Trace: design.sv:21416:17
				write_pointer_n = write_pointer_q;
			end
		end
	end
	// Trace: design.sv:21422:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21423:9
		if (~rst_ni) begin
			// Trace: design.sv:21424:13
			read_pointer_q <= 1'sb0;
			// Trace: design.sv:21425:13
			write_pointer_q <= 1'sb0;
			// Trace: design.sv:21426:13
			status_cnt_q <= 1'sb0;
		end
		else
			// Trace: design.sv:21428:13
			if (flush_i) begin
				// Trace: design.sv:21429:17
				read_pointer_q <= 1'sb0;
				// Trace: design.sv:21430:17
				write_pointer_q <= 1'sb0;
				// Trace: design.sv:21431:17
				status_cnt_q <= 1'sb0;
			end
			else begin
				// Trace: design.sv:21433:17
				read_pointer_q <= read_pointer_n;
				// Trace: design.sv:21434:17
				write_pointer_q <= write_pointer_n;
				// Trace: design.sv:21435:17
				status_cnt_q <= status_cnt_n;
			end
	// Trace: design.sv:21440:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21441:9
		if (~rst_ni)
			// Trace: design.sv:21442:13
			mem_q <= 1'sb0;
		else if (!gate_clock)
			// Trace: design.sv:21444:13
			mem_q <= mem_n;
	initial _sv2v_0 = 0;
endmodule
module fifo_v3_78C92 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	reg _sv2v_0;
	// Trace: design.sv:21324:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:21325:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:21326:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:21327:20
	// removed localparam type dtype
	// Trace: design.sv:21329:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:21331:5
	input wire clk_i;
	// Trace: design.sv:21332:5
	input wire rst_ni;
	// Trace: design.sv:21333:5
	input wire flush_i;
	// Trace: design.sv:21334:5
	input wire testmode_i;
	// Trace: design.sv:21336:5
	output wire full_o;
	// Trace: design.sv:21337:5
	output wire empty_o;
	// Trace: design.sv:21338:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:21340:5
	input wire data_i;
	// Trace: design.sv:21341:5
	input wire push_i;
	// Trace: design.sv:21343:5
	output reg data_o;
	// Trace: design.sv:21344:5
	input wire pop_i;
	// Trace: design.sv:21348:5
	localparam [31:0] FifoDepth = (DEPTH > 0 ? DEPTH : 1);
	// Trace: design.sv:21350:5
	reg gate_clock;
	// Trace: design.sv:21352:5
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	// Trace: design.sv:21355:5
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	// Trace: design.sv:21357:5
	reg [FifoDepth - 1:0] mem_n;
	reg [FifoDepth - 1:0] mem_q;
	// Trace: design.sv:21359:5
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	// Trace: design.sv:21361:5
	generate
		if (DEPTH == 0) begin : gen_pass_through
			// Trace: design.sv:21362:9
			assign empty_o = ~push_i;
			// Trace: design.sv:21363:9
			assign full_o = ~pop_i;
		end
		else begin : gen_fifo
			// Trace: design.sv:21365:9
			assign full_o = status_cnt_q == FifoDepth[ADDR_DEPTH:0];
			// Trace: design.sv:21366:9
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	// Trace: design.sv:21371:5
	always @(*) begin : read_write_comb
		if (_sv2v_0)
			;
		// Trace: design.sv:21373:9
		read_pointer_n = read_pointer_q;
		// Trace: design.sv:21374:9
		write_pointer_n = write_pointer_q;
		// Trace: design.sv:21375:9
		status_cnt_n = status_cnt_q;
		// Trace: design.sv:21376:9
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q]);
		// Trace: design.sv:21377:9
		mem_n = mem_q;
		// Trace: design.sv:21378:9
		gate_clock = 1'b1;
		// Trace: design.sv:21381:9
		if (push_i && ~full_o) begin
			// Trace: design.sv:21383:13
			mem_n[write_pointer_q] = data_i;
			// Trace: design.sv:21385:13
			gate_clock = 1'b0;
			// Trace: design.sv:21387:13
			if (write_pointer_q == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21388:17
				write_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21390:17
				write_pointer_n = write_pointer_q + 1;
			// Trace: design.sv:21392:13
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			// Trace: design.sv:21398:13
			if (read_pointer_n == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21399:17
				read_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21401:17
				read_pointer_n = read_pointer_q + 1;
			// Trace: design.sv:21403:13
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			// Trace: design.sv:21408:13
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			// Trace: design.sv:21412:13
			data_o = data_i;
			// Trace: design.sv:21413:13
			if (pop_i) begin
				// Trace: design.sv:21414:17
				status_cnt_n = status_cnt_q;
				// Trace: design.sv:21415:17
				read_pointer_n = read_pointer_q;
				// Trace: design.sv:21416:17
				write_pointer_n = write_pointer_q;
			end
		end
	end
	// Trace: design.sv:21422:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21423:9
		if (~rst_ni) begin
			// Trace: design.sv:21424:13
			read_pointer_q <= 1'sb0;
			// Trace: design.sv:21425:13
			write_pointer_q <= 1'sb0;
			// Trace: design.sv:21426:13
			status_cnt_q <= 1'sb0;
		end
		else
			// Trace: design.sv:21428:13
			if (flush_i) begin
				// Trace: design.sv:21429:17
				read_pointer_q <= 1'sb0;
				// Trace: design.sv:21430:17
				write_pointer_q <= 1'sb0;
				// Trace: design.sv:21431:17
				status_cnt_q <= 1'sb0;
			end
			else begin
				// Trace: design.sv:21433:17
				read_pointer_q <= read_pointer_n;
				// Trace: design.sv:21434:17
				write_pointer_q <= write_pointer_n;
				// Trace: design.sv:21435:17
				status_cnt_q <= status_cnt_n;
			end
	// Trace: design.sv:21440:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21441:9
		if (~rst_ni)
			// Trace: design.sv:21442:13
			mem_q <= 1'sb0;
		else if (!gate_clock)
			// Trace: design.sv:21444:13
			mem_q <= mem_n;
	initial _sv2v_0 = 0;
endmodule
module fifo_v3_DAF99_42EF4 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	// removed localparam type dtype_T_DataWidth_type
	// removed localparam type dtype_T_NumBanks_type
	parameter [31:0] dtype_T_DataWidth = 0;
	parameter [31:0] dtype_T_NumBanks = 0;
	reg _sv2v_0;
	// Trace: design.sv:21324:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:21325:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:21326:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:21327:20
	// removed localparam type dtype
	// Trace: design.sv:21329:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:21331:5
	input wire clk_i;
	// Trace: design.sv:21332:5
	input wire rst_ni;
	// Trace: design.sv:21333:5
	input wire flush_i;
	// Trace: design.sv:21334:5
	input wire testmode_i;
	// Trace: design.sv:21336:5
	output wire full_o;
	// Trace: design.sv:21337:5
	output wire empty_o;
	// Trace: design.sv:21338:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:21340:5
	input wire [(dtype_T_DataWidth / dtype_T_NumBanks) - 1:0] data_i;
	// Trace: design.sv:21341:5
	input wire push_i;
	// Trace: design.sv:21343:5
	output reg [(dtype_T_DataWidth / dtype_T_NumBanks) - 1:0] data_o;
	// Trace: design.sv:21344:5
	input wire pop_i;
	// Trace: design.sv:21348:5
	localparam [31:0] FifoDepth = (DEPTH > 0 ? DEPTH : 1);
	// Trace: design.sv:21350:5
	reg gate_clock;
	// Trace: design.sv:21352:5
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	// Trace: design.sv:21355:5
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	// Trace: design.sv:21357:5
	reg [(FifoDepth * (dtype_T_DataWidth / dtype_T_NumBanks)) - 1:0] mem_n;
	reg [(FifoDepth * (dtype_T_DataWidth / dtype_T_NumBanks)) - 1:0] mem_q;
	// Trace: design.sv:21359:5
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	// Trace: design.sv:21361:5
	generate
		if (DEPTH == 0) begin : gen_pass_through
			// Trace: design.sv:21362:9
			assign empty_o = ~push_i;
			// Trace: design.sv:21363:9
			assign full_o = ~pop_i;
		end
		else begin : gen_fifo
			// Trace: design.sv:21365:9
			assign full_o = status_cnt_q == FifoDepth[ADDR_DEPTH:0];
			// Trace: design.sv:21366:9
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	// Trace: design.sv:21371:5
	always @(*) begin : read_write_comb
		if (_sv2v_0)
			;
		// Trace: design.sv:21373:9
		read_pointer_n = read_pointer_q;
		// Trace: design.sv:21374:9
		write_pointer_n = write_pointer_q;
		// Trace: design.sv:21375:9
		status_cnt_n = status_cnt_q;
		// Trace: design.sv:21376:9
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q * (dtype_T_DataWidth / dtype_T_NumBanks)+:dtype_T_DataWidth / dtype_T_NumBanks]);
		// Trace: design.sv:21377:9
		mem_n = mem_q;
		// Trace: design.sv:21378:9
		gate_clock = 1'b1;
		// Trace: design.sv:21381:9
		if (push_i && ~full_o) begin
			// Trace: design.sv:21383:13
			mem_n[write_pointer_q * (dtype_T_DataWidth / dtype_T_NumBanks)+:dtype_T_DataWidth / dtype_T_NumBanks] = data_i;
			// Trace: design.sv:21385:13
			gate_clock = 1'b0;
			// Trace: design.sv:21387:13
			if (write_pointer_q == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21388:17
				write_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21390:17
				write_pointer_n = write_pointer_q + 1;
			// Trace: design.sv:21392:13
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			// Trace: design.sv:21398:13
			if (read_pointer_n == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				// Trace: design.sv:21399:17
				read_pointer_n = 1'sb0;
			else
				// Trace: design.sv:21401:17
				read_pointer_n = read_pointer_q + 1;
			// Trace: design.sv:21403:13
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			// Trace: design.sv:21408:13
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			// Trace: design.sv:21412:13
			data_o = data_i;
			// Trace: design.sv:21413:13
			if (pop_i) begin
				// Trace: design.sv:21414:17
				status_cnt_n = status_cnt_q;
				// Trace: design.sv:21415:17
				read_pointer_n = read_pointer_q;
				// Trace: design.sv:21416:17
				write_pointer_n = write_pointer_q;
			end
		end
	end
	// Trace: design.sv:21422:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21423:9
		if (~rst_ni) begin
			// Trace: design.sv:21424:13
			read_pointer_q <= 1'sb0;
			// Trace: design.sv:21425:13
			write_pointer_q <= 1'sb0;
			// Trace: design.sv:21426:13
			status_cnt_q <= 1'sb0;
		end
		else
			// Trace: design.sv:21428:13
			if (flush_i) begin
				// Trace: design.sv:21429:17
				read_pointer_q <= 1'sb0;
				// Trace: design.sv:21430:17
				write_pointer_q <= 1'sb0;
				// Trace: design.sv:21431:17
				status_cnt_q <= 1'sb0;
			end
			else begin
				// Trace: design.sv:21433:17
				read_pointer_q <= read_pointer_n;
				// Trace: design.sv:21434:17
				write_pointer_q <= write_pointer_n;
				// Trace: design.sv:21435:17
				status_cnt_q <= status_cnt_n;
			end
	// Trace: design.sv:21440:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:21441:9
		if (~rst_ni)
			// Trace: design.sv:21442:13
			mem_q <= 1'sb0;
		else if (!gate_clock)
			// Trace: design.sv:21444:13
			mem_q <= mem_n;
	initial _sv2v_0 = 0;
endmodule
module gray_to_binary (
	A,
	Z
);
	// Trace: design.sv:21480:15
	parameter signed [31:0] N = -1;
	// Trace: design.sv:21482:5
	input wire [N - 1:0] A;
	// Trace: design.sv:21483:5
	output wire [N - 1:0] Z;
	// Trace: design.sv:21485:5
	genvar _gv_i_7;
	generate
		for (_gv_i_7 = 0; _gv_i_7 < N; _gv_i_7 = _gv_i_7 + 1) begin : genblk1
			localparam i = _gv_i_7;
			// Trace: design.sv:21486:9
			assign Z[i] = ^A[N - 1:i];
		end
	endgenerate
endmodule
module isochronous_4phase_handshake (
	src_clk_i,
	src_rst_ni,
	src_valid_i,
	src_ready_o,
	dst_clk_i,
	dst_rst_ni,
	dst_valid_o,
	dst_ready_i
);
	// Trace: design.sv:21531:3
	input wire src_clk_i;
	// Trace: design.sv:21532:3
	input wire src_rst_ni;
	// Trace: design.sv:21533:3
	input wire src_valid_i;
	// Trace: design.sv:21534:3
	output wire src_ready_o;
	// Trace: design.sv:21535:3
	input wire dst_clk_i;
	// Trace: design.sv:21536:3
	input wire dst_rst_ni;
	// Trace: design.sv:21537:3
	output wire dst_valid_o;
	// Trace: design.sv:21538:3
	input wire dst_ready_i;
	// Trace: design.sv:21541:3
	reg src_req_q;
	reg src_ack_q;
	// Trace: design.sv:21542:3
	reg dst_req_q;
	reg dst_ack_q;
	// Trace: macro expansion of FFL at design.sv:21545:141
	always @(posedge src_clk_i or negedge src_rst_ni)
		// Trace: macro expansion of FFL at design.sv:21545:238
		if (!src_rst_ni)
			// Trace: macro expansion of FFL at design.sv:21545:335
			src_req_q <= 1'b0;
		else
			// Trace: macro expansion of FFL at design.sv:21545:525
			if (src_valid_i && src_ready_o)
				// Trace: macro expansion of FFL at design.sv:21545:622
				src_req_q <= ~src_req_q;
	// Trace: macro expansion of FF at design.sv:21547:102
	always @(posedge src_clk_i or negedge src_rst_ni)
		// Trace: macro expansion of FF at design.sv:21547:190
		if (!src_rst_ni)
			// Trace: macro expansion of FF at design.sv:21547:278
			src_ack_q <= 1'b0;
		else
			// Trace: macro expansion of FF at design.sv:21547:450
			src_ack_q <= dst_ack_q;
	// Trace: design.sv:21549:3
	assign src_ready_o = src_req_q == src_ack_q;
	// Trace: macro expansion of FFL at design.sv:21552:141
	always @(posedge dst_clk_i or negedge dst_rst_ni)
		// Trace: macro expansion of FFL at design.sv:21552:238
		if (!dst_rst_ni)
			// Trace: macro expansion of FFL at design.sv:21552:335
			dst_ack_q <= 1'b0;
		else
			// Trace: macro expansion of FFL at design.sv:21552:525
			if (dst_valid_o && dst_ready_i)
				// Trace: macro expansion of FFL at design.sv:21552:622
				dst_ack_q <= ~dst_ack_q;
	// Trace: macro expansion of FF at design.sv:21554:102
	always @(posedge dst_clk_i or negedge dst_rst_ni)
		// Trace: macro expansion of FF at design.sv:21554:190
		if (!dst_rst_ni)
			// Trace: macro expansion of FF at design.sv:21554:278
			dst_req_q <= 1'b0;
		else
			// Trace: macro expansion of FF at design.sv:21554:450
			dst_req_q <= src_req_q;
	// Trace: design.sv:21556:3
	assign dst_valid_o = dst_req_q != dst_ack_q;
endmodule
module isochronous_spill_register (
	src_clk_i,
	src_rst_ni,
	src_valid_i,
	src_ready_o,
	src_data_i,
	dst_clk_i,
	dst_rst_ni,
	dst_valid_o,
	dst_ready_i,
	dst_data_o
);
	reg _sv2v_0;
	// Trace: design.sv:21610:18
	// removed localparam type T
	// Trace: design.sv:21612:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:21615:3
	input wire src_clk_i;
	// Trace: design.sv:21617:3
	input wire src_rst_ni;
	// Trace: design.sv:21619:3
	input wire src_valid_i;
	// Trace: design.sv:21621:3
	output wire src_ready_o;
	// Trace: design.sv:21623:3
	input wire src_data_i;
	// Trace: design.sv:21625:3
	input wire dst_clk_i;
	// Trace: design.sv:21627:3
	input wire dst_rst_ni;
	// Trace: design.sv:21629:3
	output wire dst_valid_o;
	// Trace: design.sv:21631:3
	input wire dst_ready_i;
	// Trace: design.sv:21633:3
	output wire dst_data_o;
	// Trace: design.sv:21636:3
	generate
		if (Bypass) begin : gen_bypass
			// Trace: design.sv:21637:5
			assign dst_valid_o = src_valid_i;
			// Trace: design.sv:21638:5
			assign src_ready_o = dst_ready_i;
			// Trace: design.sv:21639:5
			assign dst_data_o = src_data_i;
		end
		else begin : gen_isochronous_spill_register
			// Trace: design.sv:21647:5
			reg [1:0] rd_pointer_q;
			reg [1:0] wr_pointer_q;
			// Trace: macro expansion of FFL at design.sv:21649:148
			always @(posedge src_clk_i or negedge src_rst_ni)
				// Trace: macro expansion of FFL at design.sv:21649:245
				if (!src_rst_ni)
					// Trace: macro expansion of FFL at design.sv:21649:342
					wr_pointer_q <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:21649:532
					if (src_valid_i && src_ready_o)
						// Trace: macro expansion of FFL at design.sv:21649:629
						wr_pointer_q <= wr_pointer_q + 1;
			// Trace: macro expansion of FFL at design.sv:21651:148
			always @(posedge dst_clk_i or negedge dst_rst_ni)
				// Trace: macro expansion of FFL at design.sv:21651:245
				if (!dst_rst_ni)
					// Trace: macro expansion of FFL at design.sv:21651:342
					rd_pointer_q <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:21651:532
					if (dst_valid_o && dst_ready_i)
						// Trace: macro expansion of FFL at design.sv:21651:629
						rd_pointer_q <= rd_pointer_q + 1;
			// Trace: design.sv:21653:5
			reg [1:0] mem_d;
			reg [1:0] mem_q;
			// Trace: macro expansion of FFLNR at design.sv:21654:63
			always @(posedge src_clk_i)
				// Trace: macro expansion of FFLNR at design.sv:21654:105
				if (src_valid_i && src_ready_o)
					// Trace: macro expansion of FFLNR at design.sv:21654:147
					mem_q <= mem_d;
			// Trace: design.sv:21655:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:21656:7
				mem_d = mem_q;
				// Trace: design.sv:21657:7
				mem_d[wr_pointer_q[0]] = src_data_i;
			end
			// Trace: design.sv:21660:5
			assign src_ready_o = (rd_pointer_q ^ wr_pointer_q) != 2'b10;
			// Trace: design.sv:21662:5
			assign dst_valid_o = (rd_pointer_q ^ wr_pointer_q) != {2 {1'sb0}};
			// Trace: design.sv:21663:5
			assign dst_data_o = mem_q[rd_pointer_q[0]];
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module lfsr (
	clk_i,
	rst_ni,
	en_i,
	out_o
);
	reg _sv2v_0;
	// Trace: design.sv:21702:13
	parameter [31:0] LfsrWidth = 64;
	// Trace: design.sv:21703:13
	parameter [31:0] OutWidth = 8;
	// Trace: design.sv:21704:13
	parameter [LfsrWidth - 1:0] RstVal = 1'sb1;
	// Trace: design.sv:21707:13
	parameter [31:0] CipherLayers = 0;
	// Trace: design.sv:21708:13
	parameter [0:0] CipherReg = 1'b1;
	// Trace: design.sv:21710:3
	input wire clk_i;
	// Trace: design.sv:21711:3
	input wire rst_ni;
	// Trace: design.sv:21712:3
	input wire en_i;
	// Trace: design.sv:21713:3
	output wire [OutWidth - 1:0] out_o;
	// Trace: design.sv:21719:1
	localparam [4159:256] Masks = 3904'hc000000000000001e0000000000000039000000000000007e00000000000000fa00000000000001fd00000000000003fc000000000000064b0000000000000d8f0000000000001296000000000000249600000000000043570000000000008679000000000001030e00000000000206cd00000000000403fe00000000000807b800000000001004b200000000002006a800000000004004b20000000000800b8700000000010004f3000000000200072d00000000040006ae00000000080009e300000000100005830000000020000c9200000000400005b60000000080000ea600000001000007a30000000200000abf0000000400000842000000080000123e000000100000074e0000002000000ae9000000400000086a0000008000001213000001000000077e000002000000123b0000040000000877000008000000108d0000100000000ae90000200000000e9f00004000000008a6000080000000191e000100000000090e0002000000000fb30004000000000d7d00080000000016a50010000000000b4b00200000000010af0040000000000dde008000000000181a0100000000000b65020000000000102d0400000000000cd508000000000024c11000000000000ef620000000000013634000000000000fcd80000000000019e2;
	// Trace: design.sv:21791:1
	localparam [63:0] Sbox4 = 64'h21748fe3da09b65c;
	// Trace: design.sv:21797:1
	localparam [383:0] Perm = 384'hfef7cffae78ef6d74df2c70ceeb6cbeaa68ae69649e28608de75c7da6586d65545d24504ce34c3ca2482c61441c20400;
	// Trace: design.sv:21807:1
	function automatic [63:0] sbox4_layer;
		// Trace: design.sv:21807:45
		input reg [63:0] in;
		// Trace: design.sv:21808:3
		reg [63:0] out;
		begin
			// Trace: design.sv:21811:3
			out[0+:4] = Sbox4[in[0+:4] * 4+:4];
			// Trace: design.sv:21812:3
			out[4+:4] = Sbox4[in[4+:4] * 4+:4];
			// Trace: design.sv:21813:3
			out[8+:4] = Sbox4[in[8+:4] * 4+:4];
			// Trace: design.sv:21814:3
			out[12+:4] = Sbox4[in[12+:4] * 4+:4];
			// Trace: design.sv:21816:3
			out[16+:4] = Sbox4[in[16+:4] * 4+:4];
			// Trace: design.sv:21817:3
			out[20+:4] = Sbox4[in[20+:4] * 4+:4];
			// Trace: design.sv:21818:3
			out[24+:4] = Sbox4[in[24+:4] * 4+:4];
			// Trace: design.sv:21819:3
			out[28+:4] = Sbox4[in[28+:4] * 4+:4];
			// Trace: design.sv:21821:3
			out[32+:4] = Sbox4[in[32+:4] * 4+:4];
			// Trace: design.sv:21822:3
			out[36+:4] = Sbox4[in[36+:4] * 4+:4];
			// Trace: design.sv:21823:3
			out[40+:4] = Sbox4[in[40+:4] * 4+:4];
			// Trace: design.sv:21824:3
			out[44+:4] = Sbox4[in[44+:4] * 4+:4];
			// Trace: design.sv:21826:3
			out[48+:4] = Sbox4[in[48+:4] * 4+:4];
			// Trace: design.sv:21827:3
			out[52+:4] = Sbox4[in[52+:4] * 4+:4];
			// Trace: design.sv:21828:3
			out[56+:4] = Sbox4[in[56+:4] * 4+:4];
			// Trace: design.sv:21829:3
			out[60+:4] = Sbox4[in[60+:4] * 4+:4];
			// Trace: design.sv:21830:3
			sbox4_layer = out;
		end
	endfunction
	// Trace: design.sv:21833:1
	function automatic [63:0] perm_layer;
		// Trace: design.sv:21833:44
		input reg [63:0] in;
		// Trace: design.sv:21834:3
		reg [63:0] out;
		begin
			// Trace: design.sv:21837:3
			out[Perm[0+:6]] = in[0];
			// Trace: design.sv:21838:3
			out[Perm[6+:6]] = in[1];
			// Trace: design.sv:21839:3
			out[Perm[12+:6]] = in[2];
			// Trace: design.sv:21840:3
			out[Perm[18+:6]] = in[3];
			// Trace: design.sv:21841:3
			out[Perm[24+:6]] = in[4];
			// Trace: design.sv:21842:3
			out[Perm[30+:6]] = in[5];
			// Trace: design.sv:21843:3
			out[Perm[36+:6]] = in[6];
			// Trace: design.sv:21844:3
			out[Perm[42+:6]] = in[7];
			// Trace: design.sv:21845:3
			out[Perm[48+:6]] = in[8];
			// Trace: design.sv:21846:3
			out[Perm[54+:6]] = in[9];
			// Trace: design.sv:21848:3
			out[Perm[60+:6]] = in[10];
			// Trace: design.sv:21849:3
			out[Perm[66+:6]] = in[11];
			// Trace: design.sv:21850:3
			out[Perm[72+:6]] = in[12];
			// Trace: design.sv:21851:3
			out[Perm[78+:6]] = in[13];
			// Trace: design.sv:21852:3
			out[Perm[84+:6]] = in[14];
			// Trace: design.sv:21853:3
			out[Perm[90+:6]] = in[15];
			// Trace: design.sv:21854:3
			out[Perm[96+:6]] = in[16];
			// Trace: design.sv:21855:3
			out[Perm[102+:6]] = in[17];
			// Trace: design.sv:21856:3
			out[Perm[108+:6]] = in[18];
			// Trace: design.sv:21857:3
			out[Perm[114+:6]] = in[19];
			// Trace: design.sv:21859:3
			out[Perm[120+:6]] = in[20];
			// Trace: design.sv:21860:3
			out[Perm[126+:6]] = in[21];
			// Trace: design.sv:21861:3
			out[Perm[132+:6]] = in[22];
			// Trace: design.sv:21862:3
			out[Perm[138+:6]] = in[23];
			// Trace: design.sv:21863:3
			out[Perm[144+:6]] = in[24];
			// Trace: design.sv:21864:3
			out[Perm[150+:6]] = in[25];
			// Trace: design.sv:21865:3
			out[Perm[156+:6]] = in[26];
			// Trace: design.sv:21866:3
			out[Perm[162+:6]] = in[27];
			// Trace: design.sv:21867:3
			out[Perm[168+:6]] = in[28];
			// Trace: design.sv:21868:3
			out[Perm[174+:6]] = in[29];
			// Trace: design.sv:21870:3
			out[Perm[180+:6]] = in[30];
			// Trace: design.sv:21871:3
			out[Perm[186+:6]] = in[31];
			// Trace: design.sv:21872:3
			out[Perm[192+:6]] = in[32];
			// Trace: design.sv:21873:3
			out[Perm[198+:6]] = in[33];
			// Trace: design.sv:21874:3
			out[Perm[204+:6]] = in[34];
			// Trace: design.sv:21875:3
			out[Perm[210+:6]] = in[35];
			// Trace: design.sv:21876:3
			out[Perm[216+:6]] = in[36];
			// Trace: design.sv:21877:3
			out[Perm[222+:6]] = in[37];
			// Trace: design.sv:21878:3
			out[Perm[228+:6]] = in[38];
			// Trace: design.sv:21879:3
			out[Perm[234+:6]] = in[39];
			// Trace: design.sv:21881:3
			out[Perm[240+:6]] = in[40];
			// Trace: design.sv:21882:3
			out[Perm[246+:6]] = in[41];
			// Trace: design.sv:21883:3
			out[Perm[252+:6]] = in[42];
			// Trace: design.sv:21884:3
			out[Perm[258+:6]] = in[43];
			// Trace: design.sv:21885:3
			out[Perm[264+:6]] = in[44];
			// Trace: design.sv:21886:3
			out[Perm[270+:6]] = in[45];
			// Trace: design.sv:21887:3
			out[Perm[276+:6]] = in[46];
			// Trace: design.sv:21888:3
			out[Perm[282+:6]] = in[47];
			// Trace: design.sv:21889:3
			out[Perm[288+:6]] = in[48];
			// Trace: design.sv:21890:3
			out[Perm[294+:6]] = in[49];
			// Trace: design.sv:21892:3
			out[Perm[300+:6]] = in[50];
			// Trace: design.sv:21893:3
			out[Perm[306+:6]] = in[51];
			// Trace: design.sv:21894:3
			out[Perm[312+:6]] = in[52];
			// Trace: design.sv:21895:3
			out[Perm[318+:6]] = in[53];
			// Trace: design.sv:21896:3
			out[Perm[324+:6]] = in[54];
			// Trace: design.sv:21897:3
			out[Perm[330+:6]] = in[55];
			// Trace: design.sv:21898:3
			out[Perm[336+:6]] = in[56];
			// Trace: design.sv:21899:3
			out[Perm[342+:6]] = in[57];
			// Trace: design.sv:21900:3
			out[Perm[348+:6]] = in[58];
			// Trace: design.sv:21901:3
			out[Perm[354+:6]] = in[59];
			// Trace: design.sv:21903:3
			out[Perm[360+:6]] = in[60];
			// Trace: design.sv:21904:3
			out[Perm[366+:6]] = in[61];
			// Trace: design.sv:21905:3
			out[Perm[372+:6]] = in[62];
			// Trace: design.sv:21906:3
			out[Perm[378+:6]] = in[63];
			// Trace: design.sv:21907:3
			perm_layer = out;
		end
	endfunction
	// Trace: design.sv:21914:1
	wire [LfsrWidth - 1:0] lfsr_d;
	reg [LfsrWidth - 1:0] lfsr_q;
	// Trace: design.sv:21915:1
	assign lfsr_d = (en_i ? (lfsr_q >> 1) ^ ({LfsrWidth {lfsr_q[0]}} & Masks[((68 - LfsrWidth) * 64) + (LfsrWidth - 1)-:LfsrWidth]) : lfsr_q);
	// Trace: design.sv:21918:1
	function automatic [LfsrWidth - 1:0] sv2v_cast_AC421;
		input reg [LfsrWidth - 1:0] inp;
		sv2v_cast_AC421 = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:21920:3
		if (!rst_ni)
			// Trace: design.sv:21921:5
			lfsr_q <= sv2v_cast_AC421(RstVal);
		else
			// Trace: design.sv:21923:5
			lfsr_q <= lfsr_d;
	end
	// Trace: design.sv:21931:1
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	generate
		if (CipherLayers > $unsigned(0)) begin : g_cipher_layers
			// Trace: design.sv:21932:3
			reg [63:0] ciph_layer;
			// Trace: design.sv:21933:3
			localparam [31:0] NumRepl = (64 + LfsrWidth) / LfsrWidth;
			// Trace: design.sv:21935:3
			always @(*) begin : p_ciph_layer
				// Trace: design.sv:21936:5
				reg [63:0] tmp;
				if (_sv2v_0)
					;
				// Trace: design.sv:21937:5
				tmp = sv2v_cast_64({NumRepl {lfsr_q}});
				// Trace: design.sv:21938:5
				begin : sv2v_autoblock_1
					// Trace: design.sv:21938:9
					reg [31:0] k;
					// Trace: design.sv:21938:9
					for (k = 0; k < CipherLayers; k = k + 1)
						begin
							// Trace: design.sv:21939:7
							tmp = perm_layer(sbox4_layer(tmp));
						end
				end
				// Trace: design.sv:21941:5
				ciph_layer = tmp;
			end
			if (CipherReg) begin : g_cipher_reg
				// Trace: design.sv:21946:5
				wire [OutWidth - 1:0] out_d;
				reg [OutWidth - 1:0] out_q;
				// Trace: design.sv:21948:5
				assign out_d = (en_i ? ciph_layer[OutWidth - 1:0] : out_q);
				// Trace: design.sv:21949:5
				assign out_o = out_q[OutWidth - 1:0];
				// Trace: design.sv:21951:5
				always @(posedge clk_i or negedge rst_ni) begin : p_regs
					// Trace: design.sv:21952:7
					if (!rst_ni)
						// Trace: design.sv:21953:9
						out_q <= 1'sb0;
					else
						// Trace: design.sv:21955:9
						out_q <= out_d;
				end
			end
			else begin : g_no_out_reg
				// Trace: design.sv:21960:5
				assign out_o = ciph_layer[OutWidth - 1:0];
			end
		end
		else begin : g_no_cipher_layers
			// Trace: design.sv:21965:3
			assign out_o = lfsr_q[OutWidth - 1:0];
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module lfsr_16bit (
	clk_i,
	rst_ni,
	en_i,
	refill_way_oh,
	refill_way_bin
);
	reg _sv2v_0;
	// Trace: design.sv:22015:15
	parameter [15:0] SEED = 8'b00000000;
	// Trace: design.sv:22016:15
	parameter [31:0] WIDTH = 16;
	// Trace: design.sv:22018:5
	input wire clk_i;
	// Trace: design.sv:22019:5
	input wire rst_ni;
	// Trace: design.sv:22020:5
	input wire en_i;
	// Trace: design.sv:22021:5
	output reg [WIDTH - 1:0] refill_way_oh;
	// Trace: design.sv:22022:5
	output reg [$clog2(WIDTH) - 1:0] refill_way_bin;
	// Trace: design.sv:22025:5
	localparam [31:0] LogWidth = $clog2(WIDTH);
	// Trace: design.sv:22027:5
	reg [15:0] shift_d;
	reg [15:0] shift_q;
	// Trace: design.sv:22030:5
	always @(*) begin : sv2v_autoblock_1
		// Trace: design.sv:22032:9
		reg shift_in;
		if (_sv2v_0)
			;
		// Trace: design.sv:22033:9
		shift_in = !(((shift_q[15] ^ shift_q[12]) ^ shift_q[5]) ^ shift_q[1]);
		// Trace: design.sv:22035:9
		shift_d = shift_q;
		// Trace: design.sv:22037:9
		if (en_i)
			// Trace: design.sv:22038:13
			shift_d = {shift_q[14:0], shift_in};
		// Trace: design.sv:22041:9
		refill_way_oh = 'b0;
		// Trace: design.sv:22042:9
		refill_way_oh[shift_q[LogWidth - 1:0]] = 1'b1;
		// Trace: design.sv:22043:9
		refill_way_bin = shift_q;
	end
	// Trace: design.sv:22046:5
	always @(posedge clk_i or negedge rst_ni) begin : proc_
		// Trace: design.sv:22047:9
		if (~rst_ni)
			// Trace: design.sv:22048:13
			shift_q <= SEED;
		else
			// Trace: design.sv:22050:13
			shift_q <= shift_d;
	end
	initial _sv2v_0 = 0;
endmodule
module lfsr_8bit (
	clk_i,
	rst_ni,
	en_i,
	refill_way_oh,
	refill_way_bin
);
	reg _sv2v_0;
	// Trace: design.sv:22081:13
	parameter [7:0] SEED = 8'b00000000;
	// Trace: design.sv:22082:13
	parameter [31:0] WIDTH = 8;
	// Trace: design.sv:22084:3
	input wire clk_i;
	// Trace: design.sv:22085:3
	input wire rst_ni;
	// Trace: design.sv:22086:3
	input wire en_i;
	// Trace: design.sv:22087:3
	output reg [WIDTH - 1:0] refill_way_oh;
	// Trace: design.sv:22088:3
	output reg [$clog2(WIDTH) - 1:0] refill_way_bin;
	// Trace: design.sv:22091:3
	localparam [31:0] LogWidth = $clog2(WIDTH);
	// Trace: design.sv:22093:3
	reg [7:0] shift_d;
	reg [7:0] shift_q;
	// Trace: design.sv:22095:3
	always @(*) begin : sv2v_autoblock_1
		// Trace: design.sv:22097:5
		reg shift_in;
		if (_sv2v_0)
			;
		// Trace: design.sv:22098:5
		shift_in = !(((shift_q[7] ^ shift_q[3]) ^ shift_q[2]) ^ shift_q[1]);
		// Trace: design.sv:22100:5
		shift_d = shift_q;
		// Trace: design.sv:22102:5
		if (en_i)
			// Trace: design.sv:22102:15
			shift_d = {shift_q[6:0], shift_in};
		// Trace: design.sv:22105:5
		refill_way_oh = 'b0;
		// Trace: design.sv:22106:5
		refill_way_oh[shift_q[LogWidth - 1:0]] = 1'b1;
		// Trace: design.sv:22107:5
		refill_way_bin = shift_q;
	end
	// Trace: design.sv:22110:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_
		// Trace: design.sv:22111:5
		if (~rst_ni)
			// Trace: design.sv:22112:7
			shift_q <= SEED;
		else
			// Trace: design.sv:22114:7
			shift_q <= shift_d;
	end
	initial _sv2v_0 = 0;
endmodule
module mv_filter (
	clk_i,
	rst_ni,
	sample_i,
	clear_i,
	d_i,
	q_o
);
	reg _sv2v_0;
	// Trace: design.sv:22140:15
	parameter [31:0] WIDTH = 4;
	// Trace: design.sv:22141:15
	parameter [31:0] THRESHOLD = 10;
	// Trace: design.sv:22143:5
	input wire clk_i;
	// Trace: design.sv:22144:5
	input wire rst_ni;
	// Trace: design.sv:22145:5
	input wire sample_i;
	// Trace: design.sv:22146:5
	input wire clear_i;
	// Trace: design.sv:22147:5
	input wire d_i;
	// Trace: design.sv:22148:5
	output wire q_o;
	// Trace: design.sv:22150:5
	reg [WIDTH - 1:0] counter_q;
	reg [WIDTH - 1:0] counter_d;
	// Trace: design.sv:22151:5
	reg d;
	reg q;
	// Trace: design.sv:22153:5
	assign q_o = q;
	// Trace: design.sv:22155:5
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:22156:9
		counter_d = counter_q;
		// Trace: design.sv:22157:9
		d = q;
		// Trace: design.sv:22159:9
		if (counter_q >= THRESHOLD[WIDTH - 1:0])
			// Trace: design.sv:22160:13
			d = 1'b1;
		else if (sample_i && d_i)
			// Trace: design.sv:22162:13
			counter_d = counter_q + 1;
		if (clear_i) begin
			// Trace: design.sv:22167:13
			counter_d = 1'sb0;
			// Trace: design.sv:22168:13
			d = 1'b0;
		end
	end
	// Trace: design.sv:22172:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:22173:9
		if (~rst_ni) begin
			// Trace: design.sv:22174:13
			counter_q <= 1'sb0;
			// Trace: design.sv:22175:13
			q <= 1'b0;
		end
		else begin
			// Trace: design.sv:22177:13
			counter_q <= counter_d;
			// Trace: design.sv:22178:13
			q <= d;
		end
	initial _sv2v_0 = 0;
endmodule
module onehot_to_bin (
	onehot,
	bin
);
	// Trace: design.sv:22195:15
	parameter [31:0] ONEHOT_WIDTH = 16;
	// Trace: design.sv:22197:15
	parameter [31:0] BIN_WIDTH = (ONEHOT_WIDTH == 1 ? 1 : $clog2(ONEHOT_WIDTH));
	// Trace: design.sv:22199:5
	input wire [ONEHOT_WIDTH - 1:0] onehot;
	// Trace: design.sv:22200:5
	output wire [BIN_WIDTH - 1:0] bin;
	// Trace: design.sv:22203:5
	genvar _gv_j_6;
	generate
		for (_gv_j_6 = 0; _gv_j_6 < BIN_WIDTH; _gv_j_6 = _gv_j_6 + 1) begin : gen_jl
			localparam j = _gv_j_6;
			// Trace: design.sv:22204:9
			wire [ONEHOT_WIDTH - 1:0] tmp_mask;
			genvar _gv_i_8;
			for (_gv_i_8 = 0; _gv_i_8 < ONEHOT_WIDTH; _gv_i_8 = _gv_i_8 + 1) begin : gen_il
				localparam i = _gv_i_8;
				// Trace: design.sv:22206:17
				wire [BIN_WIDTH - 1:0] tmp_i;
				// Trace: design.sv:22207:17
				assign tmp_i = i;
				// Trace: design.sv:22208:17
				assign tmp_mask[i] = tmp_i[j];
			end
			// Trace: design.sv:22210:9
			assign bin[j] = |(tmp_mask & onehot);
		end
	endgenerate
endmodule
module plru_tree (
	clk_i,
	rst_ni,
	used_i,
	plru_o
);
	reg _sv2v_0;
	// Trace: design.sv:22237:13
	parameter [31:0] ENTRIES = 16;
	// Trace: design.sv:22239:3
	input wire clk_i;
	// Trace: design.sv:22240:3
	input wire rst_ni;
	// Trace: design.sv:22241:3
	input wire [ENTRIES - 1:0] used_i;
	// Trace: design.sv:22242:3
	output reg [ENTRIES - 1:0] plru_o;
	// Trace: design.sv:22245:5
	localparam [31:0] LogEntries = $clog2(ENTRIES);
	// Trace: design.sv:22247:5
	reg [(2 * (ENTRIES - 1)) - 1:0] plru_tree_q;
	reg [(2 * (ENTRIES - 1)) - 1:0] plru_tree_d;
	// Trace: design.sv:22249:5
	always @(*) begin : plru_replacement
		if (_sv2v_0)
			;
		// Trace: design.sv:22250:9
		plru_tree_d = plru_tree_q;
		// Trace: design.sv:22274:9
		begin : sv2v_autoblock_1
			// Trace: design.sv:22274:14
			reg [31:0] i;
			// Trace: design.sv:22274:14
			for (i = 0; i < ENTRIES; i = i + 1)
				begin : sv2v_autoblock_2
					// Trace: design.sv:22275:13
					reg [31:0] idx_base;
					reg [31:0] shift;
					reg [31:0] new_index;
					// Trace: design.sv:22277:13
					if (used_i[i])
						// Trace: design.sv:22279:17
						begin : sv2v_autoblock_3
							// Trace: design.sv:22279:22
							reg [31:0] lvl;
							// Trace: design.sv:22279:22
							for (lvl = 0; lvl < LogEntries; lvl = lvl + 1)
								begin
									// Trace: design.sv:22280:19
									idx_base = $unsigned((2 ** lvl) - 1);
									// Trace: design.sv:22282:19
									shift = LogEntries - lvl;
									// Trace: design.sv:22284:19
									new_index = ~((i >> (shift - 1)) & 1);
									// Trace: design.sv:22285:19
									plru_tree_d[idx_base + (i >> shift)] = new_index[0];
								end
						end
				end
		end
		begin : sv2v_autoblock_4
			// Trace: design.sv:22303:14
			reg [31:0] i;
			// Trace: design.sv:22303:14
			for (i = 0; i < ENTRIES; i = i + 1)
				begin : sv2v_autoblock_5
					// Trace: design.sv:22304:13
					reg en;
					// Trace: design.sv:22305:13
					reg [31:0] idx_base;
					reg [31:0] shift;
					reg [31:0] new_index;
					// Trace: design.sv:22306:13
					en = 1'b1;
					// Trace: design.sv:22307:13
					begin : sv2v_autoblock_6
						// Trace: design.sv:22307:18
						reg [31:0] lvl;
						// Trace: design.sv:22307:18
						for (lvl = 0; lvl < LogEntries; lvl = lvl + 1)
							begin
								// Trace: design.sv:22308:17
								idx_base = $unsigned((2 ** lvl) - 1);
								// Trace: design.sv:22310:17
								shift = LogEntries - lvl;
								// Trace: design.sv:22312:17
								new_index = (i >> (shift - 1)) & 1;
								// Trace: design.sv:22313:17
								if (new_index[0])
									// Trace: design.sv:22314:19
									en = en & plru_tree_q[idx_base + (i >> shift)];
								else
									// Trace: design.sv:22316:19
									en = en & ~plru_tree_q[idx_base + (i >> shift)];
							end
					end
					// Trace: design.sv:22319:13
					plru_o[i] = en;
				end
		end
	end
	// Trace: design.sv:22323:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:22324:9
		if (!rst_ni)
			// Trace: design.sv:22325:13
			plru_tree_q <= 1'sb0;
		else
			// Trace: design.sv:22327:13
			plru_tree_q <= plru_tree_d;
	initial _sv2v_0 = 0;
endmodule
module popcount (
	data_i,
	popcount_o
);
	reg _sv2v_0;
	// Trace: design.sv:22359:15
	parameter [31:0] INPUT_WIDTH = 256;
	// Trace: design.sv:22360:16
	localparam [31:0] PopcountWidth = $clog2(INPUT_WIDTH) + 1;
	// Trace: design.sv:22362:5
	input wire [INPUT_WIDTH - 1:0] data_i;
	// Trace: design.sv:22363:5
	output wire [PopcountWidth - 1:0] popcount_o;
	// Trace: design.sv:22366:4
	localparam [31:0] PaddedWidth = 1 << $clog2(INPUT_WIDTH);
	// Trace: design.sv:22368:4
	reg [PaddedWidth - 1:0] padded_input;
	// Trace: design.sv:22369:4
	wire [PopcountWidth - 2:0] left_child_result;
	wire [PopcountWidth - 2:0] right_child_result;
	// Trace: design.sv:22372:4
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:22373:6
		padded_input = 1'sb0;
		// Trace: design.sv:22374:6
		padded_input[INPUT_WIDTH - 1:0] = data_i;
	end
	// Trace: design.sv:22378:4
	generate
		if (INPUT_WIDTH == 1) begin : gen_single_node
			// Trace: design.sv:22379:6
			assign left_child_result = 1'b0;
			// Trace: design.sv:22380:6
			assign right_child_result = padded_input[0];
		end
		else if (INPUT_WIDTH == 2) begin : gen_leaf_node
			// Trace: design.sv:22382:6
			assign left_child_result = padded_input[1];
			// Trace: design.sv:22383:6
			assign right_child_result = padded_input[0];
		end
		else begin : gen_non_leaf_node
			// Trace: design.sv:22385:6
			popcount #(.INPUT_WIDTH(PaddedWidth / 2)) left_child(
				.data_i(padded_input[PaddedWidth - 1:PaddedWidth / 2]),
				.popcount_o(left_child_result)
			);
			// Trace: design.sv:22390:6
			popcount #(.INPUT_WIDTH(PaddedWidth / 2)) right_child(
				.data_i(padded_input[(PaddedWidth / 2) - 1:0]),
				.popcount_o(right_child_result)
			);
		end
	endgenerate
	// Trace: design.sv:22397:4
	assign popcount_o = left_child_result + right_child_result;
	initial _sv2v_0 = 0;
endmodule
module rr_arb_tree (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	req_o,
	gnt_i,
	data_o,
	idx_o
);
	// Trace: design.sv:22448:13
	parameter [31:0] NumIn = 64;
	// Trace: design.sv:22450:13
	parameter [31:0] DataWidth = 32;
	// Trace: design.sv:22452:26
	// removed localparam type DataType
	// Trace: design.sv:22459:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: design.sv:22466:13
	parameter [0:0] AxiVldRdy = 1'b0;
	// Trace: design.sv:22473:13
	parameter [0:0] LockIn = 1'b0;
	// Trace: design.sv:22477:13
	parameter [0:0] FairArb = 1'b1;
	// Trace: design.sv:22480:13
	parameter [31:0] IdxWidth = (NumIn > 32'd1 ? $unsigned($clog2(NumIn)) : 32'd1);
	// Trace: design.sv:22483:26
	// removed localparam type idx_t
	// Trace: design.sv:22486:3
	input wire clk_i;
	// Trace: design.sv:22488:3
	input wire rst_ni;
	// Trace: design.sv:22490:3
	input wire flush_i;
	// Trace: design.sv:22492:3
	input wire [IdxWidth - 1:0] rr_i;
	// Trace: design.sv:22494:3
	input wire [NumIn - 1:0] req_i;
	// Trace: design.sv:22497:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: design.sv:22500:3
	input wire [(NumIn * DataWidth) - 1:0] data_i;
	// Trace: design.sv:22502:3
	output wire req_o;
	// Trace: design.sv:22504:3
	input wire gnt_i;
	// Trace: design.sv:22506:3
	output wire [DataWidth - 1:0] data_o;
	// Trace: design.sv:22508:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:22521:3
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	function automatic [DataWidth - 1:0] sv2v_cast_8536A;
		input reg [DataWidth - 1:0] inp;
		sv2v_cast_8536A = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : gen_pass_through
			// Trace: design.sv:22522:5
			assign req_o = req_i[0];
			// Trace: design.sv:22523:5
			assign gnt_o[0] = gnt_i;
			// Trace: design.sv:22524:5
			assign data_o = data_i[0+:DataWidth];
			// Trace: design.sv:22525:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_arbiter
			// Trace: design.sv:22528:5
			localparam [31:0] NumLevels = $unsigned($clog2(NumIn));
			// Trace: design.sv:22531:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * IdxWidth) - 1 : ((3 - (2 ** NumLevels)) * IdxWidth) + ((((2 ** NumLevels) - 2) * IdxWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * IdxWidth)] index_nodes;
			// Trace: design.sv:22532:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * DataWidth) - 1 : ((3 - (2 ** NumLevels)) * DataWidth) + ((((2 ** NumLevels) - 2) * DataWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * DataWidth)] data_nodes;
			// Trace: design.sv:22533:5
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			// Trace: design.sv:22534:5
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			// Trace: design.sv:22536:5
			reg [IdxWidth - 1:0] rr_q;
			// Trace: design.sv:22537:5
			wire [NumIn - 1:0] req_d;
			// Trace: design.sv:22540:5
			assign req_o = req_nodes[0];
			// Trace: design.sv:22541:5
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * DataWidth+:DataWidth];
			// Trace: design.sv:22542:5
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * IdxWidth+:IdxWidth];
			if (ExtPrio) begin : gen_ext_rr
				// Trace: design.sv:22545:7
				wire [IdxWidth:1] sv2v_tmp_0900B;
				assign sv2v_tmp_0900B = rr_i;
				always @(*) rr_q = sv2v_tmp_0900B;
				// Trace: design.sv:22546:7
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				// Trace: design.sv:22548:7
				wire [IdxWidth - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					// Trace: design.sv:22552:9
					wire lock_d;
					reg lock_q;
					// Trace: design.sv:22553:9
					reg [NumIn - 1:0] req_q;
					// Trace: design.sv:22555:9
					assign lock_d = req_o & ~gnt_i;
					// Trace: design.sv:22556:9
					assign req_d = (lock_q ? req_q : req_i);
					// Trace: design.sv:22558:9
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						// Trace: design.sv:22559:11
						if (!rst_ni)
							// Trace: design.sv:22560:13
							lock_q <= 1'sb0;
						else
							// Trace: design.sv:22562:13
							if (flush_i)
								// Trace: design.sv:22563:15
								lock_q <= 1'sb0;
							else
								// Trace: design.sv:22565:15
								lock_q <= lock_d;
					end
					// Trace: design.sv:22587:9
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						// Trace: design.sv:22588:11
						if (!rst_ni)
							// Trace: design.sv:22589:13
							req_q <= 1'sb0;
						else
							// Trace: design.sv:22591:13
							if (flush_i)
								// Trace: design.sv:22592:15
								req_q <= 1'sb0;
							else
								// Trace: design.sv:22594:15
								req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					// Trace: design.sv:22599:9
					assign req_d = req_i;
				end
				if (FairArb) begin : gen_fair_arb
					// Trace: design.sv:22603:9
					wire [NumIn - 1:0] upper_mask;
					wire [NumIn - 1:0] lower_mask;
					// Trace: design.sv:22604:9
					wire [IdxWidth - 1:0] upper_idx;
					wire [IdxWidth - 1:0] lower_idx;
					wire [IdxWidth - 1:0] next_idx;
					// Trace: design.sv:22605:9
					wire upper_empty;
					wire lower_empty;
					genvar _gv_i_9;
					for (_gv_i_9 = 0; _gv_i_9 < NumIn; _gv_i_9 = _gv_i_9 + 1) begin : gen_mask
						localparam i = _gv_i_9;
						// Trace: design.sv:22608:11
						assign upper_mask[i] = (i > rr_q ? req_d[i] : 1'b0);
						// Trace: design.sv:22609:11
						assign lower_mask[i] = (i <= rr_q ? req_d[i] : 1'b0);
					end
					// Trace: design.sv:22612:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_upper(
						.in_i(upper_mask),
						.cnt_o(upper_idx),
						.empty_o(upper_empty)
					);
					// Trace: design.sv:22621:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_lower(
						.in_i(lower_mask),
						.cnt_o(lower_idx),
						.empty_o()
					);
					// Trace: design.sv:22630:9
					assign next_idx = (upper_empty ? lower_idx : upper_idx);
					// Trace: design.sv:22631:9
					assign rr_d = (gnt_i && req_o ? next_idx : rr_q);
				end
				else begin : gen_unfair_arb
					// Trace: design.sv:22634:9
					assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5FDFE(NumIn - 1) ? {IdxWidth {1'sb0}} : rr_q + 1'b1) : rr_q);
				end
				// Trace: design.sv:22638:7
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					// Trace: design.sv:22639:9
					if (!rst_ni)
						// Trace: design.sv:22640:11
						rr_q <= 1'sb0;
					else
						// Trace: design.sv:22642:11
						if (flush_i)
							// Trace: design.sv:22643:13
							rr_q <= 1'sb0;
						else
							// Trace: design.sv:22645:13
							rr_q <= rr_d;
				end
			end
			// Trace: design.sv:22651:5
			assign gnt_nodes[0] = gnt_i;
			genvar _gv_level_2;
			for (_gv_level_2 = 0; $unsigned(_gv_level_2) < NumLevels; _gv_level_2 = _gv_level_2 + 1) begin : gen_levels
				localparam level = _gv_level_2;
				genvar _gv_l_4;
				for (_gv_l_4 = 0; _gv_l_4 < (2 ** level); _gv_l_4 = _gv_l_4 + 1) begin : gen_level
					localparam l = _gv_l_4;
					// Trace: design.sv:22657:9
					wire sel;
					// Trace: design.sv:22659:9
					localparam [31:0] Idx0 = ((2 ** level) - 1) + l;
					// Trace: design.sv:22660:9
					localparam [31:0] Idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : gen_reduce
							// Trace: design.sv:22666:13
							assign req_nodes[Idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							// Trace: design.sv:22669:13
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							// Trace: design.sv:22671:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(sel);
							// Trace: design.sv:22672:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * DataWidth+:DataWidth] = (sel ? data_i[((l * 2) + 1) * DataWidth+:DataWidth] : data_i[(l * 2) * DataWidth+:DataWidth]);
							// Trace: design.sv:22673:13
							assign gnt_o[l * 2] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							// Trace: design.sv:22674:13
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : gen_first
							// Trace: design.sv:22678:13
							assign req_nodes[Idx0] = req_d[l * 2];
							// Trace: design.sv:22679:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = 1'sb0;
							// Trace: design.sv:22680:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * DataWidth+:DataWidth] = data_i[(l * 2) * DataWidth+:DataWidth];
							// Trace: design.sv:22681:13
							assign gnt_o[l * 2] = gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : gen_out_of_range
							// Trace: design.sv:22685:13
							assign req_nodes[Idx0] = 1'b0;
							// Trace: design.sv:22686:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(1'sb0);
							// Trace: design.sv:22687:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * DataWidth+:DataWidth] = sv2v_cast_8536A(1'sb0);
						end
					end
					else begin : gen_other_levels
						// Trace: design.sv:22692:11
						assign req_nodes[Idx0] = req_nodes[Idx1] | req_nodes[Idx1 + 1];
						// Trace: design.sv:22695:11
						assign sel = ~req_nodes[Idx1] | (req_nodes[Idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						// Trace: design.sv:22697:11
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = (sel ? sv2v_cast_5FDFE({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5FDFE({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						// Trace: design.sv:22701:11
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * DataWidth+:DataWidth] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * DataWidth+:DataWidth] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * DataWidth+:DataWidth]);
						// Trace: design.sv:22702:11
						assign gnt_nodes[Idx1] = gnt_nodes[Idx0] & ~sel;
						// Trace: design.sv:22703:11
						assign gnt_nodes[Idx1 + 1] = gnt_nodes[Idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_0C7DB_08AEF (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	req_o,
	gnt_i,
	data_o,
	idx_o
);
	// removed localparam type DataType_payload_t_DataWidth_type
	parameter [31:0] DataType_payload_t_DataWidth = 0;
	// Trace: design.sv:22448:13
	parameter [31:0] NumIn = 64;
	// Trace: design.sv:22450:13
	parameter [31:0] DataWidth = 32;
	// Trace: design.sv:22452:26
	// removed localparam type DataType
	// Trace: design.sv:22459:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: design.sv:22466:13
	parameter [0:0] AxiVldRdy = 1'b0;
	// Trace: design.sv:22473:13
	parameter [0:0] LockIn = 1'b0;
	// Trace: design.sv:22477:13
	parameter [0:0] FairArb = 1'b1;
	// Trace: design.sv:22480:13
	parameter [31:0] IdxWidth = (NumIn > 32'd1 ? $unsigned($clog2(NumIn)) : 32'd1);
	// Trace: design.sv:22483:26
	// removed localparam type idx_t
	// Trace: design.sv:22486:3
	input wire clk_i;
	// Trace: design.sv:22488:3
	input wire rst_ni;
	// Trace: design.sv:22490:3
	input wire flush_i;
	// Trace: design.sv:22492:3
	input wire [IdxWidth - 1:0] rr_i;
	// Trace: design.sv:22494:3
	input wire [NumIn - 1:0] req_i;
	// Trace: design.sv:22497:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: design.sv:22500:3
	input wire [(NumIn * DataType_payload_t_DataWidth) - 1:0] data_i;
	// Trace: design.sv:22502:3
	output wire req_o;
	// Trace: design.sv:22504:3
	input wire gnt_i;
	// Trace: design.sv:22506:3
	output wire [DataType_payload_t_DataWidth - 1:0] data_o;
	// Trace: design.sv:22508:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:22521:3
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	function automatic [DataType_payload_t_DataWidth - 1:0] sv2v_cast_9BD02;
		input reg [DataType_payload_t_DataWidth - 1:0] inp;
		sv2v_cast_9BD02 = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : gen_pass_through
			// Trace: design.sv:22522:5
			assign req_o = req_i[0];
			// Trace: design.sv:22523:5
			assign gnt_o[0] = gnt_i;
			// Trace: design.sv:22524:5
			assign data_o = data_i[0+:DataType_payload_t_DataWidth];
			// Trace: design.sv:22525:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_arbiter
			// Trace: design.sv:22528:5
			localparam [31:0] NumLevels = $unsigned($clog2(NumIn));
			// Trace: design.sv:22531:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * IdxWidth) - 1 : ((3 - (2 ** NumLevels)) * IdxWidth) + ((((2 ** NumLevels) - 2) * IdxWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * IdxWidth)] index_nodes;
			// Trace: design.sv:22532:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * DataType_payload_t_DataWidth) - 1 : ((3 - (2 ** NumLevels)) * DataType_payload_t_DataWidth) + ((((2 ** NumLevels) - 2) * DataType_payload_t_DataWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * DataType_payload_t_DataWidth)] data_nodes;
			// Trace: design.sv:22533:5
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			// Trace: design.sv:22534:5
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			// Trace: design.sv:22536:5
			reg [IdxWidth - 1:0] rr_q;
			// Trace: design.sv:22537:5
			wire [NumIn - 1:0] req_d;
			// Trace: design.sv:22540:5
			assign req_o = req_nodes[0];
			// Trace: design.sv:22541:5
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth];
			// Trace: design.sv:22542:5
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * IdxWidth+:IdxWidth];
			if (ExtPrio) begin : gen_ext_rr
				// Trace: design.sv:22545:7
				wire [IdxWidth:1] sv2v_tmp_0900B;
				assign sv2v_tmp_0900B = rr_i;
				always @(*) rr_q = sv2v_tmp_0900B;
				// Trace: design.sv:22546:7
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				// Trace: design.sv:22548:7
				wire [IdxWidth - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					// Trace: design.sv:22552:9
					wire lock_d;
					reg lock_q;
					// Trace: design.sv:22553:9
					reg [NumIn - 1:0] req_q;
					// Trace: design.sv:22555:9
					assign lock_d = req_o & ~gnt_i;
					// Trace: design.sv:22556:9
					assign req_d = (lock_q ? req_q : req_i);
					// Trace: design.sv:22558:9
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						// Trace: design.sv:22559:11
						if (!rst_ni)
							// Trace: design.sv:22560:13
							lock_q <= 1'sb0;
						else
							// Trace: design.sv:22562:13
							if (flush_i)
								// Trace: design.sv:22563:15
								lock_q <= 1'sb0;
							else
								// Trace: design.sv:22565:15
								lock_q <= lock_d;
					end
					// Trace: design.sv:22587:9
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						// Trace: design.sv:22588:11
						if (!rst_ni)
							// Trace: design.sv:22589:13
							req_q <= 1'sb0;
						else
							// Trace: design.sv:22591:13
							if (flush_i)
								// Trace: design.sv:22592:15
								req_q <= 1'sb0;
							else
								// Trace: design.sv:22594:15
								req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					// Trace: design.sv:22599:9
					assign req_d = req_i;
				end
				if (FairArb) begin : gen_fair_arb
					// Trace: design.sv:22603:9
					wire [NumIn - 1:0] upper_mask;
					wire [NumIn - 1:0] lower_mask;
					// Trace: design.sv:22604:9
					wire [IdxWidth - 1:0] upper_idx;
					wire [IdxWidth - 1:0] lower_idx;
					wire [IdxWidth - 1:0] next_idx;
					// Trace: design.sv:22605:9
					wire upper_empty;
					wire lower_empty;
					genvar _gv_i_9;
					for (_gv_i_9 = 0; _gv_i_9 < NumIn; _gv_i_9 = _gv_i_9 + 1) begin : gen_mask
						localparam i = _gv_i_9;
						// Trace: design.sv:22608:11
						assign upper_mask[i] = (i > rr_q ? req_d[i] : 1'b0);
						// Trace: design.sv:22609:11
						assign lower_mask[i] = (i <= rr_q ? req_d[i] : 1'b0);
					end
					// Trace: design.sv:22612:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_upper(
						.in_i(upper_mask),
						.cnt_o(upper_idx),
						.empty_o(upper_empty)
					);
					// Trace: design.sv:22621:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_lower(
						.in_i(lower_mask),
						.cnt_o(lower_idx),
						.empty_o()
					);
					// Trace: design.sv:22630:9
					assign next_idx = (upper_empty ? lower_idx : upper_idx);
					// Trace: design.sv:22631:9
					assign rr_d = (gnt_i && req_o ? next_idx : rr_q);
				end
				else begin : gen_unfair_arb
					// Trace: design.sv:22634:9
					assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5FDFE(NumIn - 1) ? {IdxWidth {1'sb0}} : rr_q + 1'b1) : rr_q);
				end
				// Trace: design.sv:22638:7
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					// Trace: design.sv:22639:9
					if (!rst_ni)
						// Trace: design.sv:22640:11
						rr_q <= 1'sb0;
					else
						// Trace: design.sv:22642:11
						if (flush_i)
							// Trace: design.sv:22643:13
							rr_q <= 1'sb0;
						else
							// Trace: design.sv:22645:13
							rr_q <= rr_d;
				end
			end
			// Trace: design.sv:22651:5
			assign gnt_nodes[0] = gnt_i;
			genvar _gv_level_2;
			for (_gv_level_2 = 0; $unsigned(_gv_level_2) < NumLevels; _gv_level_2 = _gv_level_2 + 1) begin : gen_levels
				localparam level = _gv_level_2;
				genvar _gv_l_4;
				for (_gv_l_4 = 0; _gv_l_4 < (2 ** level); _gv_l_4 = _gv_l_4 + 1) begin : gen_level
					localparam l = _gv_l_4;
					// Trace: design.sv:22657:9
					wire sel;
					// Trace: design.sv:22659:9
					localparam [31:0] Idx0 = ((2 ** level) - 1) + l;
					// Trace: design.sv:22660:9
					localparam [31:0] Idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : gen_reduce
							// Trace: design.sv:22666:13
							assign req_nodes[Idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							// Trace: design.sv:22669:13
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							// Trace: design.sv:22671:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(sel);
							// Trace: design.sv:22672:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth] = (sel ? data_i[((l * 2) + 1) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth] : data_i[(l * 2) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth]);
							// Trace: design.sv:22673:13
							assign gnt_o[l * 2] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							// Trace: design.sv:22674:13
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : gen_first
							// Trace: design.sv:22678:13
							assign req_nodes[Idx0] = req_d[l * 2];
							// Trace: design.sv:22679:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = 1'sb0;
							// Trace: design.sv:22680:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth] = data_i[(l * 2) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth];
							// Trace: design.sv:22681:13
							assign gnt_o[l * 2] = gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : gen_out_of_range
							// Trace: design.sv:22685:13
							assign req_nodes[Idx0] = 1'b0;
							// Trace: design.sv:22686:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(1'sb0);
							// Trace: design.sv:22687:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth] = sv2v_cast_9BD02(1'sb0);
						end
					end
					else begin : gen_other_levels
						// Trace: design.sv:22692:11
						assign req_nodes[Idx0] = req_nodes[Idx1] | req_nodes[Idx1 + 1];
						// Trace: design.sv:22695:11
						assign sel = ~req_nodes[Idx1] | (req_nodes[Idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						// Trace: design.sv:22697:11
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = (sel ? sv2v_cast_5FDFE({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5FDFE({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						// Trace: design.sv:22701:11
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * DataType_payload_t_DataWidth+:DataType_payload_t_DataWidth]);
						// Trace: design.sv:22702:11
						assign gnt_nodes[Idx1] = gnt_nodes[Idx0] & ~sel;
						// Trace: design.sv:22703:11
						assign gnt_nodes[Idx1 + 1] = gnt_nodes[Idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_3ECCC_46CA0 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	req_o,
	gnt_i,
	data_o,
	idx_o
);
	// removed localparam type DataType_Width_type
	parameter [31:0] DataType_Width = 0;
	// Trace: design.sv:22448:13
	parameter [31:0] NumIn = 64;
	// Trace: design.sv:22450:13
	parameter [31:0] DataWidth = 32;
	// Trace: design.sv:22452:26
	// removed localparam type DataType
	// Trace: design.sv:22459:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: design.sv:22466:13
	parameter [0:0] AxiVldRdy = 1'b0;
	// Trace: design.sv:22473:13
	parameter [0:0] LockIn = 1'b0;
	// Trace: design.sv:22477:13
	parameter [0:0] FairArb = 1'b1;
	// Trace: design.sv:22480:13
	parameter [31:0] IdxWidth = (NumIn > 32'd1 ? $unsigned($clog2(NumIn)) : 32'd1);
	// Trace: design.sv:22483:26
	// removed localparam type idx_t
	// Trace: design.sv:22486:3
	input wire clk_i;
	// Trace: design.sv:22488:3
	input wire rst_ni;
	// Trace: design.sv:22490:3
	input wire flush_i;
	// Trace: design.sv:22492:3
	input wire [IdxWidth - 1:0] rr_i;
	// Trace: design.sv:22494:3
	input wire [NumIn - 1:0] req_i;
	// Trace: design.sv:22497:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: design.sv:22500:3
	input wire [((DataType_Width + 6) >= 0 ? (NumIn * (DataType_Width + 7)) - 1 : (NumIn * (1 - (DataType_Width + 6))) + (DataType_Width + 5)):((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6)] data_i;
	// Trace: design.sv:22502:3
	output wire req_o;
	// Trace: design.sv:22504:3
	input wire gnt_i;
	// Trace: design.sv:22506:3
	output wire [DataType_Width + 6:0] data_o;
	// Trace: design.sv:22508:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:22521:3
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	function automatic [((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)) - 1:0] sv2v_cast_5FCB8;
		input reg [((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)) - 1:0] inp;
		sv2v_cast_5FCB8 = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : gen_pass_through
			// Trace: design.sv:22522:5
			assign req_o = req_i[0];
			// Trace: design.sv:22523:5
			assign gnt_o[0] = gnt_i;
			// Trace: design.sv:22524:5
			assign data_o = data_i[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + 0+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))];
			// Trace: design.sv:22525:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_arbiter
			// Trace: design.sv:22528:5
			localparam [31:0] NumLevels = $unsigned($clog2(NumIn));
			// Trace: design.sv:22531:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * IdxWidth) - 1 : ((3 - (2 ** NumLevels)) * IdxWidth) + ((((2 ** NumLevels) - 2) * IdxWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * IdxWidth)] index_nodes;
			// Trace: design.sv:22532:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? ((DataType_Width + 6) >= 0 ? (((2 ** NumLevels) - 1) * (DataType_Width + 7)) - 1 : (((2 ** NumLevels) - 1) * (1 - (DataType_Width + 6))) + (DataType_Width + 5)) : ((DataType_Width + 6) >= 0 ? ((3 - (2 ** NumLevels)) * (DataType_Width + 7)) + ((((2 ** NumLevels) - 2) * (DataType_Width + 7)) - 1) : ((3 - (2 ** NumLevels)) * (1 - (DataType_Width + 6))) + (((DataType_Width + 6) + (((2 ** NumLevels) - 2) * (1 - (DataType_Width + 6)))) - 1))):(((2 ** NumLevels) - 2) >= 0 ? ((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) : ((DataType_Width + 6) >= 0 ? ((2 ** NumLevels) - 2) * (DataType_Width + 7) : (DataType_Width + 6) + (((2 ** NumLevels) - 2) * (1 - (DataType_Width + 6)))))] data_nodes;
			// Trace: design.sv:22533:5
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			// Trace: design.sv:22534:5
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			// Trace: design.sv:22536:5
			reg [IdxWidth - 1:0] rr_q;
			// Trace: design.sv:22537:5
			wire [NumIn - 1:0] req_d;
			// Trace: design.sv:22540:5
			assign req_o = req_nodes[0];
			// Trace: design.sv:22541:5
			assign data_o = data_nodes[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))];
			// Trace: design.sv:22542:5
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * IdxWidth+:IdxWidth];
			if (ExtPrio) begin : gen_ext_rr
				// Trace: design.sv:22545:7
				wire [IdxWidth:1] sv2v_tmp_0900B;
				assign sv2v_tmp_0900B = rr_i;
				always @(*) rr_q = sv2v_tmp_0900B;
				// Trace: design.sv:22546:7
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				// Trace: design.sv:22548:7
				wire [IdxWidth - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					// Trace: design.sv:22552:9
					wire lock_d;
					reg lock_q;
					// Trace: design.sv:22553:9
					reg [NumIn - 1:0] req_q;
					// Trace: design.sv:22555:9
					assign lock_d = req_o & ~gnt_i;
					// Trace: design.sv:22556:9
					assign req_d = (lock_q ? req_q : req_i);
					// Trace: design.sv:22558:9
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						// Trace: design.sv:22559:11
						if (!rst_ni)
							// Trace: design.sv:22560:13
							lock_q <= 1'sb0;
						else
							// Trace: design.sv:22562:13
							if (flush_i)
								// Trace: design.sv:22563:15
								lock_q <= 1'sb0;
							else
								// Trace: design.sv:22565:15
								lock_q <= lock_d;
					end
					// Trace: design.sv:22587:9
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						// Trace: design.sv:22588:11
						if (!rst_ni)
							// Trace: design.sv:22589:13
							req_q <= 1'sb0;
						else
							// Trace: design.sv:22591:13
							if (flush_i)
								// Trace: design.sv:22592:15
								req_q <= 1'sb0;
							else
								// Trace: design.sv:22594:15
								req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					// Trace: design.sv:22599:9
					assign req_d = req_i;
				end
				if (FairArb) begin : gen_fair_arb
					// Trace: design.sv:22603:9
					wire [NumIn - 1:0] upper_mask;
					wire [NumIn - 1:0] lower_mask;
					// Trace: design.sv:22604:9
					wire [IdxWidth - 1:0] upper_idx;
					wire [IdxWidth - 1:0] lower_idx;
					wire [IdxWidth - 1:0] next_idx;
					// Trace: design.sv:22605:9
					wire upper_empty;
					wire lower_empty;
					genvar _gv_i_9;
					for (_gv_i_9 = 0; _gv_i_9 < NumIn; _gv_i_9 = _gv_i_9 + 1) begin : gen_mask
						localparam i = _gv_i_9;
						// Trace: design.sv:22608:11
						assign upper_mask[i] = (i > rr_q ? req_d[i] : 1'b0);
						// Trace: design.sv:22609:11
						assign lower_mask[i] = (i <= rr_q ? req_d[i] : 1'b0);
					end
					// Trace: design.sv:22612:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_upper(
						.in_i(upper_mask),
						.cnt_o(upper_idx),
						.empty_o(upper_empty)
					);
					// Trace: design.sv:22621:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_lower(
						.in_i(lower_mask),
						.cnt_o(lower_idx),
						.empty_o()
					);
					// Trace: design.sv:22630:9
					assign next_idx = (upper_empty ? lower_idx : upper_idx);
					// Trace: design.sv:22631:9
					assign rr_d = (gnt_i && req_o ? next_idx : rr_q);
				end
				else begin : gen_unfair_arb
					// Trace: design.sv:22634:9
					assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5FDFE(NumIn - 1) ? {IdxWidth {1'sb0}} : rr_q + 1'b1) : rr_q);
				end
				// Trace: design.sv:22638:7
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					// Trace: design.sv:22639:9
					if (!rst_ni)
						// Trace: design.sv:22640:11
						rr_q <= 1'sb0;
					else
						// Trace: design.sv:22642:11
						if (flush_i)
							// Trace: design.sv:22643:13
							rr_q <= 1'sb0;
						else
							// Trace: design.sv:22645:13
							rr_q <= rr_d;
				end
			end
			// Trace: design.sv:22651:5
			assign gnt_nodes[0] = gnt_i;
			genvar _gv_level_2;
			for (_gv_level_2 = 0; $unsigned(_gv_level_2) < NumLevels; _gv_level_2 = _gv_level_2 + 1) begin : gen_levels
				localparam level = _gv_level_2;
				genvar _gv_l_4;
				for (_gv_l_4 = 0; _gv_l_4 < (2 ** level); _gv_l_4 = _gv_l_4 + 1) begin : gen_level
					localparam l = _gv_l_4;
					// Trace: design.sv:22657:9
					wire sel;
					// Trace: design.sv:22659:9
					localparam [31:0] Idx0 = ((2 ** level) - 1) + l;
					// Trace: design.sv:22660:9
					localparam [31:0] Idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : gen_reduce
							// Trace: design.sv:22666:13
							assign req_nodes[Idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							// Trace: design.sv:22669:13
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							// Trace: design.sv:22671:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(sel);
							// Trace: design.sv:22672:13
							assign data_nodes[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))] = (sel ? data_i[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + (((l * 2) + 1) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))] : data_i[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((l * 2) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))]);
							// Trace: design.sv:22673:13
							assign gnt_o[l * 2] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							// Trace: design.sv:22674:13
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : gen_first
							// Trace: design.sv:22678:13
							assign req_nodes[Idx0] = req_d[l * 2];
							// Trace: design.sv:22679:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = 1'sb0;
							// Trace: design.sv:22680:13
							assign data_nodes[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))] = data_i[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((l * 2) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))];
							// Trace: design.sv:22681:13
							assign gnt_o[l * 2] = gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : gen_out_of_range
							// Trace: design.sv:22685:13
							assign req_nodes[Idx0] = 1'b0;
							// Trace: design.sv:22686:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(1'sb0);
							// Trace: design.sv:22687:13
							assign data_nodes[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))] = sv2v_cast_5FCB8(1'sb0);
						end
					end
					else begin : gen_other_levels
						// Trace: design.sv:22692:11
						assign req_nodes[Idx0] = req_nodes[Idx1] | req_nodes[Idx1 + 1];
						// Trace: design.sv:22695:11
						assign sel = ~req_nodes[Idx1] | (req_nodes[Idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						// Trace: design.sv:22697:11
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = (sel ? sv2v_cast_5FDFE({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5FDFE({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						// Trace: design.sv:22701:11
						assign data_nodes[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))] = (sel ? data_nodes[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))] : data_nodes[((DataType_Width + 6) >= 0 ? 0 : DataType_Width + 6) + ((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * ((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6)))+:((DataType_Width + 6) >= 0 ? DataType_Width + 7 : 1 - (DataType_Width + 6))]);
						// Trace: design.sv:22702:11
						assign gnt_nodes[Idx1] = gnt_nodes[Idx0] & ~sel;
						// Trace: design.sv:22703:11
						assign gnt_nodes[Idx1 + 1] = gnt_nodes[Idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_93F52 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	req_o,
	gnt_i,
	data_o,
	idx_o
);
	// Trace: design.sv:22448:13
	parameter [31:0] NumIn = 64;
	// Trace: design.sv:22450:13
	parameter [31:0] DataWidth = 32;
	// Trace: design.sv:22452:26
	// removed localparam type DataType
	// Trace: design.sv:22459:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: design.sv:22466:13
	parameter [0:0] AxiVldRdy = 1'b0;
	// Trace: design.sv:22473:13
	parameter [0:0] LockIn = 1'b0;
	// Trace: design.sv:22477:13
	parameter [0:0] FairArb = 1'b1;
	// Trace: design.sv:22480:13
	parameter [31:0] IdxWidth = (NumIn > 32'd1 ? $unsigned($clog2(NumIn)) : 32'd1);
	// Trace: design.sv:22483:26
	// removed localparam type idx_t
	// Trace: design.sv:22486:3
	input wire clk_i;
	// Trace: design.sv:22488:3
	input wire rst_ni;
	// Trace: design.sv:22490:3
	input wire flush_i;
	// Trace: design.sv:22492:3
	input wire [IdxWidth - 1:0] rr_i;
	// Trace: design.sv:22494:3
	input wire [NumIn - 1:0] req_i;
	// Trace: design.sv:22497:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: design.sv:22500:3
	input wire [NumIn - 1:0] data_i;
	// Trace: design.sv:22502:3
	output wire req_o;
	// Trace: design.sv:22504:3
	input wire gnt_i;
	// Trace: design.sv:22506:3
	output wire data_o;
	// Trace: design.sv:22508:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:22521:3
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : gen_pass_through
			// Trace: design.sv:22522:5
			assign req_o = req_i[0];
			// Trace: design.sv:22523:5
			assign gnt_o[0] = gnt_i;
			// Trace: design.sv:22524:5
			assign data_o = data_i[0];
			// Trace: design.sv:22525:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_arbiter
			// Trace: design.sv:22528:5
			localparam [31:0] NumLevels = $unsigned($clog2(NumIn));
			// Trace: design.sv:22531:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * IdxWidth) - 1 : ((3 - (2 ** NumLevels)) * IdxWidth) + ((((2 ** NumLevels) - 2) * IdxWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * IdxWidth)] index_nodes;
			// Trace: design.sv:22532:5
			wire [(2 ** NumLevels) - 2:0] data_nodes;
			// Trace: design.sv:22533:5
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			// Trace: design.sv:22534:5
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			// Trace: design.sv:22536:5
			reg [IdxWidth - 1:0] rr_q;
			// Trace: design.sv:22537:5
			wire [NumIn - 1:0] req_d;
			// Trace: design.sv:22540:5
			assign req_o = req_nodes[0];
			// Trace: design.sv:22541:5
			assign data_o = data_nodes[0];
			// Trace: design.sv:22542:5
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * IdxWidth+:IdxWidth];
			if (ExtPrio) begin : gen_ext_rr
				// Trace: design.sv:22545:7
				wire [IdxWidth:1] sv2v_tmp_0900B;
				assign sv2v_tmp_0900B = rr_i;
				always @(*) rr_q = sv2v_tmp_0900B;
				// Trace: design.sv:22546:7
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				// Trace: design.sv:22548:7
				wire [IdxWidth - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					// Trace: design.sv:22552:9
					wire lock_d;
					reg lock_q;
					// Trace: design.sv:22553:9
					reg [NumIn - 1:0] req_q;
					// Trace: design.sv:22555:9
					assign lock_d = req_o & ~gnt_i;
					// Trace: design.sv:22556:9
					assign req_d = (lock_q ? req_q : req_i);
					// Trace: design.sv:22558:9
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						// Trace: design.sv:22559:11
						if (!rst_ni)
							// Trace: design.sv:22560:13
							lock_q <= 1'sb0;
						else
							// Trace: design.sv:22562:13
							if (flush_i)
								// Trace: design.sv:22563:15
								lock_q <= 1'sb0;
							else
								// Trace: design.sv:22565:15
								lock_q <= lock_d;
					end
					// Trace: design.sv:22587:9
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						// Trace: design.sv:22588:11
						if (!rst_ni)
							// Trace: design.sv:22589:13
							req_q <= 1'sb0;
						else
							// Trace: design.sv:22591:13
							if (flush_i)
								// Trace: design.sv:22592:15
								req_q <= 1'sb0;
							else
								// Trace: design.sv:22594:15
								req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					// Trace: design.sv:22599:9
					assign req_d = req_i;
				end
				if (FairArb) begin : gen_fair_arb
					// Trace: design.sv:22603:9
					wire [NumIn - 1:0] upper_mask;
					wire [NumIn - 1:0] lower_mask;
					// Trace: design.sv:22604:9
					wire [IdxWidth - 1:0] upper_idx;
					wire [IdxWidth - 1:0] lower_idx;
					wire [IdxWidth - 1:0] next_idx;
					// Trace: design.sv:22605:9
					wire upper_empty;
					wire lower_empty;
					genvar _gv_i_9;
					for (_gv_i_9 = 0; _gv_i_9 < NumIn; _gv_i_9 = _gv_i_9 + 1) begin : gen_mask
						localparam i = _gv_i_9;
						// Trace: design.sv:22608:11
						assign upper_mask[i] = (i > rr_q ? req_d[i] : 1'b0);
						// Trace: design.sv:22609:11
						assign lower_mask[i] = (i <= rr_q ? req_d[i] : 1'b0);
					end
					// Trace: design.sv:22612:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_upper(
						.in_i(upper_mask),
						.cnt_o(upper_idx),
						.empty_o(upper_empty)
					);
					// Trace: design.sv:22621:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_lower(
						.in_i(lower_mask),
						.cnt_o(lower_idx),
						.empty_o()
					);
					// Trace: design.sv:22630:9
					assign next_idx = (upper_empty ? lower_idx : upper_idx);
					// Trace: design.sv:22631:9
					assign rr_d = (gnt_i && req_o ? next_idx : rr_q);
				end
				else begin : gen_unfair_arb
					// Trace: design.sv:22634:9
					assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5FDFE(NumIn - 1) ? {IdxWidth {1'sb0}} : rr_q + 1'b1) : rr_q);
				end
				// Trace: design.sv:22638:7
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					// Trace: design.sv:22639:9
					if (!rst_ni)
						// Trace: design.sv:22640:11
						rr_q <= 1'sb0;
					else
						// Trace: design.sv:22642:11
						if (flush_i)
							// Trace: design.sv:22643:13
							rr_q <= 1'sb0;
						else
							// Trace: design.sv:22645:13
							rr_q <= rr_d;
				end
			end
			// Trace: design.sv:22651:5
			assign gnt_nodes[0] = gnt_i;
			genvar _gv_level_2;
			for (_gv_level_2 = 0; $unsigned(_gv_level_2) < NumLevels; _gv_level_2 = _gv_level_2 + 1) begin : gen_levels
				localparam level = _gv_level_2;
				genvar _gv_l_4;
				for (_gv_l_4 = 0; _gv_l_4 < (2 ** level); _gv_l_4 = _gv_l_4 + 1) begin : gen_level
					localparam l = _gv_l_4;
					// Trace: design.sv:22657:9
					wire sel;
					// Trace: design.sv:22659:9
					localparam [31:0] Idx0 = ((2 ** level) - 1) + l;
					// Trace: design.sv:22660:9
					localparam [31:0] Idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : gen_reduce
							// Trace: design.sv:22666:13
							assign req_nodes[Idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							// Trace: design.sv:22669:13
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							// Trace: design.sv:22671:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(sel);
							// Trace: design.sv:22672:13
							assign data_nodes[Idx0] = (sel ? data_i[(l * 2) + 1] : data_i[l * 2]);
							// Trace: design.sv:22673:13
							assign gnt_o[l * 2] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							// Trace: design.sv:22674:13
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : gen_first
							// Trace: design.sv:22678:13
							assign req_nodes[Idx0] = req_d[l * 2];
							// Trace: design.sv:22679:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = 1'sb0;
							// Trace: design.sv:22680:13
							assign data_nodes[Idx0] = data_i[l * 2];
							// Trace: design.sv:22681:13
							assign gnt_o[l * 2] = gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : gen_out_of_range
							// Trace: design.sv:22685:13
							assign req_nodes[Idx0] = 1'b0;
							// Trace: design.sv:22686:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(1'sb0);
							// Trace: design.sv:22687:13
							assign data_nodes[Idx0] = 1'b0;
						end
					end
					else begin : gen_other_levels
						// Trace: design.sv:22692:11
						assign req_nodes[Idx0] = req_nodes[Idx1] | req_nodes[Idx1 + 1];
						// Trace: design.sv:22695:11
						assign sel = ~req_nodes[Idx1] | (req_nodes[Idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						// Trace: design.sv:22697:11
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = (sel ? sv2v_cast_5FDFE({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5FDFE({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						// Trace: design.sv:22701:11
						assign data_nodes[Idx0] = (sel ? data_nodes[Idx1 + 1] : data_nodes[Idx1]);
						// Trace: design.sv:22702:11
						assign gnt_nodes[Idx1] = gnt_nodes[Idx0] & ~sel;
						// Trace: design.sv:22703:11
						assign gnt_nodes[Idx1 + 1] = gnt_nodes[Idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_D7936_86F21 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	req_o,
	gnt_i,
	data_o,
	idx_o
);
	// removed localparam type DataType_payload_t_DataWidth_type
	// removed localparam type DataType_payload_t_IdxWidth_type
	// removed localparam type DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6_type
	parameter [31:0] DataType_payload_t_DataWidth = 0;
	parameter [31:0] DataType_payload_t_IdxWidth = 0;
	parameter integer DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 = 0;
	// Trace: design.sv:22448:13
	parameter [31:0] NumIn = 64;
	// Trace: design.sv:22450:13
	parameter [31:0] DataWidth = 32;
	// Trace: design.sv:22452:26
	// removed localparam type DataType
	// Trace: design.sv:22459:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: design.sv:22466:13
	parameter [0:0] AxiVldRdy = 1'b0;
	// Trace: design.sv:22473:13
	parameter [0:0] LockIn = 1'b0;
	// Trace: design.sv:22477:13
	parameter [0:0] FairArb = 1'b1;
	// Trace: design.sv:22480:13
	parameter [31:0] IdxWidth = (NumIn > 32'd1 ? $unsigned($clog2(NumIn)) : 32'd1);
	// Trace: design.sv:22483:26
	// removed localparam type idx_t
	// Trace: design.sv:22486:3
	input wire clk_i;
	// Trace: design.sv:22488:3
	input wire rst_ni;
	// Trace: design.sv:22490:3
	input wire flush_i;
	// Trace: design.sv:22492:3
	input wire [IdxWidth - 1:0] rr_i;
	// Trace: design.sv:22494:3
	input wire [NumIn - 1:0] req_i;
	// Trace: design.sv:22497:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: design.sv:22500:3
	input wire [(NumIn * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)) - 1:0] data_i;
	// Trace: design.sv:22502:3
	output wire req_o;
	// Trace: design.sv:22504:3
	input wire gnt_i;
	// Trace: design.sv:22506:3
	output wire [((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth) - 1:0] data_o;
	// Trace: design.sv:22508:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:22521:3
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	function automatic [((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth) - 1:0] sv2v_cast_70469;
		input reg [((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth) - 1:0] inp;
		sv2v_cast_70469 = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : gen_pass_through
			// Trace: design.sv:22522:5
			assign req_o = req_i[0];
			// Trace: design.sv:22523:5
			assign gnt_o[0] = gnt_i;
			// Trace: design.sv:22524:5
			assign data_o = data_i[0+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth];
			// Trace: design.sv:22525:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_arbiter
			// Trace: design.sv:22528:5
			localparam [31:0] NumLevels = $unsigned($clog2(NumIn));
			// Trace: design.sv:22531:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * IdxWidth) - 1 : ((3 - (2 ** NumLevels)) * IdxWidth) + ((((2 ** NumLevels) - 2) * IdxWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * IdxWidth)] index_nodes;
			// Trace: design.sv:22532:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)) - 1 : ((3 - (2 ** NumLevels)) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)) + ((((2 ** NumLevels) - 2) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth))] data_nodes;
			// Trace: design.sv:22533:5
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			// Trace: design.sv:22534:5
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			// Trace: design.sv:22536:5
			reg [IdxWidth - 1:0] rr_q;
			// Trace: design.sv:22537:5
			wire [NumIn - 1:0] req_d;
			// Trace: design.sv:22540:5
			assign req_o = req_nodes[0];
			// Trace: design.sv:22541:5
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth];
			// Trace: design.sv:22542:5
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * IdxWidth+:IdxWidth];
			if (ExtPrio) begin : gen_ext_rr
				// Trace: design.sv:22545:7
				wire [IdxWidth:1] sv2v_tmp_0900B;
				assign sv2v_tmp_0900B = rr_i;
				always @(*) rr_q = sv2v_tmp_0900B;
				// Trace: design.sv:22546:7
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				// Trace: design.sv:22548:7
				wire [IdxWidth - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					// Trace: design.sv:22552:9
					wire lock_d;
					reg lock_q;
					// Trace: design.sv:22553:9
					reg [NumIn - 1:0] req_q;
					// Trace: design.sv:22555:9
					assign lock_d = req_o & ~gnt_i;
					// Trace: design.sv:22556:9
					assign req_d = (lock_q ? req_q : req_i);
					// Trace: design.sv:22558:9
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						// Trace: design.sv:22559:11
						if (!rst_ni)
							// Trace: design.sv:22560:13
							lock_q <= 1'sb0;
						else
							// Trace: design.sv:22562:13
							if (flush_i)
								// Trace: design.sv:22563:15
								lock_q <= 1'sb0;
							else
								// Trace: design.sv:22565:15
								lock_q <= lock_d;
					end
					// Trace: design.sv:22587:9
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						// Trace: design.sv:22588:11
						if (!rst_ni)
							// Trace: design.sv:22589:13
							req_q <= 1'sb0;
						else
							// Trace: design.sv:22591:13
							if (flush_i)
								// Trace: design.sv:22592:15
								req_q <= 1'sb0;
							else
								// Trace: design.sv:22594:15
								req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					// Trace: design.sv:22599:9
					assign req_d = req_i;
				end
				if (FairArb) begin : gen_fair_arb
					// Trace: design.sv:22603:9
					wire [NumIn - 1:0] upper_mask;
					wire [NumIn - 1:0] lower_mask;
					// Trace: design.sv:22604:9
					wire [IdxWidth - 1:0] upper_idx;
					wire [IdxWidth - 1:0] lower_idx;
					wire [IdxWidth - 1:0] next_idx;
					// Trace: design.sv:22605:9
					wire upper_empty;
					wire lower_empty;
					genvar _gv_i_9;
					for (_gv_i_9 = 0; _gv_i_9 < NumIn; _gv_i_9 = _gv_i_9 + 1) begin : gen_mask
						localparam i = _gv_i_9;
						// Trace: design.sv:22608:11
						assign upper_mask[i] = (i > rr_q ? req_d[i] : 1'b0);
						// Trace: design.sv:22609:11
						assign lower_mask[i] = (i <= rr_q ? req_d[i] : 1'b0);
					end
					// Trace: design.sv:22612:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_upper(
						.in_i(upper_mask),
						.cnt_o(upper_idx),
						.empty_o(upper_empty)
					);
					// Trace: design.sv:22621:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_lower(
						.in_i(lower_mask),
						.cnt_o(lower_idx),
						.empty_o()
					);
					// Trace: design.sv:22630:9
					assign next_idx = (upper_empty ? lower_idx : upper_idx);
					// Trace: design.sv:22631:9
					assign rr_d = (gnt_i && req_o ? next_idx : rr_q);
				end
				else begin : gen_unfair_arb
					// Trace: design.sv:22634:9
					assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5FDFE(NumIn - 1) ? {IdxWidth {1'sb0}} : rr_q + 1'b1) : rr_q);
				end
				// Trace: design.sv:22638:7
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					// Trace: design.sv:22639:9
					if (!rst_ni)
						// Trace: design.sv:22640:11
						rr_q <= 1'sb0;
					else
						// Trace: design.sv:22642:11
						if (flush_i)
							// Trace: design.sv:22643:13
							rr_q <= 1'sb0;
						else
							// Trace: design.sv:22645:13
							rr_q <= rr_d;
				end
			end
			// Trace: design.sv:22651:5
			assign gnt_nodes[0] = gnt_i;
			genvar _gv_level_2;
			for (_gv_level_2 = 0; $unsigned(_gv_level_2) < NumLevels; _gv_level_2 = _gv_level_2 + 1) begin : gen_levels
				localparam level = _gv_level_2;
				genvar _gv_l_4;
				for (_gv_l_4 = 0; _gv_l_4 < (2 ** level); _gv_l_4 = _gv_l_4 + 1) begin : gen_level
					localparam l = _gv_l_4;
					// Trace: design.sv:22657:9
					wire sel;
					// Trace: design.sv:22659:9
					localparam [31:0] Idx0 = ((2 ** level) - 1) + l;
					// Trace: design.sv:22660:9
					localparam [31:0] Idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : gen_reduce
							// Trace: design.sv:22666:13
							assign req_nodes[Idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							// Trace: design.sv:22669:13
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							// Trace: design.sv:22671:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(sel);
							// Trace: design.sv:22672:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth] = (sel ? data_i[((l * 2) + 1) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth] : data_i[(l * 2) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth]);
							// Trace: design.sv:22673:13
							assign gnt_o[l * 2] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							// Trace: design.sv:22674:13
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : gen_first
							// Trace: design.sv:22678:13
							assign req_nodes[Idx0] = req_d[l * 2];
							// Trace: design.sv:22679:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = 1'sb0;
							// Trace: design.sv:22680:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth] = data_i[(l * 2) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth];
							// Trace: design.sv:22681:13
							assign gnt_o[l * 2] = gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : gen_out_of_range
							// Trace: design.sv:22685:13
							assign req_nodes[Idx0] = 1'b0;
							// Trace: design.sv:22686:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(1'sb0);
							// Trace: design.sv:22687:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth] = sv2v_cast_70469(1'sb0);
						end
					end
					else begin : gen_other_levels
						// Trace: design.sv:22692:11
						assign req_nodes[Idx0] = req_nodes[Idx1] | req_nodes[Idx1 + 1];
						// Trace: design.sv:22695:11
						assign sel = ~req_nodes[Idx1] | (req_nodes[Idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						// Trace: design.sv:22697:11
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = (sel ? sv2v_cast_5FDFE({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5FDFE({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						// Trace: design.sv:22701:11
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * ((DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth)+:(DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + DataType_payload_t_DataWidth) + DataType_payload_t_IdxWidth]);
						// Trace: design.sv:22702:11
						assign gnt_nodes[Idx1] = gnt_nodes[Idx0] & ~sel;
						// Trace: design.sv:22703:11
						assign gnt_nodes[Idx1 + 1] = gnt_nodes[Idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_A5EF3_DDD71 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	req_o,
	gnt_i,
	data_o,
	idx_o
);
	// removed localparam type DataType_WIDTH_type
	parameter [31:0] DataType_WIDTH = 0;
	// Trace: design.sv:22448:13
	parameter [31:0] NumIn = 64;
	// Trace: design.sv:22450:13
	parameter [31:0] DataWidth = 32;
	// Trace: design.sv:22452:26
	// removed localparam type DataType
	// Trace: design.sv:22459:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: design.sv:22466:13
	parameter [0:0] AxiVldRdy = 1'b0;
	// Trace: design.sv:22473:13
	parameter [0:0] LockIn = 1'b0;
	// Trace: design.sv:22477:13
	parameter [0:0] FairArb = 1'b1;
	// Trace: design.sv:22480:13
	parameter [31:0] IdxWidth = (NumIn > 32'd1 ? $unsigned($clog2(NumIn)) : 32'd1);
	// Trace: design.sv:22483:26
	// removed localparam type idx_t
	// Trace: design.sv:22486:3
	input wire clk_i;
	// Trace: design.sv:22488:3
	input wire rst_ni;
	// Trace: design.sv:22490:3
	input wire flush_i;
	// Trace: design.sv:22492:3
	input wire [IdxWidth - 1:0] rr_i;
	// Trace: design.sv:22494:3
	input wire [NumIn - 1:0] req_i;
	// Trace: design.sv:22497:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: design.sv:22500:3
	input wire [((DataType_WIDTH + 5) >= 0 ? (NumIn * (DataType_WIDTH + 6)) - 1 : (NumIn * (1 - (DataType_WIDTH + 5))) + (DataType_WIDTH + 4)):((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5)] data_i;
	// Trace: design.sv:22502:3
	output wire req_o;
	// Trace: design.sv:22504:3
	input wire gnt_i;
	// Trace: design.sv:22506:3
	output wire [DataType_WIDTH + 5:0] data_o;
	// Trace: design.sv:22508:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:22521:3
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	function automatic [((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)) - 1:0] sv2v_cast_7B119;
		input reg [((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)) - 1:0] inp;
		sv2v_cast_7B119 = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : gen_pass_through
			// Trace: design.sv:22522:5
			assign req_o = req_i[0];
			// Trace: design.sv:22523:5
			assign gnt_o[0] = gnt_i;
			// Trace: design.sv:22524:5
			assign data_o = data_i[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + 0+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))];
			// Trace: design.sv:22525:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_arbiter
			// Trace: design.sv:22528:5
			localparam [31:0] NumLevels = $unsigned($clog2(NumIn));
			// Trace: design.sv:22531:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * IdxWidth) - 1 : ((3 - (2 ** NumLevels)) * IdxWidth) + ((((2 ** NumLevels) - 2) * IdxWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * IdxWidth)] index_nodes;
			// Trace: design.sv:22532:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? ((DataType_WIDTH + 5) >= 0 ? (((2 ** NumLevels) - 1) * (DataType_WIDTH + 6)) - 1 : (((2 ** NumLevels) - 1) * (1 - (DataType_WIDTH + 5))) + (DataType_WIDTH + 4)) : ((DataType_WIDTH + 5) >= 0 ? ((3 - (2 ** NumLevels)) * (DataType_WIDTH + 6)) + ((((2 ** NumLevels) - 2) * (DataType_WIDTH + 6)) - 1) : ((3 - (2 ** NumLevels)) * (1 - (DataType_WIDTH + 5))) + (((DataType_WIDTH + 5) + (((2 ** NumLevels) - 2) * (1 - (DataType_WIDTH + 5)))) - 1))):(((2 ** NumLevels) - 2) >= 0 ? ((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) : ((DataType_WIDTH + 5) >= 0 ? ((2 ** NumLevels) - 2) * (DataType_WIDTH + 6) : (DataType_WIDTH + 5) + (((2 ** NumLevels) - 2) * (1 - (DataType_WIDTH + 5)))))] data_nodes;
			// Trace: design.sv:22533:5
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			// Trace: design.sv:22534:5
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			// Trace: design.sv:22536:5
			reg [IdxWidth - 1:0] rr_q;
			// Trace: design.sv:22537:5
			wire [NumIn - 1:0] req_d;
			// Trace: design.sv:22540:5
			assign req_o = req_nodes[0];
			// Trace: design.sv:22541:5
			assign data_o = data_nodes[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))];
			// Trace: design.sv:22542:5
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * IdxWidth+:IdxWidth];
			if (ExtPrio) begin : gen_ext_rr
				// Trace: design.sv:22545:7
				wire [IdxWidth:1] sv2v_tmp_0900B;
				assign sv2v_tmp_0900B = rr_i;
				always @(*) rr_q = sv2v_tmp_0900B;
				// Trace: design.sv:22546:7
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				// Trace: design.sv:22548:7
				wire [IdxWidth - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					// Trace: design.sv:22552:9
					wire lock_d;
					reg lock_q;
					// Trace: design.sv:22553:9
					reg [NumIn - 1:0] req_q;
					// Trace: design.sv:22555:9
					assign lock_d = req_o & ~gnt_i;
					// Trace: design.sv:22556:9
					assign req_d = (lock_q ? req_q : req_i);
					// Trace: design.sv:22558:9
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						// Trace: design.sv:22559:11
						if (!rst_ni)
							// Trace: design.sv:22560:13
							lock_q <= 1'sb0;
						else
							// Trace: design.sv:22562:13
							if (flush_i)
								// Trace: design.sv:22563:15
								lock_q <= 1'sb0;
							else
								// Trace: design.sv:22565:15
								lock_q <= lock_d;
					end
					// Trace: design.sv:22587:9
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						// Trace: design.sv:22588:11
						if (!rst_ni)
							// Trace: design.sv:22589:13
							req_q <= 1'sb0;
						else
							// Trace: design.sv:22591:13
							if (flush_i)
								// Trace: design.sv:22592:15
								req_q <= 1'sb0;
							else
								// Trace: design.sv:22594:15
								req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					// Trace: design.sv:22599:9
					assign req_d = req_i;
				end
				if (FairArb) begin : gen_fair_arb
					// Trace: design.sv:22603:9
					wire [NumIn - 1:0] upper_mask;
					wire [NumIn - 1:0] lower_mask;
					// Trace: design.sv:22604:9
					wire [IdxWidth - 1:0] upper_idx;
					wire [IdxWidth - 1:0] lower_idx;
					wire [IdxWidth - 1:0] next_idx;
					// Trace: design.sv:22605:9
					wire upper_empty;
					wire lower_empty;
					genvar _gv_i_9;
					for (_gv_i_9 = 0; _gv_i_9 < NumIn; _gv_i_9 = _gv_i_9 + 1) begin : gen_mask
						localparam i = _gv_i_9;
						// Trace: design.sv:22608:11
						assign upper_mask[i] = (i > rr_q ? req_d[i] : 1'b0);
						// Trace: design.sv:22609:11
						assign lower_mask[i] = (i <= rr_q ? req_d[i] : 1'b0);
					end
					// Trace: design.sv:22612:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_upper(
						.in_i(upper_mask),
						.cnt_o(upper_idx),
						.empty_o(upper_empty)
					);
					// Trace: design.sv:22621:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_lower(
						.in_i(lower_mask),
						.cnt_o(lower_idx),
						.empty_o()
					);
					// Trace: design.sv:22630:9
					assign next_idx = (upper_empty ? lower_idx : upper_idx);
					// Trace: design.sv:22631:9
					assign rr_d = (gnt_i && req_o ? next_idx : rr_q);
				end
				else begin : gen_unfair_arb
					// Trace: design.sv:22634:9
					assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5FDFE(NumIn - 1) ? {IdxWidth {1'sb0}} : rr_q + 1'b1) : rr_q);
				end
				// Trace: design.sv:22638:7
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					// Trace: design.sv:22639:9
					if (!rst_ni)
						// Trace: design.sv:22640:11
						rr_q <= 1'sb0;
					else
						// Trace: design.sv:22642:11
						if (flush_i)
							// Trace: design.sv:22643:13
							rr_q <= 1'sb0;
						else
							// Trace: design.sv:22645:13
							rr_q <= rr_d;
				end
			end
			// Trace: design.sv:22651:5
			assign gnt_nodes[0] = gnt_i;
			genvar _gv_level_2;
			for (_gv_level_2 = 0; $unsigned(_gv_level_2) < NumLevels; _gv_level_2 = _gv_level_2 + 1) begin : gen_levels
				localparam level = _gv_level_2;
				genvar _gv_l_4;
				for (_gv_l_4 = 0; _gv_l_4 < (2 ** level); _gv_l_4 = _gv_l_4 + 1) begin : gen_level
					localparam l = _gv_l_4;
					// Trace: design.sv:22657:9
					wire sel;
					// Trace: design.sv:22659:9
					localparam [31:0] Idx0 = ((2 ** level) - 1) + l;
					// Trace: design.sv:22660:9
					localparam [31:0] Idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : gen_reduce
							// Trace: design.sv:22666:13
							assign req_nodes[Idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							// Trace: design.sv:22669:13
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							// Trace: design.sv:22671:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(sel);
							// Trace: design.sv:22672:13
							assign data_nodes[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))] = (sel ? data_i[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + (((l * 2) + 1) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))] : data_i[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((l * 2) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))]);
							// Trace: design.sv:22673:13
							assign gnt_o[l * 2] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							// Trace: design.sv:22674:13
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : gen_first
							// Trace: design.sv:22678:13
							assign req_nodes[Idx0] = req_d[l * 2];
							// Trace: design.sv:22679:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = 1'sb0;
							// Trace: design.sv:22680:13
							assign data_nodes[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))] = data_i[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((l * 2) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))];
							// Trace: design.sv:22681:13
							assign gnt_o[l * 2] = gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : gen_out_of_range
							// Trace: design.sv:22685:13
							assign req_nodes[Idx0] = 1'b0;
							// Trace: design.sv:22686:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_5FDFE(1'sb0);
							// Trace: design.sv:22687:13
							assign data_nodes[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))] = sv2v_cast_7B119(1'sb0);
						end
					end
					else begin : gen_other_levels
						// Trace: design.sv:22692:11
						assign req_nodes[Idx0] = req_nodes[Idx1] | req_nodes[Idx1 + 1];
						// Trace: design.sv:22695:11
						assign sel = ~req_nodes[Idx1] | (req_nodes[Idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						// Trace: design.sv:22697:11
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = (sel ? sv2v_cast_5FDFE({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5FDFE({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						// Trace: design.sv:22701:11
						assign data_nodes[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))] = (sel ? data_nodes[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))] : data_nodes[((DataType_WIDTH + 5) >= 0 ? 0 : DataType_WIDTH + 5) + ((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * ((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5)))+:((DataType_WIDTH + 5) >= 0 ? DataType_WIDTH + 6 : 1 - (DataType_WIDTH + 5))]);
						// Trace: design.sv:22702:11
						assign gnt_nodes[Idx1] = gnt_nodes[Idx0] & ~sel;
						// Trace: design.sv:22703:11
						assign gnt_nodes[Idx1 + 1] = gnt_nodes[Idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rstgen_bypass (
	clk_i,
	rst_ni,
	rst_test_mode_ni,
	test_mode_i,
	rst_no,
	init_no
);
	// Trace: design.sv:22763:15
	parameter [31:0] NumRegs = 4;
	// Trace: design.sv:22765:5
	input wire clk_i;
	// Trace: design.sv:22766:5
	input wire rst_ni;
	// Trace: design.sv:22767:5
	input wire rst_test_mode_ni;
	// Trace: design.sv:22768:5
	input wire test_mode_i;
	// Trace: design.sv:22769:5
	output wire rst_no;
	// Trace: design.sv:22770:5
	output wire init_no;
	// Trace: design.sv:22774:5
	wire rst_n;
	// Trace: design.sv:22776:5
	reg [NumRegs - 1:0] synch_regs_q;
	// Trace: design.sv:22779:5
	tc_clk_mux2 i_tc_clk_mux2_rst_n(
		.clk0_i(rst_ni),
		.clk1_i(rst_test_mode_ni),
		.clk_sel_i(test_mode_i),
		.clk_o(rst_n)
	);
	// Trace: design.sv:22786:5
	tc_clk_mux2 i_tc_clk_mux2_rst_no(
		.clk0_i(synch_regs_q[NumRegs - 1]),
		.clk1_i(rst_test_mode_ni),
		.clk_sel_i(test_mode_i),
		.clk_o(rst_no)
	);
	// Trace: design.sv:22793:5
	tc_clk_mux2 i_tc_clk_mux2_init_no(
		.clk0_i(synch_regs_q[NumRegs - 1]),
		.clk1_i(1'b1),
		.clk_sel_i(test_mode_i),
		.clk_o(init_no)
	);
	// Trace: design.sv:22800:5
	always @(posedge clk_i or negedge rst_n)
		// Trace: design.sv:22801:9
		if (~rst_n)
			// Trace: design.sv:22802:13
			synch_regs_q <= 0;
		else
			// Trace: design.sv:22804:13
			synch_regs_q <= {synch_regs_q[NumRegs - 2:0], 1'b1};
endmodule
module serial_deglitch (
	clk_i,
	rst_ni,
	en_i,
	d_i,
	q_o
);
	reg _sv2v_0;
	// Trace: design.sv:22830:15
	parameter [31:0] SIZE = 4;
	// Trace: design.sv:22832:5
	input wire clk_i;
	// Trace: design.sv:22833:5
	input wire rst_ni;
	// Trace: design.sv:22834:5
	input wire en_i;
	// Trace: design.sv:22835:5
	input wire d_i;
	// Trace: design.sv:22836:5
	output reg q_o;
	// Trace: design.sv:22838:5
	reg [SIZE - 1:0] count_q;
	// Trace: design.sv:22839:5
	reg q;
	// Trace: design.sv:22841:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:22842:9
		if (~rst_ni) begin
			// Trace: design.sv:22843:13
			count_q <= 1'sb0;
			// Trace: design.sv:22844:13
			q <= 1'b0;
		end
		else
			// Trace: design.sv:22846:13
			if (en_i) begin
				begin
					// Trace: design.sv:22847:17
					if ((d_i == 1'b1) && (count_q != SIZE[SIZE - 1:0]))
						// Trace: design.sv:22848:21
						count_q <= count_q + 1;
					else if ((d_i == 1'b0) && (count_q != SIZE[SIZE - 1:0]))
						// Trace: design.sv:22850:21
						count_q <= count_q - 1;
				end
			end
	// Trace: design.sv:22857:5
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:22858:9
		if (count_q == SIZE[SIZE - 1:0])
			// Trace: design.sv:22859:13
			q_o = 1'b1;
		else if (count_q == 0)
			// Trace: design.sv:22861:13
			q_o = 1'b0;
	end
	initial _sv2v_0 = 0;
endmodule
module shift_reg (
	clk_i,
	rst_ni,
	d_i,
	d_o
);
	// Trace: design.sv:22881:20
	// removed localparam type dtype
	// Trace: design.sv:22882:15
	parameter [31:0] Depth = 1;
	// Trace: design.sv:22884:5
	input wire clk_i;
	// Trace: design.sv:22885:5
	input wire rst_ni;
	// Trace: design.sv:22886:5
	input wire d_i;
	// Trace: design.sv:22887:5
	output reg d_o;
	// Trace: design.sv:22891:5
	generate
		if (Depth == 0) begin : gen_pass_through
			// Trace: design.sv:22892:9
			wire [1:1] sv2v_tmp_D60D7;
			assign sv2v_tmp_D60D7 = d_i;
			always @(*) d_o = sv2v_tmp_D60D7;
		end
		else if (Depth == 1) begin : gen_register
			// Trace: design.sv:22895:9
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:22896:13
				if (~rst_ni)
					// Trace: design.sv:22897:17
					d_o <= 1'sb0;
				else
					// Trace: design.sv:22899:17
					d_o <= d_i;
		end
		else if (Depth > 1) begin : gen_shift_reg
			// Trace: design.sv:22904:9
			wire [Depth - 1:0] reg_d;
			reg [Depth - 1:0] reg_q;
			// Trace: design.sv:22905:9
			wire [1:1] sv2v_tmp_EA7F3;
			assign sv2v_tmp_EA7F3 = reg_q[Depth - 1];
			always @(*) d_o = sv2v_tmp_EA7F3;
			// Trace: design.sv:22906:9
			assign reg_d = {reg_q[Depth - 2:0], d_i};
			// Trace: design.sv:22908:9
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:22909:13
				if (~rst_ni)
					// Trace: design.sv:22910:17
					reg_q <= 1'sb0;
				else
					// Trace: design.sv:22912:17
					reg_q <= reg_d;
		end
	endgenerate
endmodule
module spill_register_flushable_02CF4_D1AAE (
	clk_i,
	rst_ni,
	valid_i,
	flush_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// removed localparam type T_T_T_WIDTH_type
	parameter [31:0] T_T_T_WIDTH = 0;
	// Trace: design.sv:22935:18
	// removed localparam type T
	// Trace: design.sv:22936:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:22938:3
	input wire clk_i;
	// Trace: design.sv:22939:3
	input wire rst_ni;
	// Trace: design.sv:22940:3
	input wire valid_i;
	// Trace: design.sv:22941:3
	input wire flush_i;
	// Trace: design.sv:22942:3
	output wire ready_o;
	// Trace: design.sv:22943:3
	input wire [T_T_T_WIDTH - 1:0] data_i;
	// Trace: design.sv:22944:3
	output wire valid_o;
	// Trace: design.sv:22945:3
	input wire ready_i;
	// Trace: design.sv:22946:3
	output wire [T_T_T_WIDTH - 1:0] data_o;
	// Trace: design.sv:22949:3
	generate
		if (Bypass) begin : gen_bypass
			// Trace: design.sv:22950:5
			assign valid_o = valid_i;
			// Trace: design.sv:22951:5
			assign ready_o = ready_i;
			// Trace: design.sv:22952:5
			assign data_o = data_i;
		end
		else begin : gen_spill_reg
			// Trace: design.sv:22955:5
			reg [T_T_T_WIDTH - 1:0] a_data_q;
			// Trace: design.sv:22956:5
			reg a_full_q;
			// Trace: design.sv:22957:5
			wire a_fill;
			wire a_drain;
			// Trace: design.sv:22959:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_data
				// Trace: design.sv:22960:7
				if (!rst_ni)
					// Trace: design.sv:22961:9
					a_data_q <= 1'sb0;
				else if (a_fill)
					// Trace: design.sv:22963:9
					a_data_q <= data_i;
			end
			// Trace: design.sv:22966:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_full
				// Trace: design.sv:22967:7
				if (!rst_ni)
					// Trace: design.sv:22968:9
					a_full_q <= 0;
				else if (a_fill || a_drain)
					// Trace: design.sv:22970:9
					a_full_q <= a_fill;
			end
			// Trace: design.sv:22974:5
			reg [T_T_T_WIDTH - 1:0] b_data_q;
			// Trace: design.sv:22975:5
			reg b_full_q;
			// Trace: design.sv:22976:5
			wire b_fill;
			wire b_drain;
			// Trace: design.sv:22978:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_data
				// Trace: design.sv:22979:7
				if (!rst_ni)
					// Trace: design.sv:22980:9
					b_data_q <= 1'sb0;
				else if (b_fill)
					// Trace: design.sv:22982:9
					b_data_q <= a_data_q;
			end
			// Trace: design.sv:22985:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_full
				// Trace: design.sv:22986:7
				if (!rst_ni)
					// Trace: design.sv:22987:9
					b_full_q <= 0;
				else if (b_fill || b_drain)
					// Trace: design.sv:22989:9
					b_full_q <= b_fill;
			end
			// Trace: design.sv:22994:5
			assign a_fill = (valid_i && ready_o) && !flush_i;
			// Trace: design.sv:22995:5
			assign a_drain = (a_full_q && !b_full_q) || flush_i;
			// Trace: design.sv:23000:5
			assign b_fill = (a_drain && !ready_i) && !flush_i;
			// Trace: design.sv:23001:5
			assign b_drain = (b_full_q && ready_i) || flush_i;
			// Trace: design.sv:23006:5
			assign ready_o = !a_full_q || !b_full_q;
			// Trace: design.sv:23009:5
			assign valid_o = a_full_q | b_full_q;
			// Trace: design.sv:23012:5
			assign data_o = (b_full_q ? b_data_q : a_data_q);
		end
	endgenerate
endmodule
module spill_register_flushable_918B4_7E477 (
	clk_i,
	rst_ni,
	valid_i,
	flush_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// removed localparam type T_T_IdxWidth_type
	// removed localparam type T_T_payload_t_DataWidth_type
	parameter [31:0] T_T_IdxWidth = 0;
	parameter [31:0] T_T_payload_t_DataWidth = 0;
	// Trace: design.sv:22935:18
	// removed localparam type T
	// Trace: design.sv:22936:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:22938:3
	input wire clk_i;
	// Trace: design.sv:22939:3
	input wire rst_ni;
	// Trace: design.sv:22940:3
	input wire valid_i;
	// Trace: design.sv:22941:3
	input wire flush_i;
	// Trace: design.sv:22942:3
	output wire ready_o;
	// Trace: design.sv:22943:3
	input wire [(T_T_payload_t_DataWidth + T_T_IdxWidth) - 1:0] data_i;
	// Trace: design.sv:22944:3
	output wire valid_o;
	// Trace: design.sv:22945:3
	input wire ready_i;
	// Trace: design.sv:22946:3
	output wire [(T_T_payload_t_DataWidth + T_T_IdxWidth) - 1:0] data_o;
	// Trace: design.sv:22949:3
	generate
		if (Bypass) begin : gen_bypass
			// Trace: design.sv:22950:5
			assign valid_o = valid_i;
			// Trace: design.sv:22951:5
			assign ready_o = ready_i;
			// Trace: design.sv:22952:5
			assign data_o = data_i;
		end
		else begin : gen_spill_reg
			// Trace: design.sv:22955:5
			reg [(T_T_payload_t_DataWidth + T_T_IdxWidth) - 1:0] a_data_q;
			// Trace: design.sv:22956:5
			reg a_full_q;
			// Trace: design.sv:22957:5
			wire a_fill;
			wire a_drain;
			// Trace: design.sv:22959:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_data
				// Trace: design.sv:22960:7
				if (!rst_ni)
					// Trace: design.sv:22961:9
					a_data_q <= 1'sb0;
				else if (a_fill)
					// Trace: design.sv:22963:9
					a_data_q <= data_i;
			end
			// Trace: design.sv:22966:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_full
				// Trace: design.sv:22967:7
				if (!rst_ni)
					// Trace: design.sv:22968:9
					a_full_q <= 0;
				else if (a_fill || a_drain)
					// Trace: design.sv:22970:9
					a_full_q <= a_fill;
			end
			// Trace: design.sv:22974:5
			reg [(T_T_payload_t_DataWidth + T_T_IdxWidth) - 1:0] b_data_q;
			// Trace: design.sv:22975:5
			reg b_full_q;
			// Trace: design.sv:22976:5
			wire b_fill;
			wire b_drain;
			// Trace: design.sv:22978:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_data
				// Trace: design.sv:22979:7
				if (!rst_ni)
					// Trace: design.sv:22980:9
					b_data_q <= 1'sb0;
				else if (b_fill)
					// Trace: design.sv:22982:9
					b_data_q <= a_data_q;
			end
			// Trace: design.sv:22985:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_full
				// Trace: design.sv:22986:7
				if (!rst_ni)
					// Trace: design.sv:22987:9
					b_full_q <= 0;
				else if (b_fill || b_drain)
					// Trace: design.sv:22989:9
					b_full_q <= b_fill;
			end
			// Trace: design.sv:22994:5
			assign a_fill = (valid_i && ready_o) && !flush_i;
			// Trace: design.sv:22995:5
			assign a_drain = (a_full_q && !b_full_q) || flush_i;
			// Trace: design.sv:23000:5
			assign b_fill = (a_drain && !ready_i) && !flush_i;
			// Trace: design.sv:23001:5
			assign b_drain = (b_full_q && ready_i) || flush_i;
			// Trace: design.sv:23006:5
			assign ready_o = !a_full_q || !b_full_q;
			// Trace: design.sv:23009:5
			assign valid_o = a_full_q | b_full_q;
			// Trace: design.sv:23012:5
			assign data_o = (b_full_q ? b_data_q : a_data_q);
		end
	endgenerate
endmodule
module spill_register_flushable_AEB2B_E8B2C (
	clk_i,
	rst_ni,
	valid_i,
	flush_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// removed localparam type T_T_IdxWidth_type
	// removed localparam type T_T_payload_t_DataWidth_type
	// removed localparam type T_T_payload_t_IdxWidth_type
	// removed localparam type T_T_payload_t_i_stream_xbar_sv2v_pfunc_944F6_type
	parameter [31:0] T_T_IdxWidth = 0;
	parameter [31:0] T_T_payload_t_DataWidth = 0;
	parameter [31:0] T_T_payload_t_IdxWidth = 0;
	parameter integer T_T_payload_t_i_stream_xbar_sv2v_pfunc_944F6 = 0;
	// Trace: design.sv:22935:18
	// removed localparam type T
	// Trace: design.sv:22936:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:22938:3
	input wire clk_i;
	// Trace: design.sv:22939:3
	input wire rst_ni;
	// Trace: design.sv:22940:3
	input wire valid_i;
	// Trace: design.sv:22941:3
	input wire flush_i;
	// Trace: design.sv:22942:3
	output wire ready_o;
	// Trace: design.sv:22943:3
	input wire [(((T_T_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + T_T_payload_t_DataWidth) + T_T_payload_t_IdxWidth) + T_T_IdxWidth) - 1:0] data_i;
	// Trace: design.sv:22944:3
	output wire valid_o;
	// Trace: design.sv:22945:3
	input wire ready_i;
	// Trace: design.sv:22946:3
	output wire [(((T_T_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + T_T_payload_t_DataWidth) + T_T_payload_t_IdxWidth) + T_T_IdxWidth) - 1:0] data_o;
	// Trace: design.sv:22949:3
	generate
		if (Bypass) begin : gen_bypass
			// Trace: design.sv:22950:5
			assign valid_o = valid_i;
			// Trace: design.sv:22951:5
			assign ready_o = ready_i;
			// Trace: design.sv:22952:5
			assign data_o = data_i;
		end
		else begin : gen_spill_reg
			// Trace: design.sv:22955:5
			reg [(((T_T_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + T_T_payload_t_DataWidth) + T_T_payload_t_IdxWidth) + T_T_IdxWidth) - 1:0] a_data_q;
			// Trace: design.sv:22956:5
			reg a_full_q;
			// Trace: design.sv:22957:5
			wire a_fill;
			wire a_drain;
			// Trace: design.sv:22959:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_data
				// Trace: design.sv:22960:7
				if (!rst_ni)
					// Trace: design.sv:22961:9
					a_data_q <= 1'sb0;
				else if (a_fill)
					// Trace: design.sv:22963:9
					a_data_q <= data_i;
			end
			// Trace: design.sv:22966:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_full
				// Trace: design.sv:22967:7
				if (!rst_ni)
					// Trace: design.sv:22968:9
					a_full_q <= 0;
				else if (a_fill || a_drain)
					// Trace: design.sv:22970:9
					a_full_q <= a_fill;
			end
			// Trace: design.sv:22974:5
			reg [(((T_T_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + T_T_payload_t_DataWidth) + T_T_payload_t_IdxWidth) + T_T_IdxWidth) - 1:0] b_data_q;
			// Trace: design.sv:22975:5
			reg b_full_q;
			// Trace: design.sv:22976:5
			wire b_fill;
			wire b_drain;
			// Trace: design.sv:22978:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_data
				// Trace: design.sv:22979:7
				if (!rst_ni)
					// Trace: design.sv:22980:9
					b_data_q <= 1'sb0;
				else if (b_fill)
					// Trace: design.sv:22982:9
					b_data_q <= a_data_q;
			end
			// Trace: design.sv:22985:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_full
				// Trace: design.sv:22986:7
				if (!rst_ni)
					// Trace: design.sv:22987:9
					b_full_q <= 0;
				else if (b_fill || b_drain)
					// Trace: design.sv:22989:9
					b_full_q <= b_fill;
			end
			// Trace: design.sv:22994:5
			assign a_fill = (valid_i && ready_o) && !flush_i;
			// Trace: design.sv:22995:5
			assign a_drain = (a_full_q && !b_full_q) || flush_i;
			// Trace: design.sv:23000:5
			assign b_fill = (a_drain && !ready_i) && !flush_i;
			// Trace: design.sv:23001:5
			assign b_drain = (b_full_q && ready_i) || flush_i;
			// Trace: design.sv:23006:5
			assign ready_o = !a_full_q || !b_full_q;
			// Trace: design.sv:23009:5
			assign valid_o = a_full_q | b_full_q;
			// Trace: design.sv:23012:5
			assign data_o = (b_full_q ? b_data_q : a_data_q);
		end
	endgenerate
endmodule
module spill_register_flushable_44288_566E2 (
	clk_i,
	rst_ni,
	valid_i,
	flush_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// removed localparam type T_T_WIDTH_type
	parameter [31:0] T_T_WIDTH = 0;
	// Trace: design.sv:22935:18
	// removed localparam type T
	// Trace: design.sv:22936:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:22938:3
	input wire clk_i;
	// Trace: design.sv:22939:3
	input wire rst_ni;
	// Trace: design.sv:22940:3
	input wire valid_i;
	// Trace: design.sv:22941:3
	input wire flush_i;
	// Trace: design.sv:22942:3
	output wire ready_o;
	// Trace: design.sv:22943:3
	input wire [T_T_WIDTH - 1:0] data_i;
	// Trace: design.sv:22944:3
	output wire valid_o;
	// Trace: design.sv:22945:3
	input wire ready_i;
	// Trace: design.sv:22946:3
	output wire [T_T_WIDTH - 1:0] data_o;
	// Trace: design.sv:22949:3
	generate
		if (Bypass) begin : gen_bypass
			// Trace: design.sv:22950:5
			assign valid_o = valid_i;
			// Trace: design.sv:22951:5
			assign ready_o = ready_i;
			// Trace: design.sv:22952:5
			assign data_o = data_i;
		end
		else begin : gen_spill_reg
			// Trace: design.sv:22955:5
			reg [T_T_WIDTH - 1:0] a_data_q;
			// Trace: design.sv:22956:5
			reg a_full_q;
			// Trace: design.sv:22957:5
			wire a_fill;
			wire a_drain;
			// Trace: design.sv:22959:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_data
				// Trace: design.sv:22960:7
				if (!rst_ni)
					// Trace: design.sv:22961:9
					a_data_q <= 1'sb0;
				else if (a_fill)
					// Trace: design.sv:22963:9
					a_data_q <= data_i;
			end
			// Trace: design.sv:22966:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_full
				// Trace: design.sv:22967:7
				if (!rst_ni)
					// Trace: design.sv:22968:9
					a_full_q <= 0;
				else if (a_fill || a_drain)
					// Trace: design.sv:22970:9
					a_full_q <= a_fill;
			end
			// Trace: design.sv:22974:5
			reg [T_T_WIDTH - 1:0] b_data_q;
			// Trace: design.sv:22975:5
			reg b_full_q;
			// Trace: design.sv:22976:5
			wire b_fill;
			wire b_drain;
			// Trace: design.sv:22978:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_data
				// Trace: design.sv:22979:7
				if (!rst_ni)
					// Trace: design.sv:22980:9
					b_data_q <= 1'sb0;
				else if (b_fill)
					// Trace: design.sv:22982:9
					b_data_q <= a_data_q;
			end
			// Trace: design.sv:22985:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_full
				// Trace: design.sv:22986:7
				if (!rst_ni)
					// Trace: design.sv:22987:9
					b_full_q <= 0;
				else if (b_fill || b_drain)
					// Trace: design.sv:22989:9
					b_full_q <= b_fill;
			end
			// Trace: design.sv:22994:5
			assign a_fill = (valid_i && ready_o) && !flush_i;
			// Trace: design.sv:22995:5
			assign a_drain = (a_full_q && !b_full_q) || flush_i;
			// Trace: design.sv:23000:5
			assign b_fill = (a_drain && !ready_i) && !flush_i;
			// Trace: design.sv:23001:5
			assign b_drain = (b_full_q && ready_i) || flush_i;
			// Trace: design.sv:23006:5
			assign ready_o = !a_full_q || !b_full_q;
			// Trace: design.sv:23009:5
			assign valid_o = a_full_q | b_full_q;
			// Trace: design.sv:23012:5
			assign data_o = (b_full_q ? b_data_q : a_data_q);
		end
	endgenerate
endmodule
module spill_register_flushable_F9055 (
	clk_i,
	rst_ni,
	valid_i,
	flush_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// Trace: design.sv:22935:18
	// removed localparam type T
	// Trace: design.sv:22936:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:22938:3
	input wire clk_i;
	// Trace: design.sv:22939:3
	input wire rst_ni;
	// Trace: design.sv:22940:3
	input wire valid_i;
	// Trace: design.sv:22941:3
	input wire flush_i;
	// Trace: design.sv:22942:3
	output wire ready_o;
	// Trace: design.sv:22943:3
	input wire [1:0] data_i;
	// Trace: design.sv:22944:3
	output wire valid_o;
	// Trace: design.sv:22945:3
	input wire ready_i;
	// Trace: design.sv:22946:3
	output wire [1:0] data_o;
	// Trace: design.sv:22949:3
	generate
		if (Bypass) begin : gen_bypass
			// Trace: design.sv:22950:5
			assign valid_o = valid_i;
			// Trace: design.sv:22951:5
			assign ready_o = ready_i;
			// Trace: design.sv:22952:5
			assign data_o = data_i;
		end
		else begin : gen_spill_reg
			// Trace: design.sv:22955:5
			reg [1:0] a_data_q;
			// Trace: design.sv:22956:5
			reg a_full_q;
			// Trace: design.sv:22957:5
			wire a_fill;
			wire a_drain;
			// Trace: design.sv:22959:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_data
				// Trace: design.sv:22960:7
				if (!rst_ni)
					// Trace: design.sv:22961:9
					a_data_q <= 1'sb0;
				else if (a_fill)
					// Trace: design.sv:22963:9
					a_data_q <= data_i;
			end
			// Trace: design.sv:22966:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_full
				// Trace: design.sv:22967:7
				if (!rst_ni)
					// Trace: design.sv:22968:9
					a_full_q <= 0;
				else if (a_fill || a_drain)
					// Trace: design.sv:22970:9
					a_full_q <= a_fill;
			end
			// Trace: design.sv:22974:5
			reg [1:0] b_data_q;
			// Trace: design.sv:22975:5
			reg b_full_q;
			// Trace: design.sv:22976:5
			wire b_fill;
			wire b_drain;
			// Trace: design.sv:22978:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_data
				// Trace: design.sv:22979:7
				if (!rst_ni)
					// Trace: design.sv:22980:9
					b_data_q <= 1'sb0;
				else if (b_fill)
					// Trace: design.sv:22982:9
					b_data_q <= a_data_q;
			end
			// Trace: design.sv:22985:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_full
				// Trace: design.sv:22986:7
				if (!rst_ni)
					// Trace: design.sv:22987:9
					b_full_q <= 0;
				else if (b_fill || b_drain)
					// Trace: design.sv:22989:9
					b_full_q <= b_fill;
			end
			// Trace: design.sv:22994:5
			assign a_fill = (valid_i && ready_o) && !flush_i;
			// Trace: design.sv:22995:5
			assign a_drain = (a_full_q && !b_full_q) || flush_i;
			// Trace: design.sv:23000:5
			assign b_fill = (a_drain && !ready_i) && !flush_i;
			// Trace: design.sv:23001:5
			assign b_drain = (b_full_q && ready_i) || flush_i;
			// Trace: design.sv:23006:5
			assign ready_o = !a_full_q || !b_full_q;
			// Trace: design.sv:23009:5
			assign valid_o = a_full_q | b_full_q;
			// Trace: design.sv:23012:5
			assign data_o = (b_full_q ? b_data_q : a_data_q);
		end
	endgenerate
endmodule
module spill_register_flushable_D072E (
	clk_i,
	rst_ni,
	valid_i,
	flush_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// Trace: design.sv:22935:18
	// removed localparam type T
	// Trace: design.sv:22936:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:22938:3
	input wire clk_i;
	// Trace: design.sv:22939:3
	input wire rst_ni;
	// Trace: design.sv:22940:3
	input wire valid_i;
	// Trace: design.sv:22941:3
	input wire flush_i;
	// Trace: design.sv:22942:3
	output wire ready_o;
	// Trace: design.sv:22943:3
	input wire data_i;
	// Trace: design.sv:22944:3
	output wire valid_o;
	// Trace: design.sv:22945:3
	input wire ready_i;
	// Trace: design.sv:22946:3
	output wire data_o;
	// Trace: design.sv:22949:3
	generate
		if (Bypass) begin : gen_bypass
			// Trace: design.sv:22950:5
			assign valid_o = valid_i;
			// Trace: design.sv:22951:5
			assign ready_o = ready_i;
			// Trace: design.sv:22952:5
			assign data_o = data_i;
		end
		else begin : gen_spill_reg
			// Trace: design.sv:22955:5
			reg a_data_q;
			// Trace: design.sv:22956:5
			reg a_full_q;
			// Trace: design.sv:22957:5
			wire a_fill;
			wire a_drain;
			// Trace: design.sv:22959:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_data
				// Trace: design.sv:22960:7
				if (!rst_ni)
					// Trace: design.sv:22961:9
					a_data_q <= 1'sb0;
				else if (a_fill)
					// Trace: design.sv:22963:9
					a_data_q <= data_i;
			end
			// Trace: design.sv:22966:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_a_full
				// Trace: design.sv:22967:7
				if (!rst_ni)
					// Trace: design.sv:22968:9
					a_full_q <= 0;
				else if (a_fill || a_drain)
					// Trace: design.sv:22970:9
					a_full_q <= a_fill;
			end
			// Trace: design.sv:22974:5
			reg b_data_q;
			// Trace: design.sv:22975:5
			reg b_full_q;
			// Trace: design.sv:22976:5
			wire b_fill;
			wire b_drain;
			// Trace: design.sv:22978:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_data
				// Trace: design.sv:22979:7
				if (!rst_ni)
					// Trace: design.sv:22980:9
					b_data_q <= 1'sb0;
				else if (b_fill)
					// Trace: design.sv:22982:9
					b_data_q <= a_data_q;
			end
			// Trace: design.sv:22985:5
			always @(posedge clk_i or negedge rst_ni) begin : ps_b_full
				// Trace: design.sv:22986:7
				if (!rst_ni)
					// Trace: design.sv:22987:9
					b_full_q <= 0;
				else if (b_fill || b_drain)
					// Trace: design.sv:22989:9
					b_full_q <= b_fill;
			end
			// Trace: design.sv:22994:5
			assign a_fill = (valid_i && ready_o) && !flush_i;
			// Trace: design.sv:22995:5
			assign a_drain = (a_full_q && !b_full_q) || flush_i;
			// Trace: design.sv:23000:5
			assign b_fill = (a_drain && !ready_i) && !flush_i;
			// Trace: design.sv:23001:5
			assign b_drain = (b_full_q && ready_i) || flush_i;
			// Trace: design.sv:23006:5
			assign ready_o = !a_full_q || !b_full_q;
			// Trace: design.sv:23009:5
			assign valid_o = a_full_q | b_full_q;
			// Trace: design.sv:23012:5
			assign data_o = (b_full_q ? b_data_q : a_data_q);
		end
	endgenerate
endmodule
module stream_demux (
	inp_valid_i,
	inp_ready_o,
	oup_sel_i,
	oup_valid_o,
	oup_ready_i
);
	reg _sv2v_0;
	// Trace: design.sv:23039:13
	parameter [31:0] N_OUP = 32'd1;
	// Trace: design.sv:23041:13
	parameter [31:0] LOG_N_OUP = (N_OUP > 32'd1 ? $unsigned($clog2(N_OUP)) : 1'b1);
	// Trace: design.sv:23043:3
	input wire inp_valid_i;
	// Trace: design.sv:23044:3
	output wire inp_ready_o;
	// Trace: design.sv:23046:3
	input wire [LOG_N_OUP - 1:0] oup_sel_i;
	// Trace: design.sv:23048:3
	output reg [N_OUP - 1:0] oup_valid_o;
	// Trace: design.sv:23049:3
	input wire [N_OUP - 1:0] oup_ready_i;
	// Trace: design.sv:23052:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:23053:5
		oup_valid_o = 1'sb0;
		// Trace: design.sv:23054:5
		oup_valid_o[oup_sel_i] = inp_valid_i;
	end
	// Trace: design.sv:23056:3
	assign inp_ready_o = oup_ready_i[oup_sel_i];
	initial _sv2v_0 = 0;
endmodule
module stream_filter (
	valid_i,
	ready_o,
	drop_i,
	valid_o,
	ready_i
);
	// Trace: design.sv:23072:5
	input wire valid_i;
	// Trace: design.sv:23073:5
	output wire ready_o;
	// Trace: design.sv:23075:5
	input wire drop_i;
	// Trace: design.sv:23077:5
	output wire valid_o;
	// Trace: design.sv:23078:5
	input wire ready_i;
	// Trace: design.sv:23081:5
	assign valid_o = (drop_i ? 1'b0 : valid_i);
	// Trace: design.sv:23082:5
	assign ready_o = (drop_i ? 1'b1 : ready_i);
endmodule
module stream_fork (
	clk_i,
	rst_ni,
	valid_i,
	ready_o,
	valid_o,
	ready_i
);
	reg _sv2v_0;
	// Trace: design.sv:23104:15
	parameter [31:0] N_OUP = 0;
	// Trace: design.sv:23106:5
	input wire clk_i;
	// Trace: design.sv:23107:5
	input wire rst_ni;
	// Trace: design.sv:23108:5
	input wire valid_i;
	// Trace: design.sv:23109:5
	output reg ready_o;
	// Trace: design.sv:23110:5
	output reg [N_OUP - 1:0] valid_o;
	// Trace: design.sv:23111:5
	input wire [N_OUP - 1:0] ready_i;
	// Trace: design.sv:23114:5
	// removed localparam type state_t
	// Trace: design.sv:23116:5
	reg [N_OUP - 1:0] oup_ready;
	wire [N_OUP - 1:0] all_ones;
	// Trace: design.sv:23119:5
	reg inp_state_d;
	reg inp_state_q;
	// Trace: design.sv:23122:5
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:23124:9
		inp_state_d = inp_state_q;
		// Trace: design.sv:23126:9
		(* full_case, parallel_case *)
		case (inp_state_q)
			1'd0:
				// Trace: design.sv:23128:17
				if (valid_i) begin
					begin
						// Trace: design.sv:23129:21
						if ((valid_o == all_ones) && (ready_i == all_ones))
							// Trace: design.sv:23131:25
							ready_o = 1'b1;
						else begin
							// Trace: design.sv:23133:25
							ready_o = 1'b0;
							// Trace: design.sv:23135:25
							inp_state_d = 1'd1;
						end
					end
				end
				else
					// Trace: design.sv:23138:21
					ready_o = 1'b0;
			1'd1:
				// Trace: design.sv:23142:17
				if (valid_i && (oup_ready == all_ones)) begin
					// Trace: design.sv:23143:21
					ready_o = 1'b1;
					// Trace: design.sv:23144:21
					inp_state_d = 1'd0;
				end
				else
					// Trace: design.sv:23146:21
					ready_o = 1'b0;
			default: begin
				// Trace: design.sv:23150:17
				inp_state_d = 1'd0;
				// Trace: design.sv:23151:17
				ready_o = 1'b0;
			end
		endcase
	end
	// Trace: design.sv:23156:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:23157:9
		if (!rst_ni)
			// Trace: design.sv:23158:13
			inp_state_q <= 1'd0;
		else
			// Trace: design.sv:23160:13
			inp_state_q <= inp_state_d;
	// Trace: design.sv:23165:5
	genvar _gv_i_10;
	generate
		for (_gv_i_10 = 0; _gv_i_10 < N_OUP; _gv_i_10 = _gv_i_10 + 1) begin : gen_oup_state
			localparam i = _gv_i_10;
			// Trace: design.sv:23166:9
			reg oup_state_d;
			reg oup_state_q;
			// Trace: design.sv:23168:9
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:23169:13
				oup_ready[i] = 1'b1;
				// Trace: design.sv:23170:13
				valid_o[i] = 1'b0;
				// Trace: design.sv:23171:13
				oup_state_d = oup_state_q;
				// Trace: design.sv:23173:13
				(* full_case, parallel_case *)
				case (oup_state_q)
					1'd0:
						// Trace: design.sv:23175:21
						if (valid_i) begin
							// Trace: design.sv:23176:25
							valid_o[i] = 1'b1;
							// Trace: design.sv:23177:25
							if (ready_i[i]) begin
								begin
									// Trace: design.sv:23178:29
									if (!ready_o)
										// Trace: design.sv:23179:33
										oup_state_d = 1'd1;
								end
							end
							else
								// Trace: design.sv:23182:29
								oup_ready[i] = 1'b0;
						end
					1'd1:
						// Trace: design.sv:23187:21
						if (valid_i && ready_o)
							// Trace: design.sv:23188:25
							oup_state_d = 1'd0;
					default:
						// Trace: design.sv:23192:21
						oup_state_d = 1'd0;
				endcase
			end
			// Trace: design.sv:23197:9
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:23198:13
				if (!rst_ni)
					// Trace: design.sv:23199:17
					oup_state_q <= 1'd0;
				else
					// Trace: design.sv:23201:17
					oup_state_q <= oup_state_d;
		end
	endgenerate
	// Trace: design.sv:23206:5
	assign all_ones = 1'sb1;
	initial _sv2v_0 = 0;
endmodule
// removed interface: STREAM_DV
module stream_join (
	inp_valid_i,
	inp_ready_o,
	oup_valid_o,
	oup_ready_i
);
	// Trace: design.sv:23285:13
	parameter [31:0] N_INP = 32'd0;
	// Trace: design.sv:23288:3
	input wire [N_INP - 1:0] inp_valid_i;
	// Trace: design.sv:23290:3
	output wire [N_INP - 1:0] inp_ready_o;
	// Trace: design.sv:23292:3
	output wire oup_valid_o;
	// Trace: design.sv:23294:3
	input wire oup_ready_i;
	// Trace: design.sv:23297:3
	assign oup_valid_o = &inp_valid_i;
	// Trace: design.sv:23298:3
	genvar _gv_i_11;
	generate
		for (_gv_i_11 = 0; _gv_i_11 < N_INP; _gv_i_11 = _gv_i_11 + 1) begin : gen_inp_ready
			localparam i = _gv_i_11;
			// Trace: design.sv:23299:5
			assign inp_ready_o[i] = oup_valid_o & oup_ready_i;
		end
	endgenerate
endmodule
module stream_mux (
	inp_data_i,
	inp_valid_i,
	inp_ready_o,
	inp_sel_i,
	oup_data_o,
	oup_valid_o,
	oup_ready_i
);
	reg _sv2v_0;
	// Trace: design.sv:23324:18
	// removed localparam type DATA_T
	// Trace: design.sv:23325:13
	parameter integer N_INP = 0;
	// Trace: design.sv:23327:13
	parameter integer LOG_N_INP = $clog2(N_INP);
	// Trace: design.sv:23329:3
	input wire [N_INP - 1:0] inp_data_i;
	// Trace: design.sv:23330:3
	input wire [N_INP - 1:0] inp_valid_i;
	// Trace: design.sv:23331:3
	output reg [N_INP - 1:0] inp_ready_o;
	// Trace: design.sv:23333:3
	input wire [LOG_N_INP - 1:0] inp_sel_i;
	// Trace: design.sv:23335:3
	output wire oup_data_o;
	// Trace: design.sv:23336:3
	output wire oup_valid_o;
	// Trace: design.sv:23337:3
	input wire oup_ready_i;
	// Trace: design.sv:23340:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:23341:5
		inp_ready_o = 1'sb0;
		// Trace: design.sv:23342:5
		inp_ready_o[inp_sel_i] = oup_ready_i;
	end
	// Trace: design.sv:23344:3
	assign oup_data_o = inp_data_i[inp_sel_i];
	// Trace: design.sv:23345:3
	assign oup_valid_o = inp_valid_i[inp_sel_i];
	initial _sv2v_0 = 0;
endmodule
module stream_throttle (
	clk_i,
	rst_ni,
	req_valid_i,
	req_valid_o,
	req_ready_i,
	req_ready_o,
	rsp_valid_i,
	rsp_ready_i,
	credit_i
);
	reg _sv2v_0;
	// Trace: design.sv:23370:15
	parameter [31:0] MaxNumPending = 1;
	// Trace: design.sv:23372:15
	function automatic [31:0] cf_math_pkg_idx_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:58:9
		cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	parameter [31:0] CntWidth = cf_math_pkg_idx_width(MaxNumPending);
	// Trace: design.sv:23374:20
	// removed localparam type credit_t
	// Trace: design.sv:23377:5
	input wire clk_i;
	// Trace: design.sv:23379:5
	input wire rst_ni;
	// Trace: design.sv:23382:5
	input wire req_valid_i;
	// Trace: design.sv:23384:5
	output wire req_valid_o;
	// Trace: design.sv:23386:5
	input wire req_ready_i;
	// Trace: design.sv:23388:5
	output wire req_ready_o;
	// Trace: design.sv:23391:5
	input wire rsp_valid_i;
	// Trace: design.sv:23393:5
	input wire rsp_ready_i;
	// Trace: design.sv:23396:5
	input wire [CntWidth - 1:0] credit_i;
	// Trace: design.sv:23401:5
	reg [CntWidth - 1:0] credit_d;
	reg [CntWidth - 1:0] credit_q;
	// Trace: design.sv:23404:5
	wire credit_available;
	// Trace: design.sv:23409:5
	always @(*) begin : proc_credit_counter
		if (_sv2v_0)
			;
		// Trace: design.sv:23412:9
		credit_d = credit_q;
		// Trace: design.sv:23415:9
		if (req_ready_o & req_valid_o)
			// Trace: design.sv:23416:13
			credit_d = credit_d + 'd1;
		if (rsp_valid_i & rsp_ready_i)
			// Trace: design.sv:23421:13
			credit_d = credit_d - 'd1;
	end
	// Trace: design.sv:23426:5
	assign credit_available = credit_q <= (credit_i - 'd1);
	// Trace: design.sv:23429:5
	assign req_valid_o = req_valid_i & credit_available;
	// Trace: design.sv:23432:5
	assign req_ready_o = req_ready_i & credit_available;
	// Trace: macro expansion of FF at design.sv:23435:47
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at design.sv:23435:135
		if (!rst_ni)
			// Trace: macro expansion of FF at design.sv:23435:223
			credit_q <= 1'sb0;
		else
			// Trace: macro expansion of FF at design.sv:23435:395
			credit_q <= credit_d;
	initial _sv2v_0 = 0;
endmodule
module sub_per_hash (
	data_i,
	hash_o,
	hash_onehot_o
);
	// Trace: design.sv:23477:13
	parameter [31:0] InpWidth = 32'd11;
	// Trace: design.sv:23478:13
	parameter [31:0] HashWidth = 32'd5;
	// Trace: design.sv:23479:13
	parameter [31:0] NoRounds = 32'd1;
	// Trace: design.sv:23480:13
	parameter [31:0] PermuteKey = 32'd299034753;
	// Trace: design.sv:23481:13
	parameter [31:0] XorKey = 32'd4094834;
	// Trace: design.sv:23484:3
	input wire [InpWidth - 1:0] data_i;
	// Trace: design.sv:23485:3
	output wire [HashWidth - 1:0] hash_o;
	// Trace: design.sv:23486:3
	output wire [(2 ** HashWidth) - 1:0] hash_onehot_o;
	// Trace: design.sv:23490:3
	// removed localparam type perm_lists_t
	// Trace: design.sv:23491:3
	wire [((NoRounds * InpWidth) * 32) - 1:0] Permutations;
	// Trace: design.sv:23492:3
	function automatic [((NoRounds * InpWidth) * 32) - 1:0] get_permutations;
		// Trace: design.sv:23534:52
		input reg [31:0] seed;
		// Trace: design.sv:23535:5
		reg [31:0] indices [0:NoRounds - 1][0:InpWidth - 1];
		// Trace: design.sv:23536:5
		reg [((NoRounds * InpWidth) * 32) - 1:0] perm_array;
		// Trace: design.sv:23537:5
		reg [63:0] A;
		// Trace: design.sv:23538:5
		reg [63:0] C;
		// Trace: design.sv:23539:5
		reg [63:0] M;
		// Trace: design.sv:23540:5
		reg [63:0] index;
		// Trace: design.sv:23541:5
		reg [63:0] advance;
		// Trace: design.sv:23542:5
		reg [63:0] rand_number;
		begin
			A = 2147483629;
			C = 2147483587;
			M = 33'sd2147483648 - 1;
			index = 0;
			advance = 0;
			rand_number = ((A * seed) + C) % M;
			// Trace: design.sv:23545:5
			begin : sv2v_autoblock_1
				// Trace: design.sv:23545:10
				reg [31:0] r;
				// Trace: design.sv:23545:10
				for (r = 0; r < NoRounds; r = r + 1)
					begin
						// Trace: design.sv:23547:7
						begin : sv2v_autoblock_2
							// Trace: design.sv:23547:12
							reg [31:0] i;
							// Trace: design.sv:23547:12
							for (i = 0; i < InpWidth; i = i + 1)
								begin
									// Trace: design.sv:23548:9
									indices[r][i] = i;
								end
						end
						begin : sv2v_autoblock_3
							// Trace: design.sv:23551:12
							reg [31:0] i;
							// Trace: design.sv:23551:12
							for (i = 0; i < InpWidth; i = i + 1)
								begin
									// Trace: design.sv:23553:9
									if (i > 0) begin
										// Trace: design.sv:23554:11
										rand_number = ((A * rand_number) + C) % M;
										// Trace: design.sv:23555:11
										index = rand_number % i;
									end
									if (i != index) begin
										// Trace: design.sv:23559:11
										perm_array[((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - i)) * 32+:32] = perm_array[((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - index)) * 32+:32];
										// Trace: design.sv:23560:11
										perm_array[((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - index)) * 32+:32] = indices[r][i];
									end
								end
						end
						// Trace: design.sv:23564:7
						rand_number = ((A * rand_number) + C) % M;
						// Trace: design.sv:23565:7
						advance = rand_number % NoRounds;
						begin : sv2v_autoblock_4
							// Trace: design.sv:23566:12
							reg [31:0] i;
							// Trace: design.sv:23566:12
							for (i = 0; i < advance; i = i + 1)
								begin
									// Trace: design.sv:23567:9
									rand_number = ((A * rand_number) + C) % M;
								end
						end
					end
			end
			get_permutations = perm_array;
		end
	endfunction
	assign Permutations = get_permutations(PermuteKey);
	// Trace: design.sv:23496:3
	// removed localparam type xor_stages_t
	// Trace: design.sv:23497:3
	wire [(((NoRounds * InpWidth) * 3) * 32) - 1:0] XorStages;
	// Trace: design.sv:23498:3
	function automatic [(((NoRounds * InpWidth) * 3) * 32) - 1:0] get_xor_stages;
		// Trace: design.sv:23579:50
		input reg [31:0] seed;
		// Trace: design.sv:23580:5
		reg [(((NoRounds * InpWidth) * 3) * 32) - 1:0] xor_array;
		// Trace: design.sv:23581:5
		reg [63:0] A;
		// Trace: design.sv:23582:5
		reg [63:0] C;
		// Trace: design.sv:23583:5
		reg [63:0] M;
		// Trace: design.sv:23584:5
		reg [63:0] index;
		// Trace: design.sv:23586:5
		reg [63:0] advance;
		// Trace: design.sv:23587:5
		reg [63:0] rand_number;
		begin
			A = 1664525;
			C = 1013904223;
			M = 34'sd4294967296;
			index = 0;
			advance = 0;
			rand_number = ((A * seed) + C) % M;
			// Trace: design.sv:23592:5
			begin : sv2v_autoblock_5
				// Trace: design.sv:23592:10
				reg [31:0] r;
				// Trace: design.sv:23592:10
				for (r = 0; r < NoRounds; r = r + 1)
					begin
						// Trace: design.sv:23594:7
						begin : sv2v_autoblock_6
							// Trace: design.sv:23594:12
							reg [31:0] i;
							// Trace: design.sv:23594:12
							for (i = 0; i < InpWidth; i = i + 1)
								begin
									// Trace: design.sv:23595:9
									rand_number = ((A * rand_number) + C) % M;
									// Trace: design.sv:23597:9
									begin : sv2v_autoblock_7
										// Trace: design.sv:23597:14
										reg [31:0] j;
										// Trace: design.sv:23597:14
										for (j = 0; j < 3; j = j + 1)
											begin
												// Trace: design.sv:23598:11
												rand_number = ((A * rand_number) + C) % M;
												// Trace: design.sv:23599:11
												index = rand_number % InpWidth;
												// Trace: design.sv:23600:11
												xor_array[((((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - i)) * 3) + (2 - j)) * 32+:32] = index;
											end
									end
								end
						end
						// Trace: design.sv:23604:7
						rand_number = ((A * rand_number) + C) % M;
						// Trace: design.sv:23605:7
						advance = rand_number % NoRounds;
						begin : sv2v_autoblock_8
							// Trace: design.sv:23606:12
							reg [31:0] i;
							// Trace: design.sv:23606:12
							for (i = 0; i < advance; i = i + 1)
								begin
									// Trace: design.sv:23607:9
									rand_number = ((A * rand_number) + C) % M;
								end
						end
					end
			end
			get_xor_stages = xor_array;
		end
	endfunction
	assign XorStages = get_xor_stages(XorKey);
	// Trace: design.sv:23501:3
	wire [(NoRounds * InpWidth) - 1:0] permuted;
	wire [(NoRounds * InpWidth) - 1:0] xored;
	// Trace: design.sv:23504:3
	genvar _gv_r_1;
	generate
		for (_gv_r_1 = 0; _gv_r_1 < NoRounds; _gv_r_1 = _gv_r_1 + 1) begin : gen_round
			localparam r = _gv_r_1;
			genvar _gv_i_12;
			for (_gv_i_12 = 0; _gv_i_12 < InpWidth; _gv_i_12 = _gv_i_12 + 1) begin : gen_sub_per
				localparam i = _gv_i_12;
				if (r == 0) begin : gen_input
					// Trace: design.sv:23510:9
					assign permuted[(r * InpWidth) + i] = data_i[Permutations[((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - i)) * 32+:32]];
				end
				else begin : gen_permutation
					// Trace: design.sv:23512:9
					assign permuted[(r * InpWidth) + i] = permuted[((r - 1) * InpWidth) + Permutations[((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - i)) * 32+:32]];
				end
				// Trace: design.sv:23516:7
				assign xored[(r * InpWidth) + i] = (permuted[(r * InpWidth) + XorStages[((((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - i)) * 3) + 2) * 32+:32]] ^ permuted[(r * InpWidth) + XorStages[((((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - i)) * 3) + 1) * 32+:32]]) ^ permuted[(r * InpWidth) + XorStages[(((((NoRounds - 1) - r) * InpWidth) + ((InpWidth - 1) - i)) * 3) * 32+:32]];
			end
		end
	endgenerate
	// Trace: design.sv:23523:3
	assign hash_o = xored[((NoRounds - 1) * InpWidth) + (HashWidth - 1)-:HashWidth];
	// Trace: design.sv:23525:3
	assign hash_onehot_o = 1 << hash_o;
	// Trace: design.sv:23534:3
	// Trace: design.sv:23579:3
endmodule
module sync (
	clk_i,
	rst_ni,
	serial_i,
	serial_o
);
	// Trace: design.sv:23626:15
	parameter [31:0] STAGES = 2;
	// Trace: design.sv:23627:15
	parameter [0:0] ResetValue = 1'b0;
	// Trace: design.sv:23629:5
	input wire clk_i;
	// Trace: design.sv:23630:5
	input wire rst_ni;
	// Trace: design.sv:23631:5
	input wire serial_i;
	// Trace: design.sv:23632:5
	output wire serial_o;
	// Trace: design.sv:23637:4
	reg [STAGES - 1:0] reg_q;
	// Trace: design.sv:23639:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:23640:9
		if (!rst_ni)
			// Trace: design.sv:23641:13
			reg_q <= {STAGES {ResetValue}};
		else
			// Trace: design.sv:23643:13
			reg_q <= {reg_q[STAGES - 2:0], serial_i};
	// Trace: design.sv:23647:5
	assign serial_o = reg_q[STAGES - 1];
endmodule
module sync_wedge (
	clk_i,
	rst_ni,
	en_i,
	serial_i,
	r_edge_o,
	f_edge_o,
	serial_o
);
	// Trace: design.sv:23663:15
	parameter [31:0] STAGES = 2;
	// Trace: design.sv:23665:5
	input wire clk_i;
	// Trace: design.sv:23666:5
	input wire rst_ni;
	// Trace: design.sv:23667:5
	input wire en_i;
	// Trace: design.sv:23668:5
	input wire serial_i;
	// Trace: design.sv:23669:5
	output wire r_edge_o;
	// Trace: design.sv:23670:5
	output wire f_edge_o;
	// Trace: design.sv:23671:5
	output wire serial_o;
	// Trace: design.sv:23673:5
	wire clk;
	// Trace: design.sv:23674:5
	wire serial;
	reg serial_q;
	// Trace: design.sv:23676:5
	assign serial_o = serial_q;
	// Trace: design.sv:23677:5
	assign f_edge_o = ~serial & serial_q;
	// Trace: design.sv:23678:5
	assign r_edge_o = serial & ~serial_q;
	// Trace: design.sv:23680:5
	sync #(.STAGES(STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(serial_i),
		.serial_o(serial)
	);
	// Trace: design.sv:23689:5
	pulp_clock_gating i_pulp_clock_gating(
		.clk_i(clk_i),
		.en_i(en_i),
		.test_en_i(1'b0),
		.clk_o(clk)
	);
	// Trace: design.sv:23696:5
	always @(posedge clk or negedge rst_ni)
		// Trace: design.sv:23697:9
		if (!rst_ni)
			// Trace: design.sv:23698:13
			serial_q <= 1'b0;
		else
			// Trace: design.sv:23700:13
			if (en_i)
				// Trace: design.sv:23701:17
				serial_q <= serial;
endmodule
module unread (d_i);
	// Trace: design.sv:23722:5
	input wire d_i;
endmodule
module read (
	d_i,
	d_o
);
	// Trace: design.sv:23737:15
	parameter [31:0] Width = 1;
	// Trace: design.sv:23738:20
	// removed localparam type T
	// Trace: design.sv:23740:5
	input wire [Width - 1:0] d_i;
	// Trace: design.sv:23741:5
	output wire [Width - 1:0] d_o;
	// Trace: design.sv:23744:3
	assign d_o = d_i;
endmodule
// removed package "cdc_reset_ctrlr_pkg"
module cdc_2phase_D7A8F_A47F6 (
	src_rst_ni,
	src_clk_i,
	src_data_i,
	src_valid_i,
	src_ready_o,
	dst_rst_ni,
	dst_clk_i,
	dst_data_o,
	dst_valid_o,
	dst_ready_i
);
	// removed localparam type T_PtrWidth_type
	parameter signed [31:0] T_PtrWidth = 0;
	// Trace: design.sv:23817:18
	// removed localparam type T
	// Trace: design.sv:23819:3
	input wire src_rst_ni;
	// Trace: design.sv:23820:3
	input wire src_clk_i;
	// Trace: design.sv:23821:3
	input wire [T_PtrWidth - 1:0] src_data_i;
	// Trace: design.sv:23822:3
	input wire src_valid_i;
	// Trace: design.sv:23823:3
	output wire src_ready_o;
	// Trace: design.sv:23825:3
	input wire dst_rst_ni;
	// Trace: design.sv:23826:3
	input wire dst_clk_i;
	// Trace: design.sv:23827:3
	output wire [T_PtrWidth - 1:0] dst_data_o;
	// Trace: design.sv:23828:3
	output wire dst_valid_o;
	// Trace: design.sv:23829:3
	input wire dst_ready_i;
	// Trace: design.sv:23833:4
	wire async_req;
	// Trace: design.sv:23834:4
	wire async_ack;
	// Trace: design.sv:23835:4
	wire [T_PtrWidth - 1:0] async_data;
	// Trace: design.sv:23838:3
	cdc_2phase_src_F2E4A_14906 #(.T_T_PtrWidth(T_PtrWidth)) i_src(
		.rst_ni(src_rst_ni),
		.clk_i(src_clk_i),
		.data_i(src_data_i),
		.valid_i(src_valid_i),
		.ready_o(src_ready_o),
		.async_req_o(async_req),
		.async_ack_i(async_ack),
		.async_data_o(async_data)
	);
	// Trace: design.sv:23850:3
	cdc_2phase_dst_ED4EB_75D31 #(.T_T_PtrWidth(T_PtrWidth)) i_dst(
		.rst_ni(dst_rst_ni),
		.clk_i(dst_clk_i),
		.data_o(dst_data_o),
		.valid_o(dst_valid_o),
		.ready_i(dst_ready_i),
		.async_req_i(async_req),
		.async_ack_o(async_ack),
		.async_data_i(async_data)
	);
endmodule
module cdc_2phase_src_F2E4A_14906 (
	rst_ni,
	clk_i,
	data_i,
	valid_i,
	ready_o,
	async_req_o,
	async_ack_i,
	async_data_o
);
	// removed localparam type T_T_PtrWidth_type
	parameter signed [31:0] T_T_PtrWidth = 0;
	// Trace: design.sv:23866:18
	// removed localparam type T
	// Trace: design.sv:23868:3
	input wire rst_ni;
	// Trace: design.sv:23869:3
	input wire clk_i;
	// Trace: design.sv:23870:3
	input wire [T_T_PtrWidth - 1:0] data_i;
	// Trace: design.sv:23871:3
	input wire valid_i;
	// Trace: design.sv:23872:3
	output wire ready_o;
	// Trace: design.sv:23873:3
	output wire async_req_o;
	// Trace: design.sv:23874:3
	input wire async_ack_i;
	// Trace: design.sv:23875:3
	output wire [T_T_PtrWidth - 1:0] async_data_o;
	// Trace: design.sv:23879:3
	reg req_src_q;
	reg ack_src_q;
	reg ack_q;
	// Trace: design.sv:23881:3
	reg [T_T_PtrWidth - 1:0] data_src_q;
	// Trace: design.sv:23884:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:23885:5
		if (!rst_ni) begin
			// Trace: design.sv:23886:7
			req_src_q <= 0;
			// Trace: design.sv:23887:7
			data_src_q <= 1'sb0;
		end
		else if (valid_i && ready_o) begin
			// Trace: design.sv:23889:7
			req_src_q <= ~req_src_q;
			// Trace: design.sv:23890:7
			data_src_q <= data_i;
		end
	// Trace: design.sv:23895:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:23896:5
		if (!rst_ni) begin
			// Trace: design.sv:23897:7
			ack_src_q <= 0;
			// Trace: design.sv:23898:7
			ack_q <= 0;
		end
		else begin
			// Trace: design.sv:23900:7
			ack_src_q <= async_ack_i;
			// Trace: design.sv:23901:7
			ack_q <= ack_src_q;
		end
	// Trace: design.sv:23906:3
	assign ready_o = req_src_q == ack_q;
	// Trace: design.sv:23907:3
	assign async_req_o = req_src_q;
	// Trace: design.sv:23908:3
	assign async_data_o = data_src_q;
endmodule
module cdc_2phase_dst_ED4EB_75D31 (
	rst_ni,
	clk_i,
	data_o,
	valid_o,
	ready_i,
	async_req_i,
	async_ack_o,
	async_data_i
);
	// removed localparam type T_T_PtrWidth_type
	parameter signed [31:0] T_T_PtrWidth = 0;
	// Trace: design.sv:23916:18
	// removed localparam type T
	// Trace: design.sv:23918:3
	input wire rst_ni;
	// Trace: design.sv:23919:3
	input wire clk_i;
	// Trace: design.sv:23920:3
	output wire [T_T_PtrWidth - 1:0] data_o;
	// Trace: design.sv:23921:3
	output wire valid_o;
	// Trace: design.sv:23922:3
	input wire ready_i;
	// Trace: design.sv:23923:3
	input wire async_req_i;
	// Trace: design.sv:23924:3
	output wire async_ack_o;
	// Trace: design.sv:23925:3
	input wire [T_T_PtrWidth - 1:0] async_data_i;
	// Trace: design.sv:23930:3
	reg req_dst_q;
	reg req_q0;
	reg req_q1;
	reg ack_dst_q;
	// Trace: design.sv:23932:3
	reg [T_T_PtrWidth - 1:0] data_dst_q;
	// Trace: design.sv:23935:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:23936:5
		if (!rst_ni)
			// Trace: design.sv:23937:7
			ack_dst_q <= 0;
		else if (valid_o && ready_i)
			// Trace: design.sv:23939:7
			ack_dst_q <= ~ack_dst_q;
	// Trace: design.sv:23945:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:23946:5
		if (!rst_ni)
			// Trace: design.sv:23947:7
			data_dst_q <= 1'sb0;
		else if ((req_q0 != req_q1) && !valid_o)
			// Trace: design.sv:23949:7
			data_dst_q <= async_data_i;
	// Trace: design.sv:23954:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:23955:5
		if (!rst_ni) begin
			// Trace: design.sv:23956:7
			req_dst_q <= 0;
			// Trace: design.sv:23957:7
			req_q0 <= 0;
			// Trace: design.sv:23958:7
			req_q1 <= 0;
		end
		else begin
			// Trace: design.sv:23960:7
			req_dst_q <= async_req_i;
			// Trace: design.sv:23961:7
			req_q0 <= req_dst_q;
			// Trace: design.sv:23962:7
			req_q1 <= req_q0;
		end
	// Trace: design.sv:23967:3
	assign valid_o = ack_dst_q != req_q1;
	// Trace: design.sv:23968:3
	assign data_o = data_dst_q;
	// Trace: design.sv:23969:3
	assign async_ack_o = ack_dst_q;
endmodule
module cdc_4phase (
	src_rst_ni,
	src_clk_i,
	src_data_i,
	src_valid_i,
	src_ready_o,
	dst_rst_ni,
	dst_clk_i,
	dst_data_o,
	dst_valid_o,
	dst_ready_i
);
	// Trace: design.sv:24009:18
	// removed localparam type T
	// Trace: design.sv:24010:13
	parameter [0:0] DECOUPLED = 1'b1;
	// Trace: design.sv:24011:13
	parameter [0:0] SEND_RESET_MSG = 1'b0;
	// Trace: design.sv:24012:13
	parameter [0:0] RESET_MSG = 1'b0;
	// Trace: design.sv:24014:3
	input wire src_rst_ni;
	// Trace: design.sv:24015:3
	input wire src_clk_i;
	// Trace: design.sv:24016:3
	input wire src_data_i;
	// Trace: design.sv:24017:3
	input wire src_valid_i;
	// Trace: design.sv:24018:3
	output wire src_ready_o;
	// Trace: design.sv:24020:3
	input wire dst_rst_ni;
	// Trace: design.sv:24021:3
	input wire dst_clk_i;
	// Trace: design.sv:24022:3
	output wire dst_data_o;
	// Trace: design.sv:24023:3
	output wire dst_valid_o;
	// Trace: design.sv:24024:3
	input wire dst_ready_i;
	// Trace: design.sv:24028:4
	wire async_req;
	// Trace: design.sv:24029:4
	wire async_ack;
	// Trace: design.sv:24030:4
	wire async_data;
	// Trace: design.sv:24033:3
	cdc_4phase_src_48DA8 #(
		.DECOUPLED(DECOUPLED),
		.SEND_RESET_MSG(SEND_RESET_MSG),
		.RESET_MSG(RESET_MSG)
	) i_src(
		.rst_ni(src_rst_ni),
		.clk_i(src_clk_i),
		.data_i(src_data_i),
		.valid_i(src_valid_i),
		.ready_o(src_ready_o),
		.async_req_o(async_req),
		.async_ack_i(async_ack),
		.async_data_o(async_data)
	);
	// Trace: design.sv:24050:3
	cdc_4phase_dst_D4479 #(.DECOUPLED(DECOUPLED)) i_dst(
		.rst_ni(dst_rst_ni),
		.clk_i(dst_clk_i),
		.data_o(dst_data_o),
		.valid_o(dst_valid_o),
		.ready_i(dst_ready_i),
		.async_req_i(async_req),
		.async_ack_o(async_ack),
		.async_data_i(async_data)
	);
endmodule
module cdc_4phase_src_DFE1F (
	rst_ni,
	clk_i,
	data_i,
	valid_i,
	ready_o,
	async_req_o,
	async_ack_i,
	async_data_o
);
	reg _sv2v_0;
	// Trace: design.sv:24065:18
	// removed localparam type T
	// Trace: design.sv:24066:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:24067:13
	parameter [0:0] DECOUPLED = 1'b1;
	// Trace: design.sv:24068:13
	parameter [0:0] SEND_RESET_MSG = 1'b0;
	// Trace: design.sv:24069:13
	parameter [1:0] RESET_MSG = 2'b00;
	// Trace: design.sv:24071:3
	input wire rst_ni;
	// Trace: design.sv:24072:3
	input wire clk_i;
	// Trace: design.sv:24073:3
	input wire [1:0] data_i;
	// Trace: design.sv:24074:3
	input wire valid_i;
	// Trace: design.sv:24075:3
	output reg ready_o;
	// Trace: design.sv:24076:3
	output wire async_req_o;
	// Trace: design.sv:24077:3
	input wire async_ack_i;
	// Trace: design.sv:24078:3
	output wire [1:0] async_data_o;
	// Trace: design.sv:24082:3
	reg req_src_d;
	reg req_src_q;
	// Trace: design.sv:24084:3
	reg [1:0] data_src_d;
	reg [1:0] data_src_q;
	// Trace: design.sv:24086:3
	wire ack_synced;
	// Trace: design.sv:24088:3
	// removed localparam type state_e
	// Trace: design.sv:24089:3
	reg [1:0] state_d;
	reg [1:0] state_q;
	// Trace: design.sv:24092:3
	sync #(.STAGES(SYNC_STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(async_ack_i),
		.serial_o(ack_synced)
	);
	// Trace: design.sv:24102:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:24103:5
		state_d = state_q;
		// Trace: design.sv:24104:5
		req_src_d = 1'b0;
		// Trace: design.sv:24105:5
		data_src_d = data_src_q;
		// Trace: design.sv:24106:5
		ready_o = 1'b0;
		// Trace: design.sv:24107:5
		case (state_q)
			2'd0: begin
				// Trace: design.sv:24111:9
				if (DECOUPLED)
					// Trace: design.sv:24112:11
					ready_o = 1'b1;
				else
					// Trace: design.sv:24114:11
					ready_o = 1'b0;
				if (valid_i) begin
					// Trace: design.sv:24118:11
					data_src_d = data_i;
					// Trace: design.sv:24119:11
					req_src_d = 1'b1;
					// Trace: design.sv:24120:11
					state_d = 2'd1;
				end
			end
			2'd1: begin
				// Trace: design.sv:24124:9
				req_src_d = 1'b1;
				// Trace: design.sv:24125:9
				if (ack_synced == 1'b1) begin
					// Trace: design.sv:24126:11
					req_src_d = 1'b0;
					// Trace: design.sv:24127:11
					state_d = 2'd2;
				end
			end
			2'd2:
				// Trace: design.sv:24131:9
				if (ack_synced == 1'b0) begin
					// Trace: design.sv:24132:11
					state_d = 2'd0;
					// Trace: design.sv:24133:11
					if (!DECOUPLED)
						// Trace: design.sv:24134:13
						ready_o = 1'b1;
				end
			default:
				// Trace: design.sv:24139:9
				state_d = 2'd0;
		endcase
	end
	// Trace: design.sv:24144:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:24145:5
		if (!rst_ni)
			// Trace: design.sv:24146:7
			state_q <= 2'd0;
		else
			// Trace: design.sv:24148:7
			state_q <= state_d;
	// Trace: design.sv:24153:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:24154:5
		if (!rst_ni) begin
			begin
				// Trace: design.sv:24155:7
				if (SEND_RESET_MSG) begin
					// Trace: design.sv:24156:9
					req_src_q <= 1'b1;
					// Trace: design.sv:24157:9
					data_src_q <= RESET_MSG;
				end
				else begin
					// Trace: design.sv:24159:9
					req_src_q <= 1'b0;
					// Trace: design.sv:24160:9
					data_src_q <= 2'b00;
				end
			end
		end
		else begin
			// Trace: design.sv:24163:7
			req_src_q <= req_src_d;
			// Trace: design.sv:24164:7
			data_src_q <= data_src_d;
		end
	// Trace: design.sv:24169:3
	assign async_req_o = req_src_q;
	// Trace: design.sv:24170:3
	assign async_data_o = data_src_q;
	initial _sv2v_0 = 0;
endmodule
module cdc_4phase_src_48DA8 (
	rst_ni,
	clk_i,
	data_i,
	valid_i,
	ready_o,
	async_req_o,
	async_ack_i,
	async_data_o
);
	reg _sv2v_0;
	// Trace: design.sv:24065:18
	// removed localparam type T
	// Trace: design.sv:24066:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:24067:13
	parameter [0:0] DECOUPLED = 1'b1;
	// Trace: design.sv:24068:13
	parameter [0:0] SEND_RESET_MSG = 1'b0;
	// Trace: design.sv:24069:13
	parameter [0:0] RESET_MSG = 1'b0;
	// Trace: design.sv:24071:3
	input wire rst_ni;
	// Trace: design.sv:24072:3
	input wire clk_i;
	// Trace: design.sv:24073:3
	input wire data_i;
	// Trace: design.sv:24074:3
	input wire valid_i;
	// Trace: design.sv:24075:3
	output reg ready_o;
	// Trace: design.sv:24076:3
	output wire async_req_o;
	// Trace: design.sv:24077:3
	input wire async_ack_i;
	// Trace: design.sv:24078:3
	output wire async_data_o;
	// Trace: design.sv:24082:3
	reg req_src_d;
	reg req_src_q;
	// Trace: design.sv:24084:3
	reg data_src_d;
	reg data_src_q;
	// Trace: design.sv:24086:3
	wire ack_synced;
	// Trace: design.sv:24088:3
	// removed localparam type state_e
	// Trace: design.sv:24089:3
	reg [1:0] state_d;
	reg [1:0] state_q;
	// Trace: design.sv:24092:3
	sync #(.STAGES(SYNC_STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(async_ack_i),
		.serial_o(ack_synced)
	);
	// Trace: design.sv:24102:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:24103:5
		state_d = state_q;
		// Trace: design.sv:24104:5
		req_src_d = 1'b0;
		// Trace: design.sv:24105:5
		data_src_d = data_src_q;
		// Trace: design.sv:24106:5
		ready_o = 1'b0;
		// Trace: design.sv:24107:5
		case (state_q)
			2'd0: begin
				// Trace: design.sv:24111:9
				if (DECOUPLED)
					// Trace: design.sv:24112:11
					ready_o = 1'b1;
				else
					// Trace: design.sv:24114:11
					ready_o = 1'b0;
				if (valid_i) begin
					// Trace: design.sv:24118:11
					data_src_d = data_i;
					// Trace: design.sv:24119:11
					req_src_d = 1'b1;
					// Trace: design.sv:24120:11
					state_d = 2'd1;
				end
			end
			2'd1: begin
				// Trace: design.sv:24124:9
				req_src_d = 1'b1;
				// Trace: design.sv:24125:9
				if (ack_synced == 1'b1) begin
					// Trace: design.sv:24126:11
					req_src_d = 1'b0;
					// Trace: design.sv:24127:11
					state_d = 2'd2;
				end
			end
			2'd2:
				// Trace: design.sv:24131:9
				if (ack_synced == 1'b0) begin
					// Trace: design.sv:24132:11
					state_d = 2'd0;
					// Trace: design.sv:24133:11
					if (!DECOUPLED)
						// Trace: design.sv:24134:13
						ready_o = 1'b1;
				end
			default:
				// Trace: design.sv:24139:9
				state_d = 2'd0;
		endcase
	end
	// Trace: design.sv:24144:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:24145:5
		if (!rst_ni)
			// Trace: design.sv:24146:7
			state_q <= 2'd0;
		else
			// Trace: design.sv:24148:7
			state_q <= state_d;
	// Trace: design.sv:24153:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:24154:5
		if (!rst_ni) begin
			begin
				// Trace: design.sv:24155:7
				if (SEND_RESET_MSG) begin
					// Trace: design.sv:24156:9
					req_src_q <= 1'b1;
					// Trace: design.sv:24157:9
					data_src_q <= RESET_MSG;
				end
				else begin
					// Trace: design.sv:24159:9
					req_src_q <= 1'b0;
					// Trace: design.sv:24160:9
					data_src_q <= 1'b0;
				end
			end
		end
		else begin
			// Trace: design.sv:24163:7
			req_src_q <= req_src_d;
			// Trace: design.sv:24164:7
			data_src_q <= data_src_d;
		end
	// Trace: design.sv:24169:3
	assign async_req_o = req_src_q;
	// Trace: design.sv:24170:3
	assign async_data_o = data_src_q;
	initial _sv2v_0 = 0;
endmodule
module cdc_4phase_dst_A46CE (
	rst_ni,
	clk_i,
	data_o,
	valid_o,
	ready_i,
	async_req_i,
	async_ack_o,
	async_data_i
);
	reg _sv2v_0;
	// Trace: design.sv:24178:18
	// removed localparam type T
	// Trace: design.sv:24179:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:24180:13
	parameter [0:0] DECOUPLED = 1;
	// Trace: design.sv:24182:3
	input wire rst_ni;
	// Trace: design.sv:24183:3
	input wire clk_i;
	// Trace: design.sv:24184:3
	output wire [1:0] data_o;
	// Trace: design.sv:24185:3
	output wire valid_o;
	// Trace: design.sv:24186:3
	input wire ready_i;
	// Trace: design.sv:24187:3
	input wire async_req_i;
	// Trace: design.sv:24188:3
	output wire async_ack_o;
	// Trace: design.sv:24189:3
	input wire [1:0] async_data_i;
	// Trace: design.sv:24193:3
	reg ack_dst_d;
	reg ack_dst_q;
	// Trace: design.sv:24195:3
	wire req_synced;
	// Trace: design.sv:24197:3
	reg data_valid;
	// Trace: design.sv:24199:3
	wire output_ready;
	// Trace: design.sv:24202:3
	// removed localparam type state_e
	// Trace: design.sv:24203:3
	reg [1:0] state_d;
	reg [1:0] state_q;
	// Trace: design.sv:24206:3
	sync #(.STAGES(SYNC_STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(async_req_i),
		.serial_o(req_synced)
	);
	// Trace: design.sv:24216:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:24217:5
		state_d = state_q;
		// Trace: design.sv:24218:5
		data_valid = 1'b0;
		// Trace: design.sv:24219:5
		ack_dst_d = 1'b0;
		// Trace: design.sv:24221:5
		case (state_q)
			2'd0:
				// Trace: design.sv:24224:9
				if (req_synced == 1'b1) begin
					// Trace: design.sv:24225:11
					data_valid = 1'b1;
					// Trace: design.sv:24226:11
					if (output_ready == 1'b1)
						// Trace: design.sv:24227:13
						state_d = 2'd2;
					else
						// Trace: design.sv:24229:13
						state_d = 2'd1;
				end
			2'd1: begin
				// Trace: design.sv:24235:9
				data_valid = 1'b1;
				// Trace: design.sv:24236:9
				if (output_ready == 1'b1) begin
					// Trace: design.sv:24237:11
					state_d = 2'd2;
					// Trace: design.sv:24238:11
					ack_dst_d = 1'b1;
				end
			end
			2'd2: begin
				// Trace: design.sv:24243:9
				ack_dst_d = 1'b1;
				// Trace: design.sv:24244:9
				if (req_synced == 1'b0) begin
					// Trace: design.sv:24245:11
					ack_dst_d = 1'b0;
					// Trace: design.sv:24246:11
					state_d = 2'd0;
				end
			end
			default:
				// Trace: design.sv:24251:9
				state_d = 2'd0;
		endcase
	end
	// Trace: design.sv:24256:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:24257:5
		if (!rst_ni)
			// Trace: design.sv:24258:7
			state_q <= 2'd0;
		else
			// Trace: design.sv:24260:7
			state_q <= state_d;
	// Trace: design.sv:24265:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:24266:5
		if (!rst_ni)
			// Trace: design.sv:24267:7
			ack_dst_q <= 1'b0;
		else
			// Trace: design.sv:24269:7
			ack_dst_q <= ack_dst_d;
	// Trace: design.sv:24273:3
	generate
		if (DECOUPLED) begin : gen_decoupled
			// Trace: design.sv:24276:5
			spill_register_8294E #(.Bypass(1'b0)) i_spill_register(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.valid_i(data_valid),
				.ready_o(output_ready),
				.data_i(async_data_i),
				.valid_o(valid_o),
				.ready_i(ready_i),
				.data_o(data_o)
			);
		end
		else begin : gen_not_decoupled
			// Trace: design.sv:24290:5
			assign valid_o = data_valid;
			// Trace: design.sv:24291:5
			assign output_ready = ready_i;
			// Trace: design.sv:24292:5
			assign data_o = async_data_i;
		end
	endgenerate
	// Trace: design.sv:24296:3
	assign async_ack_o = ack_dst_q;
	initial _sv2v_0 = 0;
endmodule
module cdc_4phase_dst_D4479 (
	rst_ni,
	clk_i,
	data_o,
	valid_o,
	ready_i,
	async_req_i,
	async_ack_o,
	async_data_i
);
	reg _sv2v_0;
	// Trace: design.sv:24178:18
	// removed localparam type T
	// Trace: design.sv:24179:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:24180:13
	parameter [0:0] DECOUPLED = 1;
	// Trace: design.sv:24182:3
	input wire rst_ni;
	// Trace: design.sv:24183:3
	input wire clk_i;
	// Trace: design.sv:24184:3
	output wire data_o;
	// Trace: design.sv:24185:3
	output wire valid_o;
	// Trace: design.sv:24186:3
	input wire ready_i;
	// Trace: design.sv:24187:3
	input wire async_req_i;
	// Trace: design.sv:24188:3
	output wire async_ack_o;
	// Trace: design.sv:24189:3
	input wire async_data_i;
	// Trace: design.sv:24193:3
	reg ack_dst_d;
	reg ack_dst_q;
	// Trace: design.sv:24195:3
	wire req_synced;
	// Trace: design.sv:24197:3
	reg data_valid;
	// Trace: design.sv:24199:3
	wire output_ready;
	// Trace: design.sv:24202:3
	// removed localparam type state_e
	// Trace: design.sv:24203:3
	reg [1:0] state_d;
	reg [1:0] state_q;
	// Trace: design.sv:24206:3
	sync #(.STAGES(SYNC_STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(async_req_i),
		.serial_o(req_synced)
	);
	// Trace: design.sv:24216:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:24217:5
		state_d = state_q;
		// Trace: design.sv:24218:5
		data_valid = 1'b0;
		// Trace: design.sv:24219:5
		ack_dst_d = 1'b0;
		// Trace: design.sv:24221:5
		case (state_q)
			2'd0:
				// Trace: design.sv:24224:9
				if (req_synced == 1'b1) begin
					// Trace: design.sv:24225:11
					data_valid = 1'b1;
					// Trace: design.sv:24226:11
					if (output_ready == 1'b1)
						// Trace: design.sv:24227:13
						state_d = 2'd2;
					else
						// Trace: design.sv:24229:13
						state_d = 2'd1;
				end
			2'd1: begin
				// Trace: design.sv:24235:9
				data_valid = 1'b1;
				// Trace: design.sv:24236:9
				if (output_ready == 1'b1) begin
					// Trace: design.sv:24237:11
					state_d = 2'd2;
					// Trace: design.sv:24238:11
					ack_dst_d = 1'b1;
				end
			end
			2'd2: begin
				// Trace: design.sv:24243:9
				ack_dst_d = 1'b1;
				// Trace: design.sv:24244:9
				if (req_synced == 1'b0) begin
					// Trace: design.sv:24245:11
					ack_dst_d = 1'b0;
					// Trace: design.sv:24246:11
					state_d = 2'd0;
				end
			end
			default:
				// Trace: design.sv:24251:9
				state_d = 2'd0;
		endcase
	end
	// Trace: design.sv:24256:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:24257:5
		if (!rst_ni)
			// Trace: design.sv:24258:7
			state_q <= 2'd0;
		else
			// Trace: design.sv:24260:7
			state_q <= state_d;
	// Trace: design.sv:24265:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:24266:5
		if (!rst_ni)
			// Trace: design.sv:24267:7
			ack_dst_q <= 1'b0;
		else
			// Trace: design.sv:24269:7
			ack_dst_q <= ack_dst_d;
	// Trace: design.sv:24273:3
	generate
		if (DECOUPLED) begin : gen_decoupled
			// Trace: design.sv:24276:5
			spill_register_736F9 #(.Bypass(1'b0)) i_spill_register(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.valid_i(data_valid),
				.ready_o(output_ready),
				.data_i(async_data_i),
				.valid_o(valid_o),
				.ready_i(ready_i),
				.data_o(data_o)
			);
		end
		else begin : gen_not_decoupled
			// Trace: design.sv:24290:5
			assign valid_o = data_valid;
			// Trace: design.sv:24291:5
			assign output_ready = ready_i;
			// Trace: design.sv:24292:5
			assign data_o = async_data_i;
		end
	endgenerate
	// Trace: design.sv:24296:3
	assign async_ack_o = ack_dst_q;
	initial _sv2v_0 = 0;
endmodule
module addr_decode_6EF7A (
	addr_i,
	addr_map_i,
	idx_o,
	dec_valid_o,
	dec_error_o,
	en_default_idx_i,
	default_idx_i
);
	reg _sv2v_0;
	// Trace: design.sv:24334:13
	parameter [31:0] NoIndices = 32'd0;
	// Trace: design.sv:24336:13
	parameter [31:0] NoRules = 32'd0;
	// Trace: design.sv:24338:26
	// removed localparam type addr_t
	// Trace: design.sv:24356:26
	// removed localparam type rule_t
	// Trace: design.sv:24358:13
	parameter [0:0] Napot = 0;
	// Trace: design.sv:24362:13
	function automatic [31:0] cf_math_pkg_idx_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:58:9
		cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	parameter [31:0] IdxWidth = cf_math_pkg_idx_width(NoIndices);
	// Trace: design.sv:24366:26
	// removed localparam type idx_t
	// Trace: design.sv:24369:3
	input wire [31:0] addr_i;
	// Trace: design.sv:24371:3
	input wire [(NoRules * 96) - 1:0] addr_map_i;
	// Trace: design.sv:24373:3
	output reg [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:24375:3
	output reg dec_valid_o;
	// Trace: design.sv:24377:3
	output reg dec_error_o;
	// Trace: design.sv:24381:3
	input wire en_default_idx_i;
	// Trace: design.sv:24387:3
	input wire [IdxWidth - 1:0] default_idx_i;
	// Trace: design.sv:24390:3
	reg [NoRules - 1:0] matched_rules;
	// Trace: design.sv:24392:3
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:24394:5
		matched_rules = 1'sb0;
		// Trace: design.sv:24395:5
		dec_valid_o = 1'b0;
		// Trace: design.sv:24396:5
		dec_error_o = (en_default_idx_i ? 1'b0 : 1'b1);
		// Trace: design.sv:24397:5
		idx_o = (en_default_idx_i ? default_idx_i : {IdxWidth {1'sb0}});
		// Trace: design.sv:24400:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:24400:10
			reg [31:0] i;
			// Trace: design.sv:24400:10
			for (i = 0; i < NoRules; i = i + 1)
				begin
					// Trace: design.sv:24401:7
					if (((!Napot && (addr_i >= addr_map_i[(i * 96) + 63-:32])) && ((addr_i < addr_map_i[(i * 96) + 31-:32]) || (addr_map_i[(i * 96) + 31-:32] == {32 {1'sb0}}))) || (Napot && ((addr_map_i[(i * 96) + 63-:32] & addr_map_i[(i * 96) + 31-:32]) == (addr_i & addr_map_i[(i * 96) + 31-:32])))) begin
						// Trace: design.sv:24407:9
						matched_rules[i] = 1'b1;
						// Trace: design.sv:24408:9
						dec_valid_o = 1'b1;
						// Trace: design.sv:24409:9
						dec_error_o = 1'b0;
						// Trace: design.sv:24410:9
						idx_o = sv2v_cast_5FDFE(addr_map_i[(i * 96) + 95-:32]);
					end
				end
		end
	end
	initial _sv2v_0 = 0;
endmodule
module addr_decode_133FF (
	addr_i,
	addr_map_i,
	idx_o,
	dec_valid_o,
	dec_error_o,
	en_default_idx_i,
	default_idx_i
);
	reg _sv2v_0;
	// Trace: design.sv:24334:13
	parameter [31:0] NoIndices = 32'd0;
	// Trace: design.sv:24336:13
	parameter [31:0] NoRules = 32'd0;
	// Trace: design.sv:24338:26
	// removed localparam type addr_t
	// Trace: design.sv:24356:26
	// removed localparam type rule_t
	// Trace: design.sv:24358:13
	parameter [0:0] Napot = 0;
	// Trace: design.sv:24362:13
	function automatic [31:0] cf_math_pkg_idx_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:58:9
		cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	parameter [31:0] IdxWidth = cf_math_pkg_idx_width(NoIndices);
	// Trace: design.sv:24366:26
	// removed localparam type idx_t
	// Trace: design.sv:24369:3
	input wire addr_i;
	// Trace: design.sv:24371:3
	input wire [(NoRules * 34) - 1:0] addr_map_i;
	// Trace: design.sv:24373:3
	output reg [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:24375:3
	output reg dec_valid_o;
	// Trace: design.sv:24377:3
	output reg dec_error_o;
	// Trace: design.sv:24381:3
	input wire en_default_idx_i;
	// Trace: design.sv:24387:3
	input wire [IdxWidth - 1:0] default_idx_i;
	// Trace: design.sv:24390:3
	reg [NoRules - 1:0] matched_rules;
	// Trace: design.sv:24392:3
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:24394:5
		matched_rules = 1'sb0;
		// Trace: design.sv:24395:5
		dec_valid_o = 1'b0;
		// Trace: design.sv:24396:5
		dec_error_o = (en_default_idx_i ? 1'b0 : 1'b1);
		// Trace: design.sv:24397:5
		idx_o = (en_default_idx_i ? default_idx_i : {IdxWidth {1'sb0}});
		// Trace: design.sv:24400:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:24400:10
			reg [31:0] i;
			// Trace: design.sv:24400:10
			for (i = 0; i < NoRules; i = i + 1)
				begin
					// Trace: design.sv:24401:7
					if (((!Napot && (addr_i >= addr_map_i[(i * 34) + 1])) && ((addr_i < addr_map_i[i * 34]) || (addr_map_i[i * 34] == 1'b0))) || (Napot && ((addr_map_i[(i * 34) + 1] & addr_map_i[i * 34]) == (addr_i & addr_map_i[i * 34])))) begin
						// Trace: design.sv:24407:9
						matched_rules[i] = 1'b1;
						// Trace: design.sv:24408:9
						dec_valid_o = 1'b1;
						// Trace: design.sv:24409:9
						dec_error_o = 1'b0;
						// Trace: design.sv:24410:9
						idx_o = sv2v_cast_5FDFE(addr_map_i[(i * 34) + 33-:32]);
					end
				end
		end
	end
	initial _sv2v_0 = 0;
endmodule
module addr_decode_napot (
	addr_i,
	addr_map_i,
	idx_o,
	dec_valid_o,
	dec_error_o,
	en_default_idx_i,
	default_idx_i
);
	// Trace: design.sv:24500:13
	parameter [31:0] NoIndices = 32'd0;
	// Trace: design.sv:24502:13
	parameter [31:0] NoRules = 32'd0;
	// Trace: design.sv:24504:26
	// removed localparam type addr_t
	// Trace: design.sv:24517:26
	// removed localparam type rule_t
	// Trace: design.sv:24521:13
	function automatic [31:0] cf_math_pkg_idx_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:58:9
		cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	parameter [31:0] IdxWidth = cf_math_pkg_idx_width(NoIndices);
	// Trace: design.sv:24525:26
	// removed localparam type idx_t
	// Trace: design.sv:24528:3
	input wire addr_i;
	// Trace: design.sv:24530:3
	input wire [NoRules - 1:0] addr_map_i;
	// Trace: design.sv:24532:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: design.sv:24534:3
	output wire dec_valid_o;
	// Trace: design.sv:24536:3
	output wire dec_error_o;
	// Trace: design.sv:24540:3
	input wire en_default_idx_i;
	// Trace: design.sv:24546:3
	input wire [IdxWidth - 1:0] default_idx_i;
	// Trace: design.sv:24550:3
	// removed localparam type rule_range_t
	// Trace: design.sv:24556:3
	addr_decode_133FF #(
		.NoIndices(NoIndices),
		.NoRules(NoRules),
		.Napot(1)
	) i_addr_decode(
		.addr_i(addr_i),
		.addr_map_i(addr_map_i),
		.idx_o(idx_o),
		.dec_valid_o(dec_valid_o),
		.dec_error_o(dec_error_o),
		.en_default_idx_i(en_default_idx_i),
		.default_idx_i(default_idx_i)
	);
endmodule
module cb_filter (
	clk_i,
	rst_ni,
	look_data_i,
	look_valid_o,
	incr_data_i,
	incr_valid_i,
	decr_data_i,
	decr_valid_i,
	filter_clear_i,
	filter_usage_o,
	filter_full_o,
	filter_empty_o,
	filter_error_o
);
	reg _sv2v_0;
	// Trace: design.sv:24616:13
	parameter [31:0] KHashes = 32'd3;
	// Trace: design.sv:24617:13
	parameter [31:0] HashWidth = 32'd4;
	// Trace: design.sv:24618:13
	parameter [31:0] HashRounds = 32'd1;
	// Trace: design.sv:24619:13
	parameter [31:0] InpWidth = 32'd32;
	// Trace: design.sv:24620:13
	parameter [31:0] BucketWidth = 32'd4;
	// Trace: design.sv:24622:13
	// removed localparam type cb_filter_pkg_cb_seed_t
	localparam [191:0] cb_filter_pkg_EgSeeds = 192'h11d2e881003e7b72012ff886000f318100047df403e20e8f;
	parameter [(KHashes * 64) - 1:0] Seeds = cb_filter_pkg_EgSeeds;
	// Trace: design.sv:24624:3
	input wire clk_i;
	// Trace: design.sv:24625:3
	input wire rst_ni;
	// Trace: design.sv:24627:3
	input wire [InpWidth - 1:0] look_data_i;
	// Trace: design.sv:24628:3
	output wire look_valid_o;
	// Trace: design.sv:24630:3
	input wire [InpWidth - 1:0] incr_data_i;
	// Trace: design.sv:24631:3
	input wire incr_valid_i;
	// Trace: design.sv:24633:3
	input wire [InpWidth - 1:0] decr_data_i;
	// Trace: design.sv:24634:3
	input wire decr_valid_i;
	// Trace: design.sv:24636:3
	input wire filter_clear_i;
	// Trace: design.sv:24637:3
	output wire [HashWidth - 1:0] filter_usage_o;
	// Trace: design.sv:24638:3
	output wire filter_full_o;
	// Trace: design.sv:24639:3
	output wire filter_empty_o;
	// Trace: design.sv:24640:3
	output wire filter_error_o;
	// Trace: design.sv:24643:3
	localparam [31:0] NoCounters = 2 ** HashWidth;
	// Trace: design.sv:24646:3
	wire [NoCounters - 1:0] look_ind;
	// Trace: design.sv:24647:3
	wire [NoCounters - 1:0] incr_ind;
	// Trace: design.sv:24648:3
	wire [NoCounters - 1:0] decr_ind;
	// Trace: design.sv:24650:3
	reg [NoCounters - 1:0] bucket_en;
	// Trace: design.sv:24651:3
	wire [NoCounters - 1:0] bucket_down;
	// Trace: design.sv:24652:3
	wire [NoCounters - 1:0] bucket_occupied;
	// Trace: design.sv:24653:3
	wire [NoCounters - 1:0] bucket_overflow;
	// Trace: design.sv:24654:3
	wire [NoCounters - 1:0] bucket_full;
	// Trace: design.sv:24655:3
	wire [NoCounters - 1:0] bucket_empty;
	// Trace: design.sv:24657:3
	wire [NoCounters - 1:0] data_in_bucket;
	// Trace: design.sv:24659:3
	wire cnt_en;
	// Trace: design.sv:24660:3
	wire cnt_down;
	// Trace: design.sv:24661:3
	wire cnt_overflow;
	// Trace: design.sv:24666:3
	hash_block #(
		.NoHashes(KHashes),
		.InpWidth(InpWidth),
		.HashWidth(HashWidth),
		.NoRounds(HashRounds),
		.Seeds(Seeds)
	) i_look_hashes(
		.data_i(look_data_i),
		.indicator_o(look_ind)
	);
	// Trace: design.sv:24676:3
	assign data_in_bucket = look_ind & bucket_occupied;
	// Trace: design.sv:24677:3
	assign look_valid_o = (data_in_bucket == look_ind ? 1'b1 : 1'b0);
	// Trace: design.sv:24682:3
	hash_block #(
		.NoHashes(KHashes),
		.InpWidth(InpWidth),
		.HashWidth(HashWidth),
		.NoRounds(HashRounds),
		.Seeds(Seeds)
	) i_incr_hashes(
		.data_i(incr_data_i),
		.indicator_o(incr_ind)
	);
	// Trace: design.sv:24696:3
	hash_block #(
		.NoHashes(KHashes),
		.InpWidth(InpWidth),
		.HashWidth(HashWidth),
		.NoRounds(HashRounds),
		.Seeds(Seeds)
	) i_decr_hashes(
		.data_i(decr_data_i),
		.indicator_o(decr_ind)
	);
	// Trace: design.sv:24710:3
	assign bucket_down = (decr_valid_i ? decr_ind : {NoCounters {1'sb0}});
	// Trace: design.sv:24712:3
	always @(*) begin : proc_bucket_control
		if (_sv2v_0)
			;
		// Trace: design.sv:24713:5
		case ({incr_valid_i, decr_valid_i})
			2'b00:
				// Trace: design.sv:24714:15
				bucket_en = 1'sb0;
			2'b10:
				// Trace: design.sv:24715:15
				bucket_en = incr_ind;
			2'b01:
				// Trace: design.sv:24716:15
				bucket_en = decr_ind;
			2'b11:
				// Trace: design.sv:24717:15
				bucket_en = incr_ind ^ decr_ind;
			default:
				// Trace: design.sv:24718:16
				bucket_en = 1'sb0;
		endcase
	end
	// Trace: design.sv:24725:3
	genvar _gv_i_13;
	generate
		for (_gv_i_13 = 0; _gv_i_13 < NoCounters; _gv_i_13 = _gv_i_13 + 1) begin : gen_buckets
			localparam i = _gv_i_13;
			// Trace: design.sv:24726:5
			wire [BucketWidth - 1:0] bucket_content;
			// Trace: design.sv:24727:5
			// removed localparam type sv2v_uu_i_bucket_load_i
			localparam [0:0] sv2v_uu_i_bucket_ext_load_i_0 = 1'sb0;
			localparam [31:0] sv2v_uu_i_bucket_WIDTH = BucketWidth;
			// removed localparam type sv2v_uu_i_bucket_d_i
			localparam [BucketWidth - 1:0] sv2v_uu_i_bucket_ext_d_i_0 = 1'sb0;
			counter #(.WIDTH(BucketWidth)) i_bucket(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.clear_i(filter_clear_i),
				.en_i(bucket_en[i]),
				.load_i(sv2v_uu_i_bucket_ext_load_i_0),
				.down_i(bucket_down[i]),
				.d_i(sv2v_uu_i_bucket_ext_d_i_0),
				.q_o(bucket_content),
				.overflow_o(bucket_overflow[i])
			);
			// Trace: design.sv:24740:5
			assign bucket_full[i] = bucket_overflow[i] | &bucket_content;
			// Trace: design.sv:24741:5
			assign bucket_occupied[i] = |bucket_content;
			// Trace: design.sv:24742:5
			assign bucket_empty[i] = ~bucket_occupied[i];
		end
	endgenerate
	// Trace: design.sv:24748:3
	assign cnt_en = incr_valid_i ^ decr_valid_i;
	// Trace: design.sv:24749:3
	assign cnt_down = decr_valid_i;
	// Trace: design.sv:24750:3
	// removed localparam type sv2v_uu_i_tot_count_load_i
	localparam [0:0] sv2v_uu_i_tot_count_ext_load_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_tot_count_WIDTH = HashWidth;
	// removed localparam type sv2v_uu_i_tot_count_d_i
	localparam [sv2v_uu_i_tot_count_WIDTH - 1:0] sv2v_uu_i_tot_count_ext_d_i_0 = 1'sb0;
	counter #(.WIDTH(HashWidth)) i_tot_count(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clear_i(filter_clear_i),
		.en_i(cnt_en),
		.load_i(sv2v_uu_i_tot_count_ext_load_i_0),
		.down_i(cnt_down),
		.d_i(sv2v_uu_i_tot_count_ext_d_i_0),
		.q_o(filter_usage_o),
		.overflow_o(cnt_overflow)
	);
	// Trace: design.sv:24767:3
	assign filter_full_o = |bucket_full;
	// Trace: design.sv:24768:3
	assign filter_empty_o = &bucket_empty;
	// Trace: design.sv:24769:3
	assign filter_error_o = |bucket_overflow | cnt_overflow;
	initial _sv2v_0 = 0;
endmodule
module hash_block (
	data_i,
	indicator_o
);
	reg _sv2v_0;
	// Trace: design.sv:24774:13
	parameter [31:0] NoHashes = 32'd3;
	// Trace: design.sv:24775:13
	parameter [31:0] InpWidth = 32'd11;
	// Trace: design.sv:24776:13
	parameter [31:0] HashWidth = 32'd5;
	// Trace: design.sv:24777:13
	parameter [31:0] NoRounds = 32'd1;
	// Trace: design.sv:24778:13
	// removed localparam type cb_filter_pkg_cb_seed_t
	localparam [191:0] cb_filter_pkg_EgSeeds = 192'h11d2e881003e7b72012ff886000f318100047df403e20e8f;
	parameter [(NoHashes * 64) - 1:0] Seeds = cb_filter_pkg_EgSeeds;
	// Trace: design.sv:24780:3
	input wire [InpWidth - 1:0] data_i;
	// Trace: design.sv:24781:3
	output reg [(2 ** HashWidth) - 1:0] indicator_o;
	// Trace: design.sv:24784:3
	wire [(NoHashes * (2 ** HashWidth)) - 1:0] hashes;
	// Trace: design.sv:24786:3
	genvar _gv_i_14;
	generate
		for (_gv_i_14 = 0; _gv_i_14 < NoHashes; _gv_i_14 = _gv_i_14 + 1) begin : gen_hashes
			localparam i = _gv_i_14;
			// Trace: design.sv:24787:5
			sub_per_hash #(
				.InpWidth(InpWidth),
				.HashWidth(HashWidth),
				.NoRounds(NoRounds),
				.PermuteKey(Seeds[(i * 64) + 63-:32]),
				.XorKey(Seeds[(i * 64) + 31-:32])
			) i_hash(
				.data_i(data_i),
				.hash_o(),
				.hash_onehot_o(hashes[i * (2 ** HashWidth)+:2 ** HashWidth])
			);
		end
	endgenerate
	// Trace: design.sv:24801:3
	always @(*) begin : proc_hash_or
		if (_sv2v_0)
			;
		// Trace: design.sv:24802:5
		indicator_o = 1'sb0;
		// Trace: design.sv:24803:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:24803:10
			reg [31:0] i;
			// Trace: design.sv:24803:10
			for (i = 0; i < (2 ** HashWidth); i = i + 1)
				begin
					// Trace: design.sv:24804:7
					begin : sv2v_autoblock_2
						// Trace: design.sv:24804:12
						reg [31:0] j;
						// Trace: design.sv:24804:12
						for (j = 0; j < NoHashes; j = j + 1)
							begin
								// Trace: design.sv:24805:9
								indicator_o[i] = indicator_o[i] | hashes[(j * (2 ** HashWidth)) + i];
							end
					end
				end
		end
	end
	initial _sv2v_0 = 0;
endmodule
module cdc_fifo_2phase (
	src_rst_ni,
	src_clk_i,
	src_data_i,
	src_valid_i,
	src_ready_o,
	dst_rst_ni,
	dst_clk_i,
	dst_data_o,
	dst_valid_o,
	dst_ready_i
);
	// Trace: design.sv:24867:18
	// removed localparam type T
	// Trace: design.sv:24869:13
	parameter signed [31:0] LOG_DEPTH = 3;
	// Trace: design.sv:24871:3
	input wire src_rst_ni;
	// Trace: design.sv:24872:3
	input wire src_clk_i;
	// Trace: design.sv:24873:3
	input wire src_data_i;
	// Trace: design.sv:24874:3
	input wire src_valid_i;
	// Trace: design.sv:24875:3
	output wire src_ready_o;
	// Trace: design.sv:24877:3
	input wire dst_rst_ni;
	// Trace: design.sv:24878:3
	input wire dst_clk_i;
	// Trace: design.sv:24879:3
	output wire dst_data_o;
	// Trace: design.sv:24880:3
	output wire dst_valid_o;
	// Trace: design.sv:24881:3
	input wire dst_ready_i;
	// Trace: design.sv:24886:3
	initial begin
		// Trace: design.sv:24887:5
		assert (LOG_DEPTH > 0) ;
	end
	// Trace: design.sv:24891:3
	localparam signed [31:0] PtrWidth = LOG_DEPTH + 1;
	// Trace: design.sv:24892:3
	// removed localparam type pointer_t
	// Trace: design.sv:24893:3
	// removed localparam type index_t
	// Trace: design.sv:24895:3
	localparam [PtrWidth - 1:0] PtrFull = 1 << LOG_DEPTH;
	// Trace: design.sv:24896:3
	localparam [PtrWidth - 1:0] PtrEmpty = 1'sb0;
	// Trace: design.sv:24903:3
	wire [LOG_DEPTH - 1:0] fifo_widx;
	wire [LOG_DEPTH - 1:0] fifo_ridx;
	// Trace: design.sv:24904:3
	wire fifo_write;
	// Trace: design.sv:24905:3
	wire fifo_wdata;
	wire fifo_rdata;
	// Trace: design.sv:24906:3
	reg fifo_data_q [0:(2 ** LOG_DEPTH) - 1];
	// Trace: design.sv:24908:3
	assign fifo_rdata = fifo_data_q[fifo_ridx];
	// Trace: design.sv:24910:3
	genvar _gv_i_15;
	generate
		for (_gv_i_15 = 0; _gv_i_15 < (2 ** LOG_DEPTH); _gv_i_15 = _gv_i_15 + 1) begin : g_word
			localparam i = _gv_i_15;
			// Trace: design.sv:24911:5
			always @(posedge src_clk_i or negedge src_rst_ni)
				// Trace: design.sv:24912:7
				if (!src_rst_ni)
					// Trace: design.sv:24913:9
					fifo_data_q[i] <= 1'sb0;
				else if (fifo_write && (fifo_widx == i))
					// Trace: design.sv:24915:9
					fifo_data_q[i] <= fifo_wdata;
		end
	endgenerate
	// Trace: design.sv:24920:3
	reg [PtrWidth - 1:0] src_wptr_q;
	wire [PtrWidth - 1:0] dst_wptr;
	wire [PtrWidth - 1:0] src_rptr;
	reg [PtrWidth - 1:0] dst_rptr_q;
	// Trace: design.sv:24922:3
	always @(posedge src_clk_i or negedge src_rst_ni)
		// Trace: design.sv:24923:5
		if (!src_rst_ni)
			// Trace: design.sv:24924:7
			src_wptr_q <= 0;
		else if (src_valid_i && src_ready_o)
			// Trace: design.sv:24926:7
			src_wptr_q <= src_wptr_q + 1;
	// Trace: design.sv:24929:3
	always @(posedge dst_clk_i or negedge dst_rst_ni)
		// Trace: design.sv:24930:5
		if (!dst_rst_ni)
			// Trace: design.sv:24931:7
			dst_rptr_q <= 0;
		else if (dst_valid_o && dst_ready_i)
			// Trace: design.sv:24933:7
			dst_rptr_q <= dst_rptr_q + 1;
	// Trace: design.sv:24940:3
	assign src_ready_o = (src_wptr_q ^ src_rptr) != PtrFull;
	// Trace: design.sv:24941:3
	assign dst_valid_o = (dst_rptr_q ^ dst_wptr) != PtrEmpty;
	// Trace: design.sv:24944:3
	cdc_2phase_D7A8F_A47F6 #(.T_PtrWidth(PtrWidth)) i_cdc_wptr(
		.src_rst_ni(src_rst_ni),
		.src_clk_i(src_clk_i),
		.src_data_i(src_wptr_q),
		.src_valid_i(1'b1),
		.src_ready_o(),
		.dst_rst_ni(dst_rst_ni),
		.dst_clk_i(dst_clk_i),
		.dst_data_o(dst_wptr),
		.dst_valid_o(),
		.dst_ready_i(1'b1)
	);
	// Trace: design.sv:24957:3
	cdc_2phase_D7A8F_A47F6 #(.T_PtrWidth(PtrWidth)) i_cdc_rptr(
		.src_rst_ni(dst_rst_ni),
		.src_clk_i(dst_clk_i),
		.src_data_i(dst_rptr_q),
		.src_valid_i(1'b1),
		.src_ready_o(),
		.dst_rst_ni(src_rst_ni),
		.dst_clk_i(src_clk_i),
		.dst_data_o(src_rptr),
		.dst_valid_o(),
		.dst_ready_i(1'b1)
	);
	// Trace: design.sv:24971:3
	assign fifo_widx = src_wptr_q;
	// Trace: design.sv:24972:3
	assign fifo_wdata = src_data_i;
	// Trace: design.sv:24973:3
	assign fifo_write = src_valid_i && src_ready_o;
	// Trace: design.sv:24974:3
	assign fifo_ridx = dst_rptr_q;
	// Trace: design.sv:24975:3
	assign dst_data_o = fifo_rdata;
endmodule
module counter (
	clk_i,
	rst_ni,
	clear_i,
	en_i,
	load_i,
	down_i,
	d_i,
	q_o,
	overflow_o
);
	// Trace: design.sv:24992:15
	parameter [31:0] WIDTH = 4;
	// Trace: design.sv:24993:15
	parameter [0:0] STICKY_OVERFLOW = 1'b0;
	// Trace: design.sv:24995:5
	input wire clk_i;
	// Trace: design.sv:24996:5
	input wire rst_ni;
	// Trace: design.sv:24997:5
	input wire clear_i;
	// Trace: design.sv:24998:5
	input wire en_i;
	// Trace: design.sv:24999:5
	input wire load_i;
	// Trace: design.sv:25000:5
	input wire down_i;
	// Trace: design.sv:25001:5
	input wire [WIDTH - 1:0] d_i;
	// Trace: design.sv:25002:5
	output wire [WIDTH - 1:0] q_o;
	// Trace: design.sv:25003:5
	output wire overflow_o;
	// Trace: design.sv:25005:5
	delta_counter #(
		.WIDTH(WIDTH),
		.STICKY_OVERFLOW(STICKY_OVERFLOW)
	) i_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clear_i(clear_i),
		.en_i(en_i),
		.load_i(load_i),
		.down_i(down_i),
		.delta_i({{WIDTH - 1 {1'b0}}, 1'b1}),
		.d_i(d_i),
		.q_o(q_o),
		.overflow_o(overflow_o)
	);
endmodule
module ecc_decode (
	data_i,
	data_o,
	syndrome_o,
	single_error_o,
	parity_error_o,
	double_error_o
);
	reg _sv2v_0;
	// removed import ecc_pkg::*;
	// Trace: design.sv:25051:14
	parameter [31:0] DataWidth = 64;
	// Trace: design.sv:25053:18
	// removed localparam type data_t
	// Trace: design.sv:25054:18
	function automatic [31:0] ecc_pkg_get_parity_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:18:53
		input reg [31:0] data_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:20:5
		reg [31:0] cw_width;
		begin
			cw_width = 2;
			// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:21:5
			while ($unsigned(2 ** cw_width) < ((cw_width + data_width) + 1)) begin
				// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:21:64
				cw_width = cw_width + 1;
			end
			ecc_pkg_get_parity_width = cw_width;
		end
	endfunction
	// removed localparam type parity_t
	// Trace: design.sv:25055:18
	function automatic [31:0] ecc_pkg_get_cw_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:26:49
		input reg [31:0] data_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:28:5
		ecc_pkg_get_cw_width = data_width + ecc_pkg_get_parity_width(data_width);
	endfunction
	// removed localparam type code_word_t
	// Trace: design.sv:25056:18
	// removed localparam type encoded_data_t
	// Trace: design.sv:25062:3
	input wire [(1 + ecc_pkg_get_cw_width(DataWidth)) - 1:0] data_i;
	// Trace: design.sv:25064:3
	output wire [DataWidth - 1:0] data_o;
	// Trace: design.sv:25066:3
	output wire [ecc_pkg_get_parity_width(DataWidth) - 1:0] syndrome_o;
	// Trace: design.sv:25068:3
	output wire single_error_o;
	// Trace: design.sv:25070:3
	output wire parity_error_o;
	// Trace: design.sv:25072:3
	output wire double_error_o;
	// Trace: design.sv:25075:3
	wire parity;
	// Trace: design.sv:25076:3
	reg [DataWidth - 1:0] data_wo_parity;
	// Trace: design.sv:25077:3
	reg [ecc_pkg_get_parity_width(DataWidth) - 1:0] syndrome;
	// Trace: design.sv:25078:3
	wire syndrome_not_zero;
	// Trace: design.sv:25079:3
	reg [ecc_pkg_get_cw_width(DataWidth) - 1:0] correct_data;
	// Trace: design.sv:25082:3
	assign parity = data_i[ecc_pkg_get_cw_width(DataWidth) + 0] ^ ^data_i[ecc_pkg_get_cw_width(DataWidth) - 1-:ecc_pkg_get_cw_width(DataWidth)];
	// Trace: design.sv:25102:3
	always @(*) begin : calculate_syndrome
		if (_sv2v_0)
			;
		// Trace: design.sv:25103:5
		syndrome = 0;
		// Trace: design.sv:25104:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:25104:10
			reg [31:0] i;
			// Trace: design.sv:25104:10
			for (i = 0; i < $unsigned(ecc_pkg_get_parity_width(DataWidth)); i = i + 1)
				begin
					// Trace: design.sv:25105:7
					begin : sv2v_autoblock_2
						// Trace: design.sv:25105:12
						reg [31:0] j;
						// Trace: design.sv:25105:12
						for (j = 0; j < $unsigned(ecc_pkg_get_cw_width(DataWidth)); j = j + 1)
							begin
								// Trace: design.sv:25106:9
								if (|($unsigned(2 ** i) & (j + 1)))
									// Trace: design.sv:25106:43
									syndrome[i] = syndrome[i] ^ data_i[(ecc_pkg_get_cw_width(DataWidth) - 1) - ((ecc_pkg_get_cw_width(DataWidth) - 1) - j)];
							end
					end
				end
		end
	end
	// Trace: design.sv:25111:3
	assign syndrome_not_zero = |syndrome;
	// Trace: design.sv:25114:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:25115:5
		correct_data = data_i[ecc_pkg_get_cw_width(DataWidth) - 1-:ecc_pkg_get_cw_width(DataWidth)];
		// Trace: design.sv:25116:5
		if (syndrome_not_zero)
			// Trace: design.sv:25117:7
			correct_data[syndrome - 1] = ~data_i[(ecc_pkg_get_cw_width(DataWidth) - 1) - ((ecc_pkg_get_cw_width(DataWidth) - 1) - (syndrome - 1))];
	end
	// Trace: design.sv:25127:3
	assign single_error_o = parity & syndrome_not_zero;
	// Trace: design.sv:25128:3
	assign parity_error_o = parity & ~syndrome_not_zero;
	// Trace: design.sv:25129:3
	assign double_error_o = ~parity & syndrome_not_zero;
	// Trace: design.sv:25132:3
	always @(*) begin : sv2v_autoblock_3
		// Trace: design.sv:25133:5
		reg [31:0] idx;
		if (_sv2v_0)
			;
		// Trace: design.sv:25134:5
		data_wo_parity = 1'sb0;
		// Trace: design.sv:25135:5
		idx = 0;
		// Trace: design.sv:25137:5
		begin : sv2v_autoblock_4
			// Trace: design.sv:25137:10
			reg [31:0] i;
			// Trace: design.sv:25137:10
			for (i = 1; i < ($unsigned(ecc_pkg_get_cw_width(DataWidth)) + 1); i = i + 1)
				begin
					// Trace: design.sv:25139:7
					if ($unsigned(2 ** $clog2(i)) != i) begin
						// Trace: design.sv:25140:9
						data_wo_parity[idx] = correct_data[i - 1];
						// Trace: design.sv:25141:9
						idx = idx + 1;
					end
				end
		end
	end
	// Trace: design.sv:25146:3
	assign data_o = data_wo_parity;
	initial _sv2v_0 = 0;
endmodule
module ecc_encode (
	data_i,
	data_o
);
	reg _sv2v_0;
	// removed import ecc_pkg::*;
	// Trace: design.sv:25172:14
	parameter [31:0] DataWidth = 64;
	// Trace: design.sv:25174:18
	// removed localparam type data_t
	// Trace: design.sv:25175:18
	function automatic [31:0] ecc_pkg_get_parity_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:18:53
		input reg [31:0] data_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:20:5
		reg [31:0] cw_width;
		begin
			cw_width = 2;
			// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:21:5
			while ($unsigned(2 ** cw_width) < ((cw_width + data_width) + 1)) begin
				// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:21:64
				cw_width = cw_width + 1;
			end
			ecc_pkg_get_parity_width = cw_width;
		end
	endfunction
	// removed localparam type parity_t
	// Trace: design.sv:25176:18
	function automatic [31:0] ecc_pkg_get_cw_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:26:49
		input reg [31:0] data_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/ecc_pkg.sv:28:5
		ecc_pkg_get_cw_width = data_width + ecc_pkg_get_parity_width(data_width);
	endfunction
	// removed localparam type code_word_t
	// Trace: design.sv:25177:18
	// removed localparam type encoded_data_t
	// Trace: design.sv:25183:3
	input wire [DataWidth - 1:0] data_i;
	// Trace: design.sv:25185:3
	output wire [(1 + ecc_pkg_get_cw_width(DataWidth)) - 1:0] data_o;
	// Trace: design.sv:25188:3
	reg [ecc_pkg_get_parity_width(DataWidth) - 1:0] parity_code_word;
	// Trace: design.sv:25189:3
	reg [ecc_pkg_get_cw_width(DataWidth) - 1:0] data;
	reg [ecc_pkg_get_cw_width(DataWidth) - 1:0] codeword;
	// Trace: design.sv:25192:3
	always @(*) begin : expand_data
		// Trace: design.sv:25193:5
		reg [31:0] idx;
		if (_sv2v_0)
			;
		// Trace: design.sv:25194:5
		data = 1'sb0;
		// Trace: design.sv:25195:5
		idx = 0;
		// Trace: design.sv:25196:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:25196:10
			reg [31:0] i;
			// Trace: design.sv:25196:10
			for (i = 1; i < ($unsigned(ecc_pkg_get_cw_width(DataWidth)) + 1); i = i + 1)
				begin
					// Trace: design.sv:25198:7
					if ($unsigned(2 ** $clog2(i)) != i) begin
						// Trace: design.sv:25199:9
						data[i - 1] = data_i[idx];
						// Trace: design.sv:25200:9
						idx = idx + 1;
					end
				end
		end
	end
	// Trace: design.sv:25206:3
	always @(*) begin : calculate_syndrome
		if (_sv2v_0)
			;
		// Trace: design.sv:25207:5
		parity_code_word = 0;
		// Trace: design.sv:25208:5
		begin : sv2v_autoblock_2
			// Trace: design.sv:25208:10
			reg [31:0] i;
			// Trace: design.sv:25208:10
			for (i = 0; i < $unsigned(ecc_pkg_get_parity_width(DataWidth)); i = i + 1)
				begin
					// Trace: design.sv:25209:7
					begin : sv2v_autoblock_3
						// Trace: design.sv:25209:12
						reg [31:0] j;
						// Trace: design.sv:25209:12
						for (j = 1; j < ($unsigned(ecc_pkg_get_cw_width(DataWidth)) + 1); j = j + 1)
							begin
								// Trace: design.sv:25210:9
								if (|($unsigned(2 ** i) & j))
									// Trace: design.sv:25210:37
									parity_code_word[i] = parity_code_word[i] ^ data[j - 1];
							end
					end
				end
		end
	end
	// Trace: design.sv:25216:3
	always @(*) begin : generate_codeword
		if (_sv2v_0)
			;
		// Trace: design.sv:25217:7
		codeword = data;
		// Trace: design.sv:25218:7
		begin : sv2v_autoblock_4
			// Trace: design.sv:25218:12
			reg [31:0] i;
			// Trace: design.sv:25218:12
			for (i = 0; i < $unsigned(ecc_pkg_get_parity_width(DataWidth)); i = i + 1)
				begin
					// Trace: design.sv:25219:9
					codeword[(2 ** i) - 1] = parity_code_word[i];
				end
		end
	end
	// Trace: design.sv:25223:3
	assign data_o[ecc_pkg_get_cw_width(DataWidth) - 1-:ecc_pkg_get_cw_width(DataWidth)] = codeword;
	// Trace: design.sv:25224:3
	assign data_o[ecc_pkg_get_cw_width(DataWidth) + 0] = ^codeword;
	initial _sv2v_0 = 0;
endmodule
module edge_detect (
	clk_i,
	rst_ni,
	d_i,
	re_o,
	fe_o
);
	// Trace: design.sv:25241:5
	input wire clk_i;
	// Trace: design.sv:25242:5
	input wire rst_ni;
	// Trace: design.sv:25243:5
	input wire d_i;
	// Trace: design.sv:25244:5
	output wire re_o;
	// Trace: design.sv:25245:5
	output wire fe_o;
	// Trace: design.sv:25248:5
	sync_wedge i_sync_wedge(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.en_i(1'b1),
		.serial_i(d_i),
		.r_edge_o(re_o),
		.f_edge_o(fe_o),
		.serial_o()
	);
endmodule
module lzc (
	in_i,
	cnt_o,
	empty_o
);
	reg _sv2v_0;
	// Trace: design.sv:25275:13
	parameter [31:0] WIDTH = 2;
	// Trace: design.sv:25277:13
	parameter [0:0] MODE = 1'b0;
	// Trace: design.sv:25281:13
	function automatic [31:0] cf_math_pkg_idx_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:58:9
		cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	parameter [31:0] CNT_WIDTH = cf_math_pkg_idx_width(WIDTH);
	// Trace: design.sv:25284:3
	input wire [WIDTH - 1:0] in_i;
	// Trace: design.sv:25286:3
	output wire [CNT_WIDTH - 1:0] cnt_o;
	// Trace: design.sv:25288:3
	output wire empty_o;
	// Trace: design.sv:25291:3
	generate
		if (WIDTH == 1) begin : gen_degenerate_lzc
			// Trace: design.sv:25293:5
			assign cnt_o[0] = !in_i[0];
			// Trace: design.sv:25294:5
			assign empty_o = !in_i[0];
		end
		else begin : gen_lzc
			// Trace: design.sv:25298:5
			localparam [31:0] NumLevels = $clog2(WIDTH);
			// Trace: design.sv:25308:5
			wire [(WIDTH * NumLevels) - 1:0] index_lut;
			// Trace: design.sv:25309:5
			wire [(2 ** NumLevels) - 1:0] sel_nodes;
			// Trace: design.sv:25310:5
			wire [((2 ** NumLevels) * NumLevels) - 1:0] index_nodes;
			// Trace: design.sv:25312:5
			reg [WIDTH - 1:0] in_tmp;
			// Trace: design.sv:25315:5
			always @(*) begin : flip_vector
				if (_sv2v_0)
					;
				// Trace: design.sv:25316:7
				begin : sv2v_autoblock_1
					// Trace: design.sv:25316:12
					reg [31:0] i;
					// Trace: design.sv:25316:12
					for (i = 0; i < WIDTH; i = i + 1)
						begin
							// Trace: design.sv:25317:9
							in_tmp[i] = (MODE ? in_i[(WIDTH - 1) - i] : in_i[i]);
						end
				end
			end
			genvar _gv_j_7;
			for (_gv_j_7 = 0; $unsigned(_gv_j_7) < WIDTH; _gv_j_7 = _gv_j_7 + 1) begin : g_index_lut
				localparam j = _gv_j_7;
				// Trace: design.sv:25322:7
				function automatic [NumLevels - 1:0] sv2v_cast_677FF;
					input reg [NumLevels - 1:0] inp;
					sv2v_cast_677FF = inp;
				endfunction
				assign index_lut[j * NumLevels+:NumLevels] = sv2v_cast_677FF($unsigned(j));
			end
			genvar _gv_level_3;
			for (_gv_level_3 = 0; $unsigned(_gv_level_3) < NumLevels; _gv_level_3 = _gv_level_3 + 1) begin : g_levels
				localparam level = _gv_level_3;
				if ($unsigned(level) == (NumLevels - 1)) begin : g_last_level
					genvar _gv_k_6;
					for (_gv_k_6 = 0; _gv_k_6 < (2 ** level); _gv_k_6 = _gv_k_6 + 1) begin : g_level
						localparam k = _gv_k_6;
						if (($unsigned(k) * 2) < (WIDTH - 1)) begin : g_reduce
							// Trace: design.sv:25330:13
							assign sel_nodes[((2 ** level) - 1) + k] = in_tmp[k * 2] | in_tmp[(k * 2) + 1];
							// Trace: design.sv:25331:13
							assign index_nodes[(((2 ** level) - 1) + k) * NumLevels+:NumLevels] = (in_tmp[k * 2] == 1'b1 ? index_lut[(k * 2) * NumLevels+:NumLevels] : index_lut[((k * 2) + 1) * NumLevels+:NumLevels]);
						end
						if (($unsigned(k) * 2) == (WIDTH - 1)) begin : g_base
							// Trace: design.sv:25337:13
							assign sel_nodes[((2 ** level) - 1) + k] = in_tmp[k * 2];
							// Trace: design.sv:25338:13
							assign index_nodes[(((2 ** level) - 1) + k) * NumLevels+:NumLevels] = index_lut[(k * 2) * NumLevels+:NumLevels];
						end
						if (($unsigned(k) * 2) > (WIDTH - 1)) begin : g_out_of_range
							// Trace: design.sv:25342:13
							assign sel_nodes[((2 ** level) - 1) + k] = 1'b0;
							// Trace: design.sv:25343:13
							assign index_nodes[(((2 ** level) - 1) + k) * NumLevels+:NumLevels] = 1'sb0;
						end
					end
				end
				else begin : g_not_last_level
					genvar _gv_l_5;
					for (_gv_l_5 = 0; _gv_l_5 < (2 ** level); _gv_l_5 = _gv_l_5 + 1) begin : g_level
						localparam l = _gv_l_5;
						// Trace: design.sv:25348:11
						assign sel_nodes[((2 ** level) - 1) + l] = sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] | sel_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) + 1];
						// Trace: design.sv:25350:11
						assign index_nodes[(((2 ** level) - 1) + l) * NumLevels+:NumLevels] = (sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] == 1'b1 ? index_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) * NumLevels+:NumLevels] : index_nodes[((((2 ** (level + 1)) - 1) + (l * 2)) + 1) * NumLevels+:NumLevels]);
					end
				end
			end
			// Trace: design.sv:25357:5
			assign cnt_o = (NumLevels > $unsigned(0) ? index_nodes[0+:NumLevels] : {$clog2(WIDTH) {1'b0}});
			// Trace: design.sv:25358:5
			assign empty_o = (NumLevels > $unsigned(0) ? ~sel_nodes[0] : ~(|in_i));
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module max_counter (
	clk_i,
	rst_ni,
	clear_i,
	clear_max_i,
	en_i,
	load_i,
	down_i,
	delta_i,
	d_i,
	q_o,
	max_o,
	overflow_o,
	overflow_max_o
);
	reg _sv2v_0;
	// Trace: design.sv:25385:15
	parameter [31:0] WIDTH = 4;
	// Trace: design.sv:25387:5
	input wire clk_i;
	// Trace: design.sv:25388:5
	input wire rst_ni;
	// Trace: design.sv:25389:5
	input wire clear_i;
	// Trace: design.sv:25390:5
	input wire clear_max_i;
	// Trace: design.sv:25391:5
	input wire en_i;
	// Trace: design.sv:25392:5
	input wire load_i;
	// Trace: design.sv:25393:5
	input wire down_i;
	// Trace: design.sv:25394:5
	input wire [WIDTH - 1:0] delta_i;
	// Trace: design.sv:25395:5
	input wire [WIDTH - 1:0] d_i;
	// Trace: design.sv:25396:5
	output wire [WIDTH - 1:0] q_o;
	// Trace: design.sv:25397:5
	output reg [WIDTH - 1:0] max_o;
	// Trace: design.sv:25398:5
	output wire overflow_o;
	// Trace: design.sv:25399:5
	output wire overflow_max_o;
	// Trace: design.sv:25401:5
	reg [WIDTH - 1:0] max_d;
	reg [WIDTH - 1:0] max_q;
	// Trace: design.sv:25402:5
	reg overflow_max_d;
	reg overflow_max_q;
	// Trace: design.sv:25404:5
	delta_counter #(
		.WIDTH(WIDTH),
		.STICKY_OVERFLOW(1'b1)
	) i_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clear_i(clear_i),
		.en_i(en_i),
		.load_i(load_i),
		.down_i(down_i),
		.delta_i(delta_i),
		.d_i(d_i),
		.q_o(q_o),
		.overflow_o(overflow_o)
	);
	// Trace: design.sv:25420:5
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:25421:9
		max_d = max_q;
		// Trace: design.sv:25422:9
		max_o = max_q;
		// Trace: design.sv:25423:9
		overflow_max_d = overflow_max_q;
		// Trace: design.sv:25424:9
		if (clear_max_i) begin
			// Trace: design.sv:25425:13
			max_d = 1'sb0;
			// Trace: design.sv:25426:13
			overflow_max_d = 1'b0;
		end
		else if (q_o > max_q) begin
			// Trace: design.sv:25428:13
			max_d = q_o;
			// Trace: design.sv:25429:13
			max_o = q_o;
			// Trace: design.sv:25430:13
			if (overflow_o)
				// Trace: design.sv:25431:17
				overflow_max_d = 1'b1;
		end
	end
	// Trace: design.sv:25436:5
	assign overflow_max_o = overflow_max_q;
	// Trace: design.sv:25438:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:25439:9
		if (!rst_ni) begin
			// Trace: design.sv:25440:12
			max_q <= 1'sb0;
			// Trace: design.sv:25441:12
			overflow_max_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:25443:12
			max_q <= max_d;
			// Trace: design.sv:25444:12
			overflow_max_q <= overflow_max_d;
		end
	initial _sv2v_0 = 0;
endmodule
module rstgen (
	clk_i,
	rst_ni,
	test_mode_i,
	rst_no,
	init_no
);
	// Trace: design.sv:25462:5
	input wire clk_i;
	// Trace: design.sv:25463:5
	input wire rst_ni;
	// Trace: design.sv:25464:5
	input wire test_mode_i;
	// Trace: design.sv:25465:5
	output wire rst_no;
	// Trace: design.sv:25466:5
	output wire init_no;
	// Trace: design.sv:25469:5
	rstgen_bypass i_rstgen_bypass(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_test_mode_ni(rst_ni),
		.test_mode_i(test_mode_i),
		.rst_no(rst_no),
		.init_no(init_no)
	);
endmodule
module spill_register_0D540_46F20 (
	clk_i,
	rst_ni,
	valid_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// removed localparam type T_IdxWidth_type
	// removed localparam type T_payload_t_DataWidth_type
	// removed localparam type T_payload_t_IdxWidth_type
	// removed localparam type T_payload_t_i_stream_xbar_sv2v_pfunc_944F6_type
	parameter [31:0] T_IdxWidth = 0;
	parameter [31:0] T_payload_t_DataWidth = 0;
	parameter [31:0] T_payload_t_IdxWidth = 0;
	parameter integer T_payload_t_i_stream_xbar_sv2v_pfunc_944F6 = 0;
	// Trace: design.sv:25496:18
	// removed localparam type T
	// Trace: design.sv:25497:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:25499:3
	input wire clk_i;
	// Trace: design.sv:25500:3
	input wire rst_ni;
	// Trace: design.sv:25501:3
	input wire valid_i;
	// Trace: design.sv:25502:3
	output wire ready_o;
	// Trace: design.sv:25503:3
	input wire [(((T_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + T_payload_t_DataWidth) + T_payload_t_IdxWidth) + T_IdxWidth) - 1:0] data_i;
	// Trace: design.sv:25504:3
	output wire valid_o;
	// Trace: design.sv:25505:3
	input wire ready_i;
	// Trace: design.sv:25506:3
	output wire [(((T_payload_t_i_stream_xbar_sv2v_pfunc_944F6 + T_payload_t_DataWidth) + T_payload_t_IdxWidth) + T_IdxWidth) - 1:0] data_o;
	// Trace: design.sv:25509:3
	spill_register_flushable_AEB2B_E8B2C #(
		.T_T_IdxWidth(T_IdxWidth),
		.T_T_payload_t_DataWidth(T_payload_t_DataWidth),
		.T_T_payload_t_IdxWidth(T_payload_t_IdxWidth),
		.T_T_payload_t_i_stream_xbar_sv2v_pfunc_944F6(T_payload_t_i_stream_xbar_sv2v_pfunc_944F6),
		.Bypass(Bypass)
	) spill_register_flushable_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.valid_i(valid_i),
		.flush_i(1'b0),
		.ready_o(ready_o),
		.data_i(data_i),
		.valid_o(valid_o),
		.ready_i(ready_i),
		.data_o(data_o)
	);
endmodule
module spill_register_1C0C7_8C0C0 (
	clk_i,
	rst_ni,
	valid_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// removed localparam type T_IdxWidth_type
	// removed localparam type T_payload_t_DataWidth_type
	parameter [31:0] T_IdxWidth = 0;
	parameter [31:0] T_payload_t_DataWidth = 0;
	// Trace: design.sv:25496:18
	// removed localparam type T
	// Trace: design.sv:25497:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:25499:3
	input wire clk_i;
	// Trace: design.sv:25500:3
	input wire rst_ni;
	// Trace: design.sv:25501:3
	input wire valid_i;
	// Trace: design.sv:25502:3
	output wire ready_o;
	// Trace: design.sv:25503:3
	input wire [(T_payload_t_DataWidth + T_IdxWidth) - 1:0] data_i;
	// Trace: design.sv:25504:3
	output wire valid_o;
	// Trace: design.sv:25505:3
	input wire ready_i;
	// Trace: design.sv:25506:3
	output wire [(T_payload_t_DataWidth + T_IdxWidth) - 1:0] data_o;
	// Trace: design.sv:25509:3
	spill_register_flushable_918B4_7E477 #(
		.T_T_IdxWidth(T_IdxWidth),
		.T_T_payload_t_DataWidth(T_payload_t_DataWidth),
		.Bypass(Bypass)
	) spill_register_flushable_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.valid_i(valid_i),
		.flush_i(1'b0),
		.ready_o(ready_o),
		.data_i(data_i),
		.valid_o(valid_o),
		.ready_i(ready_i),
		.data_o(data_o)
	);
endmodule
module spill_register_71BB7_B4D1A (
	clk_i,
	rst_ni,
	valid_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// removed localparam type T_T_WIDTH_type
	parameter [31:0] T_T_WIDTH = 0;
	// Trace: design.sv:25496:18
	// removed localparam type T
	// Trace: design.sv:25497:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:25499:3
	input wire clk_i;
	// Trace: design.sv:25500:3
	input wire rst_ni;
	// Trace: design.sv:25501:3
	input wire valid_i;
	// Trace: design.sv:25502:3
	output wire ready_o;
	// Trace: design.sv:25503:3
	input wire [T_T_WIDTH - 1:0] data_i;
	// Trace: design.sv:25504:3
	output wire valid_o;
	// Trace: design.sv:25505:3
	input wire ready_i;
	// Trace: design.sv:25506:3
	output wire [T_T_WIDTH - 1:0] data_o;
	// Trace: design.sv:25509:3
	spill_register_flushable_02CF4_D1AAE #(
		.T_T_T_WIDTH(T_T_WIDTH),
		.Bypass(Bypass)
	) spill_register_flushable_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.valid_i(valid_i),
		.flush_i(1'b0),
		.ready_o(ready_o),
		.data_i(data_i),
		.valid_o(valid_o),
		.ready_i(ready_i),
		.data_o(data_o)
	);
endmodule
module spill_register_736F9 (
	clk_i,
	rst_ni,
	valid_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// Trace: design.sv:25496:18
	// removed localparam type T
	// Trace: design.sv:25497:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:25499:3
	input wire clk_i;
	// Trace: design.sv:25500:3
	input wire rst_ni;
	// Trace: design.sv:25501:3
	input wire valid_i;
	// Trace: design.sv:25502:3
	output wire ready_o;
	// Trace: design.sv:25503:3
	input wire data_i;
	// Trace: design.sv:25504:3
	output wire valid_o;
	// Trace: design.sv:25505:3
	input wire ready_i;
	// Trace: design.sv:25506:3
	output wire data_o;
	// Trace: design.sv:25509:3
	spill_register_flushable_D072E #(.Bypass(Bypass)) spill_register_flushable_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.valid_i(valid_i),
		.flush_i(1'b0),
		.ready_o(ready_o),
		.data_i(data_i),
		.valid_o(valid_o),
		.ready_i(ready_i),
		.data_o(data_o)
	);
endmodule
module spill_register_8294E (
	clk_i,
	rst_ni,
	valid_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// Trace: design.sv:25496:18
	// removed localparam type T
	// Trace: design.sv:25497:13
	parameter [0:0] Bypass = 1'b0;
	// Trace: design.sv:25499:3
	input wire clk_i;
	// Trace: design.sv:25500:3
	input wire rst_ni;
	// Trace: design.sv:25501:3
	input wire valid_i;
	// Trace: design.sv:25502:3
	output wire ready_o;
	// Trace: design.sv:25503:3
	input wire [1:0] data_i;
	// Trace: design.sv:25504:3
	output wire valid_o;
	// Trace: design.sv:25505:3
	input wire ready_i;
	// Trace: design.sv:25506:3
	output wire [1:0] data_o;
	// Trace: design.sv:25509:3
	spill_register_flushable_F9055 #(.Bypass(Bypass)) spill_register_flushable_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.valid_i(valid_i),
		.flush_i(1'b0),
		.ready_o(ready_o),
		.data_i(data_i),
		.valid_o(valid_o),
		.ready_i(ready_i),
		.data_o(data_o)
	);
endmodule
module stream_delay (
	clk_i,
	rst_ni,
	payload_i,
	ready_o,
	valid_i,
	payload_o,
	ready_i,
	valid_o
);
	reg _sv2v_0;
	// Trace: design.sv:25539:15
	parameter [0:0] StallRandom = 0;
	// Trace: design.sv:25540:15
	parameter signed [31:0] FixedDelay = 1;
	// Trace: design.sv:25541:21
	// removed localparam type payload_t
	// Trace: design.sv:25542:15
	parameter [15:0] Seed = 1'sb0;
	// Trace: design.sv:25544:5
	input wire clk_i;
	// Trace: design.sv:25545:5
	input wire rst_ni;
	// Trace: design.sv:25547:5
	input wire payload_i;
	// Trace: design.sv:25548:5
	output reg ready_o;
	// Trace: design.sv:25549:5
	input wire valid_i;
	// Trace: design.sv:25551:5
	output wire payload_o;
	// Trace: design.sv:25552:5
	input wire ready_i;
	// Trace: design.sv:25553:5
	output reg valid_o;
	// Trace: design.sv:25556:5
	generate
		if ((FixedDelay == 0) && !StallRandom) begin : gen_pass_through
			// Trace: design.sv:25557:9
			wire [1:1] sv2v_tmp_0F16F;
			assign sv2v_tmp_0F16F = ready_i;
			always @(*) ready_o = sv2v_tmp_0F16F;
			// Trace: design.sv:25558:9
			wire [1:1] sv2v_tmp_15E2F;
			assign sv2v_tmp_15E2F = valid_i;
			always @(*) valid_o = sv2v_tmp_15E2F;
			// Trace: design.sv:25559:9
			assign payload_o = payload_i;
		end
		else begin : gen_delay
			// Trace: design.sv:25562:9
			localparam [31:0] CounterBits = 4;
			// Trace: design.sv:25564:9
			// removed localparam type state_e
			// Trace: design.sv:25568:9
			reg [1:0] state_d;
			reg [1:0] state_q;
			// Trace: design.sv:25570:9
			reg load;
			// Trace: design.sv:25571:9
			wire [3:0] count_out;
			// Trace: design.sv:25572:9
			reg en;
			// Trace: design.sv:25574:9
			wire [3:0] counter_load;
			// Trace: design.sv:25576:9
			assign payload_o = payload_i;
			// Trace: design.sv:25578:9
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:25579:13
				state_d = state_q;
				// Trace: design.sv:25580:13
				valid_o = 1'b0;
				// Trace: design.sv:25581:13
				ready_o = 1'b0;
				// Trace: design.sv:25582:13
				load = 1'b0;
				// Trace: design.sv:25583:13
				en = 1'b0;
				// Trace: design.sv:25585:13
				(* full_case, parallel_case *)
				case (state_q)
					2'd0:
						// Trace: design.sv:25587:21
						if (valid_i) begin
							// Trace: design.sv:25588:25
							load = 1'b1;
							// Trace: design.sv:25589:25
							state_d = 2'd1;
							// Trace: design.sv:25591:25
							if ((FixedDelay == 1) || (StallRandom && (counter_load == 1)))
								// Trace: design.sv:25592:29
								state_d = 2'd2;
							if (StallRandom && (counter_load == 0)) begin
								// Trace: design.sv:25596:29
								valid_o = 1'b1;
								// Trace: design.sv:25597:29
								ready_o = ready_i;
								// Trace: design.sv:25598:29
								if (ready_i)
									// Trace: design.sv:25598:42
									state_d = 2'd0;
								else
									// Trace: design.sv:25599:34
									state_d = 2'd2;
							end
						end
					2'd1: begin
						// Trace: design.sv:25604:21
						en = 1'b1;
						// Trace: design.sv:25605:21
						if (count_out == 0)
							// Trace: design.sv:25606:25
							state_d = 2'd2;
					end
					2'd2: begin
						// Trace: design.sv:25611:21
						valid_o = 1'b1;
						// Trace: design.sv:25612:21
						ready_o = ready_i;
						// Trace: design.sv:25613:21
						if (ready_i)
							// Trace: design.sv:25613:34
							state_d = 2'd0;
					end
					default:
						;
				endcase
			end
			if (StallRandom) begin : gen_random_stall
				// Trace: design.sv:25621:13
				lfsr_16bit #(
					.WIDTH(16),
					.SEED(Seed)
				) i_lfsr_16bit(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.en_i(load),
					.refill_way_oh(),
					.refill_way_bin(counter_load)
				);
			end
			else begin : gen_fixed_delay
				// Trace: design.sv:25632:13
				assign counter_load = FixedDelay;
			end
			// Trace: design.sv:25635:9
			counter #(.WIDTH(CounterBits)) i_counter(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.clear_i(1'b0),
				.en_i(en),
				.load_i(load),
				.down_i(1'b1),
				.d_i(counter_load),
				.q_o(count_out),
				.overflow_o()
			);
			// Trace: design.sv:25649:9
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:25650:13
				if (~rst_ni)
					// Trace: design.sv:25651:17
					state_q <= 2'd0;
				else
					// Trace: design.sv:25653:17
					state_q <= state_d;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module stream_fifo_7F5E8_FC84F (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	usage_o,
	data_i,
	valid_i,
	ready_o,
	data_o,
	valid_o,
	ready_i
);
	// removed localparam type T_DataWidth_type
	// removed localparam type T_NumBanks_type
	parameter [31:0] T_DataWidth = 0;
	parameter [31:0] T_NumBanks = 0;
	// Trace: design.sv:25673:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:25675:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:25677:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:25678:28
	// removed localparam type T
	// Trace: design.sv:25680:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:25682:5
	input wire clk_i;
	// Trace: design.sv:25683:5
	input wire rst_ni;
	// Trace: design.sv:25684:5
	input wire flush_i;
	// Trace: design.sv:25685:5
	input wire testmode_i;
	// Trace: design.sv:25686:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:25688:5
	input wire [(T_DataWidth / T_NumBanks) - 1:0] data_i;
	// Trace: design.sv:25689:5
	input wire valid_i;
	// Trace: design.sv:25690:5
	output wire ready_o;
	// Trace: design.sv:25692:5
	output wire [(T_DataWidth / T_NumBanks) - 1:0] data_o;
	// Trace: design.sv:25693:5
	output wire valid_o;
	// Trace: design.sv:25694:5
	input wire ready_i;
	// Trace: design.sv:25697:5
	wire push;
	wire pop;
	// Trace: design.sv:25698:5
	wire empty;
	wire full;
	// Trace: design.sv:25700:5
	assign push = valid_i & ~full;
	// Trace: design.sv:25701:5
	assign pop = ready_i & ~empty;
	// Trace: design.sv:25702:5
	assign ready_o = ~full;
	// Trace: design.sv:25703:5
	assign valid_o = ~empty;
	// Trace: design.sv:25705:5
	fifo_v3_DAF99_42EF4 #(
		.dtype_T_DataWidth(T_DataWidth),
		.dtype_T_NumBanks(T_NumBanks),
		.FALL_THROUGH(FALL_THROUGH),
		.DATA_WIDTH(DATA_WIDTH),
		.DEPTH(DEPTH)
	) fifo_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.testmode_i(testmode_i),
		.full_o(full),
		.empty_o(empty),
		.usage_o(usage_o),
		.data_i(data_i),
		.push_i(push),
		.data_o(data_o),
		.pop_i(pop)
	);
endmodule
module stream_fifo_10183 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	usage_o,
	data_i,
	valid_i,
	ready_o,
	data_o,
	valid_o,
	ready_i
);
	// Trace: design.sv:25673:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:25675:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:25677:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:25678:28
	// removed localparam type T
	// Trace: design.sv:25680:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:25682:5
	input wire clk_i;
	// Trace: design.sv:25683:5
	input wire rst_ni;
	// Trace: design.sv:25684:5
	input wire flush_i;
	// Trace: design.sv:25685:5
	input wire testmode_i;
	// Trace: design.sv:25686:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:25688:5
	input wire data_i;
	// Trace: design.sv:25689:5
	input wire valid_i;
	// Trace: design.sv:25690:5
	output wire ready_o;
	// Trace: design.sv:25692:5
	output wire data_o;
	// Trace: design.sv:25693:5
	output wire valid_o;
	// Trace: design.sv:25694:5
	input wire ready_i;
	// Trace: design.sv:25697:5
	wire push;
	wire pop;
	// Trace: design.sv:25698:5
	wire empty;
	wire full;
	// Trace: design.sv:25700:5
	assign push = valid_i & ~full;
	// Trace: design.sv:25701:5
	assign pop = ready_i & ~empty;
	// Trace: design.sv:25702:5
	assign ready_o = ~full;
	// Trace: design.sv:25703:5
	assign valid_o = ~empty;
	// Trace: design.sv:25705:5
	fifo_v3_78C92 #(
		.FALL_THROUGH(FALL_THROUGH),
		.DATA_WIDTH(DATA_WIDTH),
		.DEPTH(DEPTH)
	) fifo_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.testmode_i(testmode_i),
		.full_o(full),
		.empty_o(empty),
		.usage_o(usage_o),
		.data_i(data_i),
		.push_i(push),
		.data_o(data_o),
		.pop_i(pop)
	);
endmodule
module stream_fifo_30B4A_70D5B (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	usage_o,
	data_i,
	valid_i,
	ready_o,
	data_o,
	valid_o,
	ready_i
);
	// removed localparam type T_AddrWidth_type
	// removed localparam type T_AtopWidth_type
	// removed localparam type T_DataWidth_type
	// removed localparam type T_NumBanks_type
	parameter [31:0] T_AddrWidth = 0;
	parameter [31:0] T_AtopWidth = 0;
	parameter [31:0] T_DataWidth = 0;
	parameter [31:0] T_NumBanks = 0;
	// Trace: design.sv:25673:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:25675:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:25677:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:25678:28
	// removed localparam type T
	// Trace: design.sv:25680:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:25682:5
	input wire clk_i;
	// Trace: design.sv:25683:5
	input wire rst_ni;
	// Trace: design.sv:25684:5
	input wire flush_i;
	// Trace: design.sv:25685:5
	input wire testmode_i;
	// Trace: design.sv:25686:5
	output wire [ADDR_DEPTH - 1:0] usage_o;
	// Trace: design.sv:25688:5
	input wire [(((T_AddrWidth + (T_DataWidth / T_NumBanks)) + ((T_DataWidth / T_NumBanks) / 8)) + T_AtopWidth) + 0:0] data_i;
	// Trace: design.sv:25689:5
	input wire valid_i;
	// Trace: design.sv:25690:5
	output wire ready_o;
	// Trace: design.sv:25692:5
	output wire [(((T_AddrWidth + (T_DataWidth / T_NumBanks)) + ((T_DataWidth / T_NumBanks) / 8)) + T_AtopWidth) + 0:0] data_o;
	// Trace: design.sv:25693:5
	output wire valid_o;
	// Trace: design.sv:25694:5
	input wire ready_i;
	// Trace: design.sv:25697:5
	wire push;
	wire pop;
	// Trace: design.sv:25698:5
	wire empty;
	wire full;
	// Trace: design.sv:25700:5
	assign push = valid_i & ~full;
	// Trace: design.sv:25701:5
	assign pop = ready_i & ~empty;
	// Trace: design.sv:25702:5
	assign ready_o = ~full;
	// Trace: design.sv:25703:5
	assign valid_o = ~empty;
	// Trace: design.sv:25705:5
	fifo_v3_463D7_52D08 #(
		.dtype_T_AddrWidth(T_AddrWidth),
		.dtype_T_AtopWidth(T_AtopWidth),
		.dtype_T_DataWidth(T_DataWidth),
		.dtype_T_NumBanks(T_NumBanks),
		.FALL_THROUGH(FALL_THROUGH),
		.DATA_WIDTH(DATA_WIDTH),
		.DEPTH(DEPTH)
	) fifo_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.testmode_i(testmode_i),
		.full_o(full),
		.empty_o(empty),
		.usage_o(usage_o),
		.data_i(data_i),
		.push_i(push),
		.data_o(data_o),
		.pop_i(pop)
	);
endmodule
module stream_fork_dynamic (
	clk_i,
	rst_ni,
	valid_i,
	ready_o,
	sel_i,
	sel_valid_i,
	sel_ready_o,
	valid_o,
	ready_i
);
	reg _sv2v_0;
	// Trace: design.sv:25748:13
	parameter [31:0] N_OUP = 32'd0;
	// Trace: design.sv:25751:3
	input wire clk_i;
	// Trace: design.sv:25753:3
	input wire rst_ni;
	// Trace: design.sv:25755:3
	input wire valid_i;
	// Trace: design.sv:25757:3
	output reg ready_o;
	// Trace: design.sv:25759:3
	input wire [N_OUP - 1:0] sel_i;
	// Trace: design.sv:25761:3
	input wire sel_valid_i;
	// Trace: design.sv:25763:3
	output reg sel_ready_o;
	// Trace: design.sv:25765:3
	output reg [N_OUP - 1:0] valid_o;
	// Trace: design.sv:25767:3
	input wire [N_OUP - 1:0] ready_i;
	// Trace: design.sv:25770:3
	reg int_inp_valid;
	wire int_inp_ready;
	// Trace: design.sv:25771:3
	wire [N_OUP - 1:0] int_oup_valid;
	reg [N_OUP - 1:0] int_oup_ready;
	// Trace: design.sv:25774:3
	genvar _gv_i_16;
	generate
		for (_gv_i_16 = 0; _gv_i_16 < N_OUP; _gv_i_16 = _gv_i_16 + 1) begin : gen_oups
			localparam i = _gv_i_16;
			// Trace: design.sv:25775:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:25776:7
				valid_o[i] = 1'b0;
				// Trace: design.sv:25777:7
				int_oup_ready[i] = 1'b0;
				// Trace: design.sv:25778:7
				if (sel_valid_i) begin
					begin
						// Trace: design.sv:25779:9
						if (sel_i[i]) begin
							// Trace: design.sv:25780:11
							valid_o[i] = int_oup_valid[i];
							// Trace: design.sv:25781:11
							int_oup_ready[i] = ready_i[i];
						end
						else
							// Trace: design.sv:25783:11
							int_oup_ready[i] = 1'b1;
					end
				end
			end
		end
	endgenerate
	// Trace: design.sv:25790:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:25791:5
		int_inp_valid = 1'b0;
		// Trace: design.sv:25792:5
		ready_o = 1'b0;
		// Trace: design.sv:25793:5
		sel_ready_o = 1'b0;
		// Trace: design.sv:25794:5
		if (sel_valid_i) begin
			// Trace: design.sv:25795:7
			int_inp_valid = valid_i;
			// Trace: design.sv:25796:7
			ready_o = int_inp_ready;
			// Trace: design.sv:25797:7
			sel_ready_o = int_inp_ready;
		end
	end
	// Trace: design.sv:25801:3
	stream_fork #(.N_OUP(N_OUP)) i_fork(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.valid_i(int_inp_valid),
		.ready_o(int_inp_ready),
		.valid_o(int_oup_valid),
		.ready_i(int_oup_ready)
	);
	initial _sv2v_0 = 0;
endmodule
module clk_mux_glitch_free (
	clks_i,
	test_clk_i,
	test_en_i,
	async_rstn_i,
	async_sel_i,
	clk_o
);
	reg _sv2v_0;
	// Trace: design.sv:25868:13
	parameter [31:0] NUM_INPUTS = 2;
	// Trace: design.sv:25869:13
	parameter [31:0] NUM_SYNC_STAGES = 2;
	// Trace: design.sv:25870:14
	localparam [31:0] SelWidth = $clog2(NUM_INPUTS);
	// Trace: design.sv:25872:4
	input wire [NUM_INPUTS - 1:0] clks_i;
	// Trace: design.sv:25873:4
	input wire test_clk_i;
	// Trace: design.sv:25874:4
	input wire test_en_i;
	// Trace: design.sv:25875:4
	input wire async_rstn_i;
	// Trace: design.sv:25876:4
	input wire [SelWidth - 1:0] async_sel_i;
	// Trace: design.sv:25877:4
	output wire clk_o;
	// Trace: design.sv:25882:3
	generate
		if (NUM_INPUTS < 2) begin : genblk1
			// Trace: design.sv:25883:5
			$error("Num inputs must be parametrized to a value >= 2.");
		end
	endgenerate
	// Trace: design.sv:25911:3
	reg [NUM_INPUTS - 1:0] s_sel_onehot;
	// Trace: design.sv:25914:3
	reg [(NUM_INPUTS * 2) - 1:0] glitch_filter_d;
	reg [(NUM_INPUTS * 2) - 1:0] glitch_filter_q;
	// Trace: design.sv:25915:3
	wire [NUM_INPUTS - 1:0] s_glitch_filter_output;
	// Trace: design.sv:25916:3
	wire [NUM_INPUTS - 1:0] s_gate_enable;
	// Trace: design.sv:25917:3
	reg [NUM_INPUTS - 1:0] clock_has_been_disabled_q;
	// Trace: design.sv:25918:3
	wire [NUM_INPUTS - 1:0] s_gated_clock;
	// Trace: design.sv:25919:3
	wire s_output_clock;
	// Trace: design.sv:25923:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:25924:5
		s_sel_onehot = 1'sb0;
		// Trace: design.sv:25925:5
		s_sel_onehot[async_sel_i] = 1'b1;
	end
	// Trace: design.sv:25929:3
	genvar _gv_i_17;
	generate
		for (_gv_i_17 = 0; _gv_i_17 < NUM_INPUTS; _gv_i_17 = _gv_i_17 + 1) begin : gen_input_stages
			localparam i = _gv_i_17;
			// Trace: design.sv:25931:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:25932:7
				glitch_filter_d[i * 2] = 1'b1;
				// Trace: design.sv:25933:7
				begin : sv2v_autoblock_1
					// Trace: design.sv:25933:12
					reg signed [31:0] j;
					// Trace: design.sv:25933:12
					for (j = 0; j < NUM_INPUTS; j = j + 1)
						begin
							// Trace: design.sv:25934:9
							if (i == j)
								// Trace: design.sv:25935:11
								glitch_filter_d[i * 2] = glitch_filter_d[i * 2] & s_sel_onehot[j];
							else
								// Trace: design.sv:25937:11
								glitch_filter_d[i * 2] = glitch_filter_d[i * 2] & clock_has_been_disabled_q[j];
						end
				end
			end
			// Trace: design.sv:25941:5
			wire [1:1] sv2v_tmp_B1E63;
			assign sv2v_tmp_B1E63 = glitch_filter_q[i * 2];
			always @(*) glitch_filter_d[(i * 2) + 1] = sv2v_tmp_B1E63;
			// Trace: design.sv:25944:5
			always @(posedge clks_i[i] or negedge async_rstn_i)
				// Trace: design.sv:25945:7
				if (!async_rstn_i)
					// Trace: design.sv:25946:9
					glitch_filter_q[i * 2+:2] <= 1'sb0;
				else
					// Trace: design.sv:25948:9
					glitch_filter_q[i * 2+:2] <= glitch_filter_d[i * 2+:2];
			// Trace: design.sv:25951:5
			assign s_glitch_filter_output[i] = (glitch_filter_q[(i * 2) + 1] & glitch_filter_q[i * 2]) & glitch_filter_d[i * 2];
			// Trace: design.sv:25956:5
			sync #(.STAGES(NUM_SYNC_STAGES)) i_sync_en(
				.clk_i(clks_i[i]),
				.rst_ni(async_rstn_i),
				.serial_i(s_glitch_filter_output[i]),
				.serial_o(s_gate_enable[i])
			);
			// Trace: design.sv:25964:5
			tc_clk_gating #(.IS_FUNCTIONAL(1'b1)) i_clk_gate(
				.clk_i(clks_i[i]),
				.en_i(s_gate_enable[i]),
				.test_en_i(1'b0),
				.clk_o(s_gated_clock[i])
			);
			// Trace: design.sv:25983:5
			always @(posedge clks_i[i] or negedge async_rstn_i)
				// Trace: design.sv:25984:7
				if (!async_rstn_i)
					// Trace: design.sv:25985:9
					clock_has_been_disabled_q[i] <= 1'b0;
				else
					// Trace: design.sv:25987:9
					clock_has_been_disabled_q[i] <= ~s_gate_enable[i];
		end
	endgenerate
	// Trace: design.sv:25996:3
	clk_or_tree #(.NUM_INPUTS(NUM_INPUTS)) i_clk_or_tree(
		.clks_i(s_gated_clock),
		.clk_o(s_output_clock)
	);
	// Trace: design.sv:26002:3
	tc_clk_mux2 i_test_clk_mux(
		.clk0_i(s_output_clock),
		.clk1_i(test_clk_i),
		.clk_sel_i(test_en_i),
		.clk_o(clk_o)
	);
	initial _sv2v_0 = 0;
endmodule
module clk_or_tree (
	clks_i,
	clk_o
);
	// Trace: design.sv:26013:13
	parameter [31:0] NUM_INPUTS = 0;
	// Trace: design.sv:26015:3
	input wire [NUM_INPUTS - 1:0] clks_i;
	// Trace: design.sv:26016:3
	output wire clk_o;
	// Trace: design.sv:26019:3
	generate
		if (NUM_INPUTS < 1) begin : gen_error
			// Trace: design.sv:26020:5
			$error("Cannot parametrize clk_or with less then 1 input but was %0d", NUM_INPUTS);
		end
		else if (NUM_INPUTS == 1) begin : gen_leaf
			// Trace: design.sv:26022:5
			assign clk_o = clks_i[0];
		end
		else if (NUM_INPUTS == 2) begin : gen_leaf
			// Trace: design.sv:26024:5
			tc_clk_or2 i_clk_or2(
				.clk0_i(clks_i[0]),
				.clk1_i(clks_i[1]),
				.clk_o(clk_o)
			);
		end
		else begin : gen_recursive
			// Trace: design.sv:26030:5
			wire branch_a;
			wire branch_b;
			// Trace: design.sv:26031:5
			clk_or_tree #(.NUM_INPUTS(NUM_INPUTS / 2)) i_or_branch_a(
				.clks_i(clks_i[0+:NUM_INPUTS / 2]),
				.clk_o(branch_a)
			);
			// Trace: design.sv:26036:5
			clk_or_tree #(.NUM_INPUTS((NUM_INPUTS / 2) + (NUM_INPUTS % 2))) i_or_branch_b(
				.clks_i(clks_i[NUM_INPUTS - 1:NUM_INPUTS / 2]),
				.clk_o(branch_b)
			);
			// Trace: design.sv:26041:5
			tc_clk_or2 i_clk_or2(
				.clk0_i(branch_a),
				.clk1_i(branch_b),
				.clk_o(clk_o)
			);
		end
	endgenerate
endmodule
module cdc_reset_ctrlr (
	a_clk_i,
	a_rst_ni,
	a_clear_i,
	a_clear_o,
	a_clear_ack_i,
	a_isolate_o,
	a_isolate_ack_i,
	b_clk_i,
	b_rst_ni,
	b_clear_i,
	b_clear_o,
	b_clear_ack_i,
	b_isolate_o,
	b_isolate_ack_i
);
	// removed import cdc_reset_ctrlr_pkg::*;
	// Trace: design.sv:26163:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:26166:13
	parameter [0:0] CLEAR_ON_ASYNC_RESET = 1'b1;
	// Trace: design.sv:26169:3
	input wire a_clk_i;
	// Trace: design.sv:26170:3
	input wire a_rst_ni;
	// Trace: design.sv:26171:3
	input wire a_clear_i;
	// Trace: design.sv:26172:3
	output wire a_clear_o;
	// Trace: design.sv:26173:3
	input wire a_clear_ack_i;
	// Trace: design.sv:26174:3
	output wire a_isolate_o;
	// Trace: design.sv:26175:3
	input wire a_isolate_ack_i;
	// Trace: design.sv:26177:3
	input wire b_clk_i;
	// Trace: design.sv:26178:3
	input wire b_rst_ni;
	// Trace: design.sv:26179:3
	input wire b_clear_i;
	// Trace: design.sv:26180:3
	output wire b_clear_o;
	// Trace: design.sv:26181:3
	input wire b_clear_ack_i;
	// Trace: design.sv:26182:3
	output wire b_isolate_o;
	// Trace: design.sv:26183:3
	input wire b_isolate_ack_i;
	// Trace: design.sv:26187:3
	wire async_a2b_req;
	wire async_b2a_ack;
	// Trace: design.sv:26189:3
	// removed localparam type cdc_reset_ctrlr_pkg_clear_seq_phase_e
	wire [1:0] async_a2b_next_phase;
	// Trace: design.sv:26191:3
	wire async_b2a_req;
	wire async_a2b_ack;
	// Trace: design.sv:26193:3
	wire [1:0] async_b2a_next_phase;
	// Trace: design.sv:26195:3
	cdc_reset_ctrlr_half #(
		.SYNC_STAGES(SYNC_STAGES),
		.CLEAR_ON_ASYNC_RESET(CLEAR_ON_ASYNC_RESET)
	) i_cdc_reset_ctrlr_half_a(
		.clk_i(a_clk_i),
		.rst_ni(a_rst_ni),
		.clear_i(a_clear_i),
		.clear_o(a_clear_o),
		.clear_ack_i(a_clear_ack_i),
		.isolate_o(a_isolate_o),
		.isolate_ack_i(a_isolate_ack_i),
		.async_next_phase_o(async_a2b_next_phase),
		.async_req_o(async_a2b_req),
		.async_ack_i(async_b2a_ack),
		.async_next_phase_i(async_b2a_next_phase),
		.async_req_i(async_b2a_req),
		.async_ack_o(async_a2b_ack)
	);
	// Trace: design.sv:26214:5
	cdc_reset_ctrlr_half #(
		.SYNC_STAGES(SYNC_STAGES),
		.CLEAR_ON_ASYNC_RESET(CLEAR_ON_ASYNC_RESET)
	) i_cdc_reset_ctrlr_half_b(
		.clk_i(b_clk_i),
		.rst_ni(b_rst_ni),
		.clear_i(b_clear_i),
		.clear_o(b_clear_o),
		.clear_ack_i(b_clear_ack_i),
		.isolate_o(b_isolate_o),
		.isolate_ack_i(b_isolate_ack_i),
		.async_next_phase_o(async_b2a_next_phase),
		.async_req_o(async_b2a_req),
		.async_ack_i(async_a2b_ack),
		.async_next_phase_i(async_a2b_next_phase),
		.async_req_i(async_a2b_req),
		.async_ack_o(async_b2a_ack)
	);
endmodule
module cdc_reset_ctrlr_half (
	clk_i,
	rst_ni,
	clear_i,
	isolate_o,
	isolate_ack_i,
	clear_o,
	clear_ack_i,
	async_next_phase_o,
	async_req_o,
	async_ack_i,
	async_next_phase_i,
	async_req_i,
	async_ack_o
);
	reg _sv2v_0;
	// removed import cdc_reset_ctrlr_pkg::*;
	// Trace: design.sv:26241:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:26244:13
	parameter [0:0] CLEAR_ON_ASYNC_RESET = 1'b1;
	// Trace: design.sv:26247:3
	input wire clk_i;
	// Trace: design.sv:26248:3
	input wire rst_ni;
	// Trace: design.sv:26249:3
	input wire clear_i;
	// Trace: design.sv:26250:3
	output wire isolate_o;
	// Trace: design.sv:26251:3
	input wire isolate_ack_i;
	// Trace: design.sv:26252:3
	output wire clear_o;
	// Trace: design.sv:26253:3
	input wire clear_ack_i;
	// Trace: design.sv:26255:3
	// removed localparam type cdc_reset_ctrlr_pkg_clear_seq_phase_e
	output wire [1:0] async_next_phase_o;
	// Trace: design.sv:26256:3
	output wire async_req_o;
	// Trace: design.sv:26257:3
	input wire async_ack_i;
	// Trace: design.sv:26258:3
	input wire [1:0] async_next_phase_i;
	// Trace: design.sv:26259:3
	input wire async_req_i;
	// Trace: design.sv:26260:3
	output wire async_ack_o;
	// Trace: design.sv:26292:4
	// removed localparam type initiator_state_e
	// Trace: design.sv:26303:3
	reg [3:0] initiator_state_d;
	reg [3:0] initiator_state_q;
	// Trace: design.sv:26307:3
	reg [1:0] initiator_clear_seq_phase;
	// Trace: design.sv:26308:3
	reg initiator_phase_transition_req;
	// Trace: design.sv:26309:3
	wire initiator_phase_transition_ack;
	// Trace: design.sv:26310:3
	reg initiator_isolate_out;
	// Trace: design.sv:26311:3
	reg initiator_clear_out;
	// Trace: design.sv:26313:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:26314:5
		initiator_state_d = initiator_state_q;
		// Trace: design.sv:26315:5
		initiator_phase_transition_req = 1'b0;
		// Trace: design.sv:26316:5
		initiator_isolate_out = 1'b0;
		// Trace: design.sv:26317:5
		initiator_clear_out = 1'b0;
		// Trace: design.sv:26318:5
		initiator_clear_seq_phase = 2'd0;
		// Trace: design.sv:26320:5
		case (initiator_state_q)
			4'd0:
				// Trace: design.sv:26322:9
				if (clear_i)
					// Trace: design.sv:26323:11
					initiator_state_d = 4'd1;
			4'd1: begin
				// Trace: design.sv:26328:9
				initiator_phase_transition_req = 1'b1;
				// Trace: design.sv:26329:9
				initiator_clear_seq_phase = 2'd1;
				// Trace: design.sv:26330:9
				initiator_isolate_out = 1'b1;
				// Trace: design.sv:26331:9
				initiator_clear_out = 1'b0;
				// Trace: design.sv:26332:9
				if (initiator_phase_transition_ack && isolate_ack_i)
					// Trace: design.sv:26333:11
					initiator_state_d = 4'd4;
				else if (initiator_phase_transition_ack)
					// Trace: design.sv:26335:11
					initiator_state_d = 4'd3;
				else if (isolate_ack_i)
					// Trace: design.sv:26337:11
					initiator_state_d = 4'd2;
			end
			4'd3: begin
				// Trace: design.sv:26342:9
				initiator_isolate_out = 1'b1;
				// Trace: design.sv:26343:9
				initiator_clear_out = 1'b0;
				// Trace: design.sv:26344:9
				initiator_clear_seq_phase = 2'd1;
				// Trace: design.sv:26345:9
				if (isolate_ack_i)
					// Trace: design.sv:26346:11
					initiator_state_d = 4'd4;
			end
			4'd2: begin
				// Trace: design.sv:26351:9
				initiator_phase_transition_req = 1'b1;
				// Trace: design.sv:26352:9
				initiator_clear_seq_phase = 2'd1;
				// Trace: design.sv:26353:9
				initiator_isolate_out = 1'b1;
				// Trace: design.sv:26354:9
				initiator_clear_out = 1'b0;
				// Trace: design.sv:26355:9
				if (initiator_phase_transition_ack)
					// Trace: design.sv:26356:11
					initiator_state_d = 4'd4;
			end
			4'd4: begin
				// Trace: design.sv:26361:9
				initiator_isolate_out = 1'b1;
				// Trace: design.sv:26362:9
				initiator_clear_out = 1'b1;
				// Trace: design.sv:26363:9
				initiator_phase_transition_req = 1'b1;
				// Trace: design.sv:26364:9
				initiator_clear_seq_phase = 2'd2;
				// Trace: design.sv:26365:9
				if (initiator_phase_transition_ack && clear_ack_i)
					// Trace: design.sv:26366:11
					initiator_state_d = 4'd7;
				else if (initiator_phase_transition_ack)
					// Trace: design.sv:26368:11
					initiator_state_d = 4'd6;
				else if (clear_ack_i)
					// Trace: design.sv:26370:11
					initiator_state_d = 4'd5;
			end
			4'd6: begin
				// Trace: design.sv:26375:9
				initiator_isolate_out = 1'b1;
				// Trace: design.sv:26376:9
				initiator_clear_out = 1'b1;
				// Trace: design.sv:26377:9
				initiator_clear_seq_phase = 2'd2;
				// Trace: design.sv:26378:9
				if (clear_ack_i)
					// Trace: design.sv:26379:11
					initiator_state_d = 4'd7;
			end
			4'd5: begin
				// Trace: design.sv:26384:9
				initiator_phase_transition_req = 1'b1;
				// Trace: design.sv:26385:9
				initiator_clear_seq_phase = 2'd2;
				// Trace: design.sv:26386:9
				initiator_isolate_out = 1'b1;
				// Trace: design.sv:26387:9
				initiator_clear_out = 1'b1;
				// Trace: design.sv:26388:9
				if (initiator_phase_transition_ack)
					// Trace: design.sv:26389:11
					initiator_state_d = 4'd7;
			end
			4'd7: begin
				// Trace: design.sv:26394:9
				initiator_isolate_out = 1'b1;
				// Trace: design.sv:26395:9
				initiator_clear_out = 1'b0;
				// Trace: design.sv:26396:9
				initiator_phase_transition_req = 1'b1;
				// Trace: design.sv:26397:9
				initiator_clear_seq_phase = 2'd3;
				// Trace: design.sv:26398:9
				if (initiator_phase_transition_ack)
					// Trace: design.sv:26399:11
					initiator_state_d = 4'd8;
			end
			4'd8: begin
				// Trace: design.sv:26404:9
				initiator_isolate_out = 1'b1;
				// Trace: design.sv:26405:9
				initiator_clear_out = 1'b0;
				// Trace: design.sv:26406:9
				initiator_phase_transition_req = 1'b1;
				// Trace: design.sv:26407:9
				initiator_clear_seq_phase = 2'd0;
				// Trace: design.sv:26408:9
				if (initiator_phase_transition_ack)
					// Trace: design.sv:26409:11
					initiator_state_d = 4'd0;
			end
			default:
				// Trace: design.sv:26414:9
				initiator_state_d = 4'd1;
		endcase
	end
	// Trace: design.sv:26419:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:26420:5
		if (!rst_ni) begin
			begin
				// Trace: design.sv:26421:7
				if (CLEAR_ON_ASYNC_RESET)
					// Trace: design.sv:26422:9
					initiator_state_q <= 4'd1;
				else
					// Trace: design.sv:26425:9
					initiator_state_q <= 4'd0;
			end
		end
		else
			// Trace: design.sv:26428:7
			initiator_state_q <= initiator_state_d;
	// Trace: design.sv:26437:3
	cdc_4phase_src_DFE1F #(
		.SYNC_STAGES(2),
		.DECOUPLED(0),
		.SEND_RESET_MSG(CLEAR_ON_ASYNC_RESET),
		.RESET_MSG(2'd1)
	) i_state_transition_cdc_src(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.data_i(initiator_clear_seq_phase),
		.valid_i(initiator_phase_transition_req),
		.ready_o(initiator_phase_transition_ack),
		.async_req_o(async_req_o),
		.async_ack_i(async_ack_i),
		.async_data_o(async_next_phase_o)
	);
	// Trace: design.sv:26462:3
	reg [1:0] receiver_phase_q;
	// Trace: design.sv:26463:3
	wire [1:0] receiver_next_phase;
	// Trace: design.sv:26464:3
	wire receiver_phase_req;
	reg receiver_phase_ack;
	// Trace: design.sv:26466:3
	reg receiver_isolate_out;
	// Trace: design.sv:26467:3
	reg receiver_clear_out;
	// Trace: design.sv:26469:3
	cdc_4phase_dst_A46CE #(
		.SYNC_STAGES(2),
		.DECOUPLED(0)
	) i_state_transition_cdc_dst(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.data_o(receiver_next_phase),
		.valid_o(receiver_phase_req),
		.ready_i(receiver_phase_ack),
		.async_req_i(async_req_i),
		.async_ack_o(async_ack_o),
		.async_data_i(async_next_phase_i)
	);
	// Trace: design.sv:26486:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:26487:5
		if (!rst_ni)
			// Trace: design.sv:26488:7
			receiver_phase_q <= 2'd0;
		else if (receiver_phase_req && receiver_phase_ack)
			// Trace: design.sv:26490:7
			receiver_phase_q <= receiver_next_phase;
	// Trace: design.sv:26494:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:26495:5
		receiver_isolate_out = 1'b0;
		// Trace: design.sv:26496:5
		receiver_clear_out = 1'b0;
		// Trace: design.sv:26497:5
		receiver_phase_ack = 1'b0;
		// Trace: design.sv:26500:5
		if (receiver_phase_req)
			// Trace: design.sv:26501:7
			case (receiver_next_phase)
				2'd0: begin
					// Trace: design.sv:26503:11
					receiver_clear_out = 1'b0;
					// Trace: design.sv:26504:11
					receiver_isolate_out = 1'b0;
					// Trace: design.sv:26505:11
					receiver_phase_ack = 1'b1;
				end
				2'd1: begin
					// Trace: design.sv:26509:11
					receiver_clear_out = 1'b0;
					// Trace: design.sv:26510:11
					receiver_isolate_out = 1'b1;
					// Trace: design.sv:26512:11
					receiver_phase_ack = isolate_ack_i;
				end
				2'd2: begin
					// Trace: design.sv:26516:11
					receiver_clear_out = 1'b1;
					// Trace: design.sv:26517:11
					receiver_isolate_out = 1'b1;
					// Trace: design.sv:26519:11
					receiver_phase_ack = clear_ack_i;
				end
				2'd3: begin
					// Trace: design.sv:26523:11
					receiver_clear_out = 1'b0;
					// Trace: design.sv:26524:11
					receiver_isolate_out = 1'b1;
					// Trace: design.sv:26525:11
					receiver_phase_ack = 1'b1;
				end
				default: begin
					// Trace: design.sv:26529:11
					receiver_clear_out = 1'b0;
					// Trace: design.sv:26530:11
					receiver_isolate_out = 1'b0;
					// Trace: design.sv:26531:11
					receiver_phase_ack = 1'b0;
				end
			endcase
		else
			// Trace: design.sv:26538:7
			case (receiver_phase_q)
				2'd0: begin
					// Trace: design.sv:26540:11
					receiver_clear_out = 1'b0;
					// Trace: design.sv:26541:11
					receiver_isolate_out = 1'b0;
				end
				2'd1: begin
					// Trace: design.sv:26545:11
					receiver_clear_out = 1'b0;
					// Trace: design.sv:26546:11
					receiver_isolate_out = 1'b1;
				end
				2'd2: begin
					// Trace: design.sv:26550:11
					receiver_clear_out = 1'b1;
					// Trace: design.sv:26551:11
					receiver_isolate_out = 1'b1;
				end
				2'd3: begin
					// Trace: design.sv:26555:11
					receiver_clear_out = 1'b0;
					// Trace: design.sv:26556:11
					receiver_isolate_out = 1'b1;
				end
				default: begin
					// Trace: design.sv:26560:11
					receiver_clear_out = 1'b0;
					// Trace: design.sv:26561:11
					receiver_isolate_out = 1'b0;
					// Trace: design.sv:26562:11
					receiver_phase_ack = 1'b0;
				end
			endcase
	end
	// Trace: design.sv:26574:3
	assign clear_o = initiator_clear_out || receiver_clear_out;
	// Trace: design.sv:26575:3
	assign isolate_o = initiator_isolate_out || receiver_isolate_out;
	initial _sv2v_0 = 0;
endmodule
module cdc_fifo_gray (
	src_rst_ni,
	src_clk_i,
	src_data_i,
	src_valid_i,
	src_ready_o,
	dst_rst_ni,
	dst_clk_i,
	dst_data_o,
	dst_valid_o,
	dst_ready_i
);
	// Trace: design.sv:26681:13
	parameter [31:0] WIDTH = 1;
	// Trace: design.sv:26683:18
	// removed localparam type T
	// Trace: design.sv:26685:13
	parameter signed [31:0] LOG_DEPTH = 3;
	// Trace: design.sv:26687:13
	parameter signed [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:26689:3
	input wire src_rst_ni;
	// Trace: design.sv:26690:3
	input wire src_clk_i;
	// Trace: design.sv:26691:3
	input wire [WIDTH - 1:0] src_data_i;
	// Trace: design.sv:26692:3
	input wire src_valid_i;
	// Trace: design.sv:26693:3
	output wire src_ready_o;
	// Trace: design.sv:26695:3
	input wire dst_rst_ni;
	// Trace: design.sv:26696:3
	input wire dst_clk_i;
	// Trace: design.sv:26697:3
	output wire [WIDTH - 1:0] dst_data_o;
	// Trace: design.sv:26698:3
	output wire dst_valid_o;
	// Trace: design.sv:26699:3
	input wire dst_ready_i;
	// Trace: design.sv:26702:3
	wire [((2 ** LOG_DEPTH) * WIDTH) - 1:0] async_data;
	// Trace: design.sv:26703:3
	wire [LOG_DEPTH:0] async_wptr;
	// Trace: design.sv:26704:3
	wire [LOG_DEPTH:0] async_rptr;
	// Trace: design.sv:26706:3
	cdc_fifo_gray_src_82E7A_2EAD4 #(
		.T_WIDTH(WIDTH),
		.LOG_DEPTH(LOG_DEPTH)
	) i_src(
		.src_rst_ni(src_rst_ni),
		.src_clk_i(src_clk_i),
		.src_data_i(src_data_i),
		.src_valid_i(src_valid_i),
		.src_ready_o(src_ready_o),
		.async_data_o(async_data),
		.async_wptr_o(async_wptr),
		.async_rptr_i(async_rptr)
	);
	// Trace: design.sv:26721:3
	cdc_fifo_gray_dst_55D7B_215FD #(
		.T_WIDTH(WIDTH),
		.LOG_DEPTH(LOG_DEPTH)
	) i_dst(
		.dst_rst_ni(dst_rst_ni),
		.dst_clk_i(dst_clk_i),
		.dst_data_o(dst_data_o),
		.dst_valid_o(dst_valid_o),
		.dst_ready_i(dst_ready_i),
		.async_data_i(async_data),
		.async_wptr_i(async_wptr),
		.async_rptr_o(async_rptr)
	);
endmodule
module cdc_fifo_gray_src_82E7A_2EAD4 (
	src_rst_ni,
	src_clk_i,
	src_data_i,
	src_valid_i,
	src_ready_o,
	async_data_o,
	async_wptr_o,
	async_rptr_i
);
	// removed localparam type T_WIDTH_type
	parameter [31:0] T_WIDTH = 0;
	// Trace: design.sv:26750:18
	// removed localparam type T
	// Trace: design.sv:26751:13
	parameter signed [31:0] LOG_DEPTH = 3;
	// Trace: design.sv:26752:13
	parameter signed [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:26754:3
	input wire src_rst_ni;
	// Trace: design.sv:26755:3
	input wire src_clk_i;
	// Trace: design.sv:26756:3
	input wire [T_WIDTH - 1:0] src_data_i;
	// Trace: design.sv:26757:3
	input wire src_valid_i;
	// Trace: design.sv:26758:3
	output wire src_ready_o;
	// Trace: design.sv:26760:3
	output wire [((2 ** LOG_DEPTH) * T_WIDTH) - 1:0] async_data_o;
	// Trace: design.sv:26761:3
	output wire [LOG_DEPTH:0] async_wptr_o;
	// Trace: design.sv:26762:3
	input wire [LOG_DEPTH:0] async_rptr_i;
	// Trace: design.sv:26765:3
	localparam signed [31:0] PtrWidth = LOG_DEPTH + 1;
	// Trace: design.sv:26766:3
	localparam [PtrWidth - 1:0] PtrFull = 1 << LOG_DEPTH;
	// Trace: design.sv:26768:3
	reg [((2 ** LOG_DEPTH) * T_WIDTH) - 1:0] data_q;
	// Trace: design.sv:26769:3
	reg [PtrWidth - 1:0] wptr_q;
	wire [PtrWidth - 1:0] wptr_d;
	wire [PtrWidth - 1:0] wptr_bin;
	wire [PtrWidth - 1:0] wptr_next;
	wire [PtrWidth - 1:0] rptr;
	wire [PtrWidth - 1:0] rptr_bin;
	// Trace: design.sv:26772:3
	assign async_data_o = data_q;
	// Trace: design.sv:26773:3
	genvar _gv_i_18;
	generate
		for (_gv_i_18 = 0; _gv_i_18 < (2 ** LOG_DEPTH); _gv_i_18 = _gv_i_18 + 1) begin : gen_word
			localparam i = _gv_i_18;
			// Trace: macro expansion of FFLNR at design.sv:26775:78
			always @(posedge src_clk_i)
				// Trace: macro expansion of FFLNR at design.sv:26775:120
				if ((src_valid_i & src_ready_o) & (wptr_bin[LOG_DEPTH - 1:0] == i))
					// Trace: macro expansion of FFLNR at design.sv:26775:162
					data_q[i * T_WIDTH+:T_WIDTH] <= src_data_i;
		end
	endgenerate
	// Trace: design.sv:26779:3
	genvar _gv_i_19;
	generate
		for (_gv_i_19 = 0; _gv_i_19 < PtrWidth; _gv_i_19 = _gv_i_19 + 1) begin : gen_sync
			localparam i = _gv_i_19;
			// Trace: design.sv:26780:5
			sync #(.STAGES(SYNC_STAGES)) i_sync(
				.clk_i(src_clk_i),
				.rst_ni(src_rst_ni),
				.serial_i(async_rptr_i[i]),
				.serial_o(rptr[i])
			);
		end
	endgenerate
	// Trace: design.sv:26787:3
	gray_to_binary #(.N(PtrWidth)) i_rptr_g2b(
		.A(rptr),
		.Z(rptr_bin)
	);
	// Trace: design.sv:26790:3
	assign wptr_next = wptr_bin + 1;
	// Trace: design.sv:26791:3
	gray_to_binary #(.N(PtrWidth)) i_wptr_g2b(
		.A(wptr_q),
		.Z(wptr_bin)
	);
	// Trace: design.sv:26792:3
	binary_to_gray #(.N(PtrWidth)) i_wptr_b2g(
		.A(wptr_next),
		.Z(wptr_d)
	);
	// Trace: macro expansion of FFL at design.sv:26793:129
	always @(posedge src_clk_i or negedge src_rst_ni)
		// Trace: macro expansion of FFL at design.sv:26793:226
		if (!src_rst_ni)
			// Trace: macro expansion of FFL at design.sv:26793:323
			wptr_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at design.sv:26793:513
			if (src_valid_i & src_ready_o)
				// Trace: macro expansion of FFL at design.sv:26793:610
				wptr_q <= wptr_d;
	// Trace: design.sv:26794:3
	assign async_wptr_o = wptr_q;
	// Trace: design.sv:26800:3
	assign src_ready_o = (wptr_bin ^ rptr_bin) != PtrFull;
endmodule
module cdc_fifo_gray_dst_55D7B_215FD (
	dst_rst_ni,
	dst_clk_i,
	dst_data_o,
	dst_valid_o,
	dst_ready_i,
	async_data_i,
	async_wptr_i,
	async_rptr_o
);
	// removed localparam type T_WIDTH_type
	parameter [31:0] T_WIDTH = 0;
	// Trace: design.sv:26808:18
	// removed localparam type T
	// Trace: design.sv:26809:13
	parameter signed [31:0] LOG_DEPTH = 3;
	// Trace: design.sv:26810:13
	parameter signed [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:26812:3
	input wire dst_rst_ni;
	// Trace: design.sv:26813:3
	input wire dst_clk_i;
	// Trace: design.sv:26814:3
	output wire [T_WIDTH - 1:0] dst_data_o;
	// Trace: design.sv:26815:3
	output wire dst_valid_o;
	// Trace: design.sv:26816:3
	input wire dst_ready_i;
	// Trace: design.sv:26818:3
	input wire [((2 ** LOG_DEPTH) * T_WIDTH) - 1:0] async_data_i;
	// Trace: design.sv:26819:3
	input wire [LOG_DEPTH:0] async_wptr_i;
	// Trace: design.sv:26820:3
	output wire [LOG_DEPTH:0] async_rptr_o;
	// Trace: design.sv:26823:3
	localparam signed [31:0] PtrWidth = LOG_DEPTH + 1;
	// Trace: design.sv:26824:3
	localparam [PtrWidth - 1:0] PtrEmpty = 1'sb0;
	// Trace: design.sv:26826:3
	wire [T_WIDTH - 1:0] dst_data;
	// Trace: design.sv:26827:3
	reg [PtrWidth - 1:0] rptr_q;
	wire [PtrWidth - 1:0] rptr_d;
	wire [PtrWidth - 1:0] rptr_bin;
	wire [PtrWidth - 1:0] rptr_bin_d;
	wire [PtrWidth - 1:0] rptr_next;
	wire [PtrWidth - 1:0] wptr;
	wire [PtrWidth - 1:0] wptr_bin;
	// Trace: design.sv:26828:3
	wire dst_valid;
	wire dst_ready;
	// Trace: design.sv:26830:3
	assign dst_data = async_data_i[rptr_bin[LOG_DEPTH - 1:0] * T_WIDTH+:T_WIDTH];
	// Trace: design.sv:26833:3
	assign rptr_next = rptr_bin + 1;
	// Trace: design.sv:26834:3
	gray_to_binary #(.N(PtrWidth)) i_rptr_g2b(
		.A(rptr_q),
		.Z(rptr_bin)
	);
	// Trace: design.sv:26835:3
	binary_to_gray #(.N(PtrWidth)) i_rptr_b2g(
		.A(rptr_next),
		.Z(rptr_d)
	);
	// Trace: macro expansion of FFL at design.sv:26836:125
	always @(posedge dst_clk_i or negedge dst_rst_ni)
		// Trace: macro expansion of FFL at design.sv:26836:222
		if (!dst_rst_ni)
			// Trace: macro expansion of FFL at design.sv:26836:319
			rptr_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at design.sv:26836:509
			if (dst_valid & dst_ready)
				// Trace: macro expansion of FFL at design.sv:26836:606
				rptr_q <= rptr_d;
	// Trace: design.sv:26837:3
	assign async_rptr_o = rptr_q;
	// Trace: design.sv:26840:3
	genvar _gv_i_20;
	generate
		for (_gv_i_20 = 0; _gv_i_20 < PtrWidth; _gv_i_20 = _gv_i_20 + 1) begin : gen_sync
			localparam i = _gv_i_20;
			// Trace: design.sv:26841:5
			sync #(.STAGES(SYNC_STAGES)) i_sync(
				.clk_i(dst_clk_i),
				.rst_ni(dst_rst_ni),
				.serial_i(async_wptr_i[i]),
				.serial_o(wptr[i])
			);
		end
	endgenerate
	// Trace: design.sv:26848:3
	gray_to_binary #(.N(PtrWidth)) i_wptr_g2b(
		.A(wptr),
		.Z(wptr_bin)
	);
	// Trace: design.sv:26854:3
	assign dst_valid = (wptr_bin ^ rptr_bin) != PtrEmpty;
	// Trace: design.sv:26857:3
	spill_register_71BB7_B4D1A #(.T_T_WIDTH(T_WIDTH)) i_spill_register(
		.clk_i(dst_clk_i),
		.rst_ni(dst_rst_ni),
		.valid_i(dst_valid),
		.ready_o(dst_ready),
		.data_i(dst_data),
		.valid_o(dst_valid_o),
		.ready_i(dst_ready_i),
		.data_o(dst_data_o)
	);
endmodule
module fall_through_register (
	clk_i,
	rst_ni,
	clr_i,
	testmode_i,
	valid_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// Trace: design.sv:26886:20
	// removed localparam type T
	// Trace: design.sv:26888:5
	input wire clk_i;
	// Trace: design.sv:26889:5
	input wire rst_ni;
	// Trace: design.sv:26890:5
	input wire clr_i;
	// Trace: design.sv:26891:5
	input wire testmode_i;
	// Trace: design.sv:26893:5
	input wire valid_i;
	// Trace: design.sv:26894:5
	output wire ready_o;
	// Trace: design.sv:26895:5
	input wire data_i;
	// Trace: design.sv:26897:5
	output wire valid_o;
	// Trace: design.sv:26898:5
	input wire ready_i;
	// Trace: design.sv:26899:5
	output wire data_o;
	// Trace: design.sv:26902:5
	wire fifo_empty;
	wire fifo_full;
	// Trace: design.sv:26905:5
	fifo_v3_78C92 #(
		.FALL_THROUGH(1'b1),
		.DEPTH(1)
	) i_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(clr_i),
		.testmode_i(testmode_i),
		.full_o(fifo_full),
		.empty_o(fifo_empty),
		.usage_o(),
		.data_i(data_i),
		.push_i(valid_i & ~fifo_full),
		.data_o(data_o),
		.pop_i(ready_i & ~fifo_empty)
	);
	// Trace: design.sv:26923:5
	assign ready_o = ~fifo_full;
	// Trace: design.sv:26924:5
	assign valid_o = ~fifo_empty;
endmodule
module id_queue (
	clk_i,
	rst_ni,
	inp_id_i,
	inp_data_i,
	inp_req_i,
	inp_gnt_o,
	exists_data_i,
	exists_mask_i,
	exists_req_i,
	exists_o,
	exists_gnt_o,
	oup_id_i,
	oup_pop_i,
	oup_req_i,
	oup_data_o,
	oup_data_valid_o,
	oup_gnt_o
);
	reg _sv2v_0;
	// Trace: design.sv:26975:15
	parameter signed [31:0] ID_WIDTH = 0;
	// Trace: design.sv:26976:15
	parameter signed [31:0] CAPACITY = 0;
	// Trace: design.sv:26977:15
	parameter [0:0] FULL_BW = 0;
	// Trace: design.sv:26978:20
	// removed localparam type data_t
	// Trace: design.sv:26980:21
	// removed localparam type id_t
	// Trace: design.sv:26982:5
	input wire clk_i;
	// Trace: design.sv:26983:5
	input wire rst_ni;
	// Trace: design.sv:26985:5
	input wire [ID_WIDTH - 1:0] inp_id_i;
	// Trace: design.sv:26986:5
	input wire [31:0] inp_data_i;
	// Trace: design.sv:26987:5
	input wire inp_req_i;
	// Trace: design.sv:26988:5
	output wire inp_gnt_o;
	// Trace: design.sv:26990:5
	input wire [31:0] exists_data_i;
	// Trace: design.sv:26991:5
	input wire [31:0] exists_mask_i;
	// Trace: design.sv:26992:5
	input wire exists_req_i;
	// Trace: design.sv:26993:5
	output reg exists_o;
	// Trace: design.sv:26994:5
	output reg exists_gnt_o;
	// Trace: design.sv:26996:5
	input wire [ID_WIDTH - 1:0] oup_id_i;
	// Trace: design.sv:26997:5
	input wire oup_pop_i;
	// Trace: design.sv:26998:5
	input wire oup_req_i;
	// Trace: design.sv:26999:5
	output reg [31:0] oup_data_o;
	// Trace: design.sv:27000:5
	output reg oup_data_valid_o;
	// Trace: design.sv:27001:5
	output reg oup_gnt_o;
	// Trace: design.sv:27006:5
	localparam signed [31:0] NIds = 2 ** ID_WIDTH;
	// Trace: design.sv:27007:5
	localparam signed [31:0] HtCapacity = (NIds <= CAPACITY ? NIds : CAPACITY);
	// Trace: design.sv:27008:5
	function automatic [31:0] cf_math_pkg_idx_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:58:9
		cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	localparam [31:0] HtIdxWidth = cf_math_pkg_idx_width(HtCapacity);
	// Trace: design.sv:27009:5
	localparam [31:0] LdIdxWidth = cf_math_pkg_idx_width(CAPACITY);
	// Trace: design.sv:27012:5
	// removed localparam type ht_idx_t
	// Trace: design.sv:27015:5
	// removed localparam type ld_idx_t
	// Trace: design.sv:27018:5
	// removed localparam type head_tail_t
	// Trace: design.sv:27026:5
	// removed localparam type linked_data_t
	// Trace: design.sv:27032:5
	reg [((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (HtCapacity * (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1)) - 1 : (HtCapacity * (1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) - 1)):((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)] head_tail_d;
	reg [((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (HtCapacity * (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1)) - 1 : (HtCapacity * (1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) - 1)):((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)] head_tail_q;
	// Trace: design.sv:27034:5
	reg [(((32 + LdIdxWidth) + 0) >= 0 ? (CAPACITY * ((32 + LdIdxWidth) + 1)) - 1 : (CAPACITY * (1 - ((32 + LdIdxWidth) + 0))) + ((32 + LdIdxWidth) - 1)):(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0)] linked_data_d;
	reg [(((32 + LdIdxWidth) + 0) >= 0 ? (CAPACITY * ((32 + LdIdxWidth) + 1)) - 1 : (CAPACITY * (1 - ((32 + LdIdxWidth) + 0))) + ((32 + LdIdxWidth) - 1)):(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0)] linked_data_q;
	// Trace: design.sv:27036:5
	wire full;
	reg match_in_id_valid;
	reg match_out_id_valid;
	wire no_in_id_match;
	wire no_out_id_match;
	// Trace: design.sv:27042:5
	wire [HtCapacity - 1:0] head_tail_free;
	wire [HtCapacity - 1:0] idx_matches_in_id;
	wire [HtCapacity - 1:0] idx_matches_out_id;
	// Trace: design.sv:27046:5
	wire [CAPACITY - 1:0] exists_match;
	wire [CAPACITY - 1:0] linked_data_free;
	// Trace: design.sv:27049:5
	reg [ID_WIDTH - 1:0] match_in_id;
	reg [ID_WIDTH - 1:0] match_out_id;
	// Trace: design.sv:27051:5
	wire [HtIdxWidth - 1:0] head_tail_free_idx;
	wire [HtIdxWidth - 1:0] match_in_idx;
	wire [HtIdxWidth - 1:0] match_out_idx;
	// Trace: design.sv:27055:5
	wire [LdIdxWidth - 1:0] linked_data_free_idx;
	wire [LdIdxWidth - 1:0] oup_data_free_idx;
	// Trace: design.sv:27058:5
	reg oup_data_popped;
	reg oup_ht_popped;
	// Trace: design.sv:27062:5
	genvar _gv_i_21;
	generate
		for (_gv_i_21 = 0; _gv_i_21 < HtCapacity; _gv_i_21 = _gv_i_21 + 1) begin : gen_idx_match
			localparam i = _gv_i_21;
			// Trace: design.sv:27063:9
			assign idx_matches_in_id[i] = (match_in_id_valid && (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)))) : (((i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))))) + ((ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))) >= (LdIdxWidth + (LdIdxWidth + 1)) ? ((ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))) - (LdIdxWidth + (LdIdxWidth + 1))) + 1 : ((LdIdxWidth + (LdIdxWidth + 1)) - (ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)))) + 1)) - 1)-:((ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))) >= (LdIdxWidth + (LdIdxWidth + 1)) ? ((ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))) - (LdIdxWidth + (LdIdxWidth + 1))) + 1 : ((LdIdxWidth + (LdIdxWidth + 1)) - (ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)))) + 1)] == match_in_id)) && !head_tail_q[(i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)];
			// Trace: design.sv:27065:9
			assign idx_matches_out_id[i] = (match_out_id_valid && (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)))) : (((i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))))) + ((ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))) >= (LdIdxWidth + (LdIdxWidth + 1)) ? ((ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))) - (LdIdxWidth + (LdIdxWidth + 1))) + 1 : ((LdIdxWidth + (LdIdxWidth + 1)) - (ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)))) + 1)) - 1)-:((ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))) >= (LdIdxWidth + (LdIdxWidth + 1)) ? ((ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0))) - (LdIdxWidth + (LdIdxWidth + 1))) + 1 : ((LdIdxWidth + (LdIdxWidth + 1)) - (ID_WIDTH + (LdIdxWidth + (LdIdxWidth + 0)))) + 1)] == match_out_id)) && !head_tail_q[(i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)];
		end
	endgenerate
	// Trace: design.sv:27068:5
	assign no_in_id_match = !(|idx_matches_in_id);
	// Trace: design.sv:27069:5
	assign no_out_id_match = !(|idx_matches_out_id);
	// Trace: design.sv:27070:5
	onehot_to_bin #(.ONEHOT_WIDTH(HtCapacity)) i_id_ohb_in(
		.onehot(idx_matches_in_id),
		.bin(match_in_idx)
	);
	// Trace: design.sv:27076:5
	onehot_to_bin #(.ONEHOT_WIDTH(HtCapacity)) i_id_ohb_out(
		.onehot(idx_matches_out_id),
		.bin(match_out_idx)
	);
	// Trace: design.sv:27084:5
	genvar _gv_i_22;
	generate
		for (_gv_i_22 = 0; _gv_i_22 < HtCapacity; _gv_i_22 = _gv_i_22 + 1) begin : gen_head_tail_free
			localparam i = _gv_i_22;
			// Trace: design.sv:27085:9
			assign head_tail_free[i] = head_tail_q[(i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)];
		end
	endgenerate
	// Trace: design.sv:27087:5
	lzc #(
		.WIDTH(HtCapacity),
		.MODE(0)
	) i_ht_free_lzc(
		.in_i(head_tail_free),
		.cnt_o(head_tail_free_idx),
		.empty_o()
	);
	// Trace: design.sv:27097:5
	genvar _gv_i_23;
	generate
		for (_gv_i_23 = 0; _gv_i_23 < CAPACITY; _gv_i_23 = _gv_i_23 + 1) begin : gen_linked_data_free
			localparam i = _gv_i_23;
			// Trace: design.sv:27098:9
			assign linked_data_free[i] = linked_data_q[(i * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0)];
		end
	endgenerate
	// Trace: design.sv:27100:5
	lzc #(
		.WIDTH(CAPACITY),
		.MODE(0)
	) i_ld_free_lzc(
		.in_i(linked_data_free),
		.cnt_o(linked_data_free_idx),
		.empty_o()
	);
	// Trace: design.sv:27110:5
	assign full = !(|linked_data_free);
	// Trace: design.sv:27112:5
	assign oup_data_free_idx = head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)];
	// Trace: design.sv:27115:5
	assign inp_gnt_o = ~full || (oup_data_popped && FULL_BW);
	// Trace: design.sv:27116:5
	function automatic [ID_WIDTH - 1:0] sv2v_cast_64419;
		input reg [ID_WIDTH - 1:0] inp;
		sv2v_cast_64419 = inp;
	endfunction
	function automatic [LdIdxWidth - 1:0] sv2v_cast_1B5F4;
		input reg [LdIdxWidth - 1:0] inp;
		sv2v_cast_1B5F4 = inp;
	endfunction
	function automatic [ID_WIDTH - 1:0] sv2v_cast_37B7D;
		input reg [ID_WIDTH - 1:0] inp;
		sv2v_cast_37B7D = inp;
	endfunction
	function automatic [LdIdxWidth - 1:0] sv2v_cast_D5FF0;
		input reg [LdIdxWidth - 1:0] inp;
		sv2v_cast_D5FF0 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:27117:9
		match_in_id = 1'sb0;
		// Trace: design.sv:27118:9
		match_out_id = 1'sb0;
		// Trace: design.sv:27119:9
		match_in_id_valid = 1'b0;
		// Trace: design.sv:27120:9
		match_out_id_valid = 1'b0;
		// Trace: design.sv:27121:9
		head_tail_d = head_tail_q;
		// Trace: design.sv:27122:9
		linked_data_d = linked_data_q;
		// Trace: design.sv:27123:9
		oup_gnt_o = 1'b0;
		// Trace: design.sv:27124:9
		oup_data_o = 32'b00000000000000000000000000000000;
		// Trace: design.sv:27125:9
		oup_data_valid_o = 1'b0;
		// Trace: design.sv:27126:9
		oup_data_popped = 1'b0;
		// Trace: design.sv:27127:9
		oup_ht_popped = 1'b0;
		// Trace: design.sv:27129:9
		if (!FULL_BW) begin
			begin
				// Trace: design.sv:27130:13
				if (inp_req_i && !full) begin
					// Trace: design.sv:27131:17
					match_in_id = inp_id_i;
					// Trace: design.sv:27132:17
					match_in_id_valid = 1'b1;
					// Trace: design.sv:27134:17
					if (no_in_id_match)
						// Trace: design.sv:27135:21
						head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (head_tail_free_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] = {sv2v_cast_64419(inp_id_i), sv2v_cast_1B5F4(linked_data_free_idx), sv2v_cast_1B5F4(linked_data_free_idx), 1'b0};
					else begin
						// Trace: design.sv:27143:21
						linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] = linked_data_free_idx;
						// Trace: design.sv:27144:21
						head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] = linked_data_free_idx;
					end
					// Trace: design.sv:27146:17
					linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (linked_data_free_idx * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = {inp_data_i, sv2v_cast_1B5F4(1'sb0), 1'b0};
				end
				else if (oup_req_i) begin
					// Trace: design.sv:27152:17
					match_in_id = oup_id_i;
					// Trace: design.sv:27153:17
					match_in_id_valid = 1'b1;
					// Trace: design.sv:27154:17
					if (!no_in_id_match) begin
						// Trace: design.sv:27155:21
						oup_data_o = sv2v_cast_32(linked_data_q[(((32 + LdIdxWidth) + 0) >= 0 ? (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 32 + (LdIdxWidth + 0) : ((32 + LdIdxWidth) + 0) - (32 + (LdIdxWidth + 0))) : (((head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 32 + (LdIdxWidth + 0) : ((32 + LdIdxWidth) + 0) - (32 + (LdIdxWidth + 0)))) + ((32 + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((32 + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (32 + (LdIdxWidth + 0))) + 1)) - 1)-:((32 + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((32 + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (32 + (LdIdxWidth + 0))) + 1)]);
						// Trace: design.sv:27156:21
						oup_data_valid_o = 1'b1;
						// Trace: design.sv:27157:21
						if (oup_pop_i) begin
							// Trace: design.sv:27159:25
							linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = 1'sb0;
							// Trace: design.sv:27160:25
							linked_data_d[(head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0)] = 1'b1;
							// Trace: design.sv:27161:25
							if (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] == head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))])
								// Trace: design.sv:27162:29
								head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] = {sv2v_cast_37B7D(1'sb0), sv2v_cast_D5FF0(1'sb0), sv2v_cast_D5FF0(1'sb0), 1'b1};
							else
								// Trace: design.sv:27164:29
								head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] = linked_data_q[(((32 + LdIdxWidth) + 0) >= 0 ? (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))];
						end
					end
					// Trace: design.sv:27171:17
					oup_gnt_o = 1'b1;
				end
			end
		end
		else begin
			// Trace: design.sv:27175:13
			if (oup_req_i) begin
				// Trace: design.sv:27176:17
				match_out_id = oup_id_i;
				// Trace: design.sv:27177:17
				match_out_id_valid = 1'b1;
				// Trace: design.sv:27178:17
				if (!no_out_id_match) begin
					// Trace: design.sv:27179:21
					oup_data_o = sv2v_cast_32(linked_data_q[(((32 + LdIdxWidth) + 0) >= 0 ? (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 32 + (LdIdxWidth + 0) : ((32 + LdIdxWidth) + 0) - (32 + (LdIdxWidth + 0))) : (((head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 32 + (LdIdxWidth + 0) : ((32 + LdIdxWidth) + 0) - (32 + (LdIdxWidth + 0)))) + ((32 + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((32 + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (32 + (LdIdxWidth + 0))) + 1)) - 1)-:((32 + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((32 + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (32 + (LdIdxWidth + 0))) + 1)]);
					// Trace: design.sv:27180:21
					oup_data_valid_o = 1'b1;
					// Trace: design.sv:27181:21
					if (oup_pop_i) begin
						// Trace: design.sv:27182:25
						oup_data_popped = 1'b1;
						// Trace: design.sv:27184:25
						linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = 1'sb0;
						// Trace: design.sv:27185:25
						linked_data_d[(head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0)] = 1'b1;
						// Trace: design.sv:27186:25
						if (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] == head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))]) begin
							// Trace: design.sv:27188:29
							oup_ht_popped = 1'b1;
							// Trace: design.sv:27189:29
							head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] = {sv2v_cast_37B7D(1'sb0), sv2v_cast_D5FF0(1'sb0), sv2v_cast_D5FF0(1'sb0), 1'b1};
						end
						else
							// Trace: design.sv:27191:29
							head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] = linked_data_q[(((32 + LdIdxWidth) + 0) >= 0 ? (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0))) : (((match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + (LdIdxWidth + 0) : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + (LdIdxWidth + 0)))) + ((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)) - 1)-:((LdIdxWidth + (LdIdxWidth + 0)) >= (LdIdxWidth + 1) ? ((LdIdxWidth + (LdIdxWidth + 0)) - (LdIdxWidth + 1)) + 1 : ((LdIdxWidth + 1) - (LdIdxWidth + (LdIdxWidth + 0))) + 1)] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))];
					end
				end
				// Trace: design.sv:27198:17
				oup_gnt_o = 1'b1;
			end
			if (inp_req_i && inp_gnt_o) begin
				// Trace: design.sv:27201:17
				match_in_id = inp_id_i;
				// Trace: design.sv:27202:17
				match_in_id_valid = 1'b1;
				// Trace: design.sv:27204:17
				if (oup_ht_popped && (oup_id_i == inp_id_i)) begin
					// Trace: design.sv:27207:21
					head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] = {sv2v_cast_64419(inp_id_i), sv2v_cast_1B5F4(oup_data_free_idx), sv2v_cast_1B5F4(oup_data_free_idx), 1'b0};
					// Trace: design.sv:27213:21
					linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (oup_data_free_idx * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = {inp_data_i, sv2v_cast_1B5F4(1'sb0), 1'b0};
				end
				else if (no_in_id_match) begin
					begin
						// Trace: design.sv:27220:21
						if (oup_ht_popped) begin
							// Trace: design.sv:27221:25
							head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (match_out_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] = {sv2v_cast_64419(inp_id_i), sv2v_cast_1B5F4(oup_data_free_idx), sv2v_cast_1B5F4(oup_data_free_idx), 1'b0};
							// Trace: design.sv:27227:25
							linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (oup_data_free_idx * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = {inp_data_i, sv2v_cast_1B5F4(1'sb0), 1'b0};
						end
						else
							// Trace: design.sv:27233:25
							if (oup_data_popped) begin
								// Trace: design.sv:27234:27
								head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (head_tail_free_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] = {sv2v_cast_64419(inp_id_i), sv2v_cast_1B5F4(oup_data_free_idx), sv2v_cast_1B5F4(oup_data_free_idx), 1'b0};
								// Trace: design.sv:27240:27
								linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (oup_data_free_idx * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = {inp_data_i, sv2v_cast_1B5F4(1'sb0), 1'b0};
							end
							else begin
								// Trace: design.sv:27246:29
								head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (head_tail_free_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] = {sv2v_cast_64419(inp_id_i), sv2v_cast_1B5F4(linked_data_free_idx), sv2v_cast_1B5F4(linked_data_free_idx), 1'b0};
								// Trace: design.sv:27252:29
								linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (linked_data_free_idx * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = {inp_data_i, sv2v_cast_1B5F4(1'sb0), 1'b0};
							end
					end
				end
				else
					// Trace: design.sv:27261:21
					if (oup_data_popped) begin
						// Trace: design.sv:27262:25
						linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] = oup_data_free_idx;
						// Trace: design.sv:27263:25
						head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] = oup_data_free_idx;
						// Trace: design.sv:27264:25
						linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (oup_data_free_idx * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = {inp_data_i, sv2v_cast_1B5F4(1'sb0), 1'b0};
					end
					else begin
						// Trace: design.sv:27270:25
						linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? (head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : ((32 + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] = linked_data_free_idx;
						// Trace: design.sv:27271:25
						head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? (match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0)) : (((match_in_idx * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))) + ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? LdIdxWidth + 0 : (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) - (LdIdxWidth + 0))) + ((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))) - 1)-:((LdIdxWidth + 0) >= 1 ? LdIdxWidth + 0 : 2 - (LdIdxWidth + 0))] = linked_data_free_idx;
						// Trace: design.sv:27272:25
						linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (linked_data_free_idx * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] = {inp_data_i, sv2v_cast_1B5F4(1'sb0), 1'b0};
					end
			end
		end
	end
	// Trace: design.sv:27284:5
	genvar _gv_i_24;
	generate
		for (_gv_i_24 = 0; _gv_i_24 < CAPACITY; _gv_i_24 = _gv_i_24 + 1) begin : gen_lookup
			localparam i = _gv_i_24;
			// Trace: design.sv:27285:9
			reg [31:0] exists_match_bits;
			genvar _gv_j_8;
			for (_gv_j_8 = 0; _gv_j_8 < 32; _gv_j_8 = _gv_j_8 + 1) begin : gen_mask
				localparam j = _gv_j_8;
				// Trace: design.sv:27287:13
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:27288:17
					if (linked_data_q[(i * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0)])
						// Trace: design.sv:27289:21
						exists_match_bits[j] = 1'b0;
					else
						// Trace: design.sv:27291:21
						if (!exists_mask_i[j])
							// Trace: design.sv:27292:25
							exists_match_bits[j] = 1'b1;
						else
							// Trace: design.sv:27294:25
							exists_match_bits[j] = linked_data_q[(i * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? (32 + (LdIdxWidth + 0)) - (31 - j) : ((32 + LdIdxWidth) + 0) - ((32 + (LdIdxWidth + 0)) - (31 - j)))] == exists_data_i[j];
				end
			end
			// Trace: design.sv:27299:9
			assign exists_match[i] = &exists_match_bits;
		end
	endgenerate
	// Trace: design.sv:27301:5
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:27302:9
		exists_gnt_o = 1'b0;
		// Trace: design.sv:27303:9
		exists_o = 1'sb0;
		// Trace: design.sv:27304:9
		if (exists_req_i) begin
			// Trace: design.sv:27305:13
			exists_gnt_o = 1'b1;
			// Trace: design.sv:27306:13
			exists_o = |exists_match;
		end
	end
	// Trace: design.sv:27311:5
	genvar _gv_i_25;
	generate
		for (_gv_i_25 = 0; _gv_i_25 < HtCapacity; _gv_i_25 = _gv_i_25 + 1) begin : gen_ht_ffs
			localparam i = _gv_i_25;
			// Trace: design.sv:27312:9
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:27313:13
				if (!rst_ni)
					// Trace: design.sv:27314:17
					head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] <= {sv2v_cast_37B7D(1'sb0), sv2v_cast_D5FF0(1'sb0), sv2v_cast_D5FF0(1'sb0), 1'b1};
				else
					// Trace: design.sv:27316:17
					head_tail_q[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))] <= head_tail_d[((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? 0 : ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) + (i * ((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0)))+:((((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0) >= 0 ? ((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 1 : 1 - (((ID_WIDTH + LdIdxWidth) + LdIdxWidth) + 0))];
		end
	endgenerate
	// Trace: design.sv:27320:5
	genvar _gv_i_26;
	generate
		for (_gv_i_26 = 0; _gv_i_26 < CAPACITY; _gv_i_26 = _gv_i_26 + 1) begin : gen_data_ffs
			localparam i = _gv_i_26;
			// Trace: design.sv:27321:9
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:27322:13
				if (!rst_ni) begin
					// Trace: design.sv:27324:17
					linked_data_q[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (i * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] <= 1'sb0;
					// Trace: design.sv:27325:17
					linked_data_q[(i * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))) + (((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0)] <= 1'b1;
				end
				else
					// Trace: design.sv:27327:17
					linked_data_q[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (i * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))] <= linked_data_d[(((32 + LdIdxWidth) + 0) >= 0 ? 0 : (32 + LdIdxWidth) + 0) + (i * (((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0)))+:(((32 + LdIdxWidth) + 0) >= 0 ? (32 + LdIdxWidth) + 1 : 1 - ((32 + LdIdxWidth) + 0))];
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module stream_to_mem (
	clk_i,
	rst_ni,
	req_i,
	req_valid_i,
	req_ready_o,
	resp_o,
	resp_valid_o,
	resp_ready_i,
	mem_req_o,
	mem_req_valid_o,
	mem_req_ready_i,
	mem_resp_i,
	mem_resp_valid_i
);
	reg _sv2v_0;
	// Trace: design.sv:27363:26
	// removed localparam type mem_req_t
	// Trace: design.sv:27365:26
	// removed localparam type mem_resp_t
	// Trace: design.sv:27371:13
	parameter [31:0] BufDepth = 32'd1;
	// Trace: design.sv:27374:3
	input wire clk_i;
	// Trace: design.sv:27376:3
	input wire rst_ni;
	// Trace: design.sv:27378:3
	input wire req_i;
	// Trace: design.sv:27380:3
	input wire req_valid_i;
	// Trace: design.sv:27382:3
	output wire req_ready_o;
	// Trace: design.sv:27384:3
	output wire resp_o;
	// Trace: design.sv:27386:3
	output wire resp_valid_o;
	// Trace: design.sv:27388:3
	input wire resp_ready_i;
	// Trace: design.sv:27390:3
	output wire mem_req_o;
	// Trace: design.sv:27392:3
	output wire mem_req_valid_o;
	// Trace: design.sv:27394:3
	input wire mem_req_ready_i;
	// Trace: design.sv:27396:3
	input wire mem_resp_i;
	// Trace: design.sv:27398:3
	input wire mem_resp_valid_i;
	// Trace: design.sv:27401:3
	// removed localparam type cnt_t
	// Trace: design.sv:27403:3
	reg [$clog2(BufDepth + 1):0] cnt_d;
	reg [$clog2(BufDepth + 1):0] cnt_q;
	// Trace: design.sv:27404:3
	wire buf_ready;
	wire req_ready;
	// Trace: design.sv:27407:3
	generate
		if (BufDepth > 0) begin : gen_buf
			// Trace: design.sv:27409:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:27410:7
				cnt_d = cnt_q;
				// Trace: design.sv:27411:7
				if (req_valid_i && req_ready_o)
					// Trace: design.sv:27412:9
					cnt_d = cnt_d + 1;
				if (resp_valid_o && resp_ready_i)
					// Trace: design.sv:27415:9
					cnt_d = cnt_d - 1;
			end
			// Trace: design.sv:27421:5
			assign req_ready = (cnt_q < BufDepth) | (resp_valid_o & resp_ready_i);
			// Trace: design.sv:27424:5
			assign req_ready_o = mem_req_ready_i & req_ready;
			// Trace: design.sv:27425:5
			assign mem_req_valid_o = req_valid_i & req_ready;
			// Trace: design.sv:27428:5
			stream_fifo_10183 #(
				.FALL_THROUGH(1'b1),
				.DEPTH(BufDepth)
			) i_resp_buf(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(1'b0),
				.data_i(mem_resp_i),
				.valid_i(mem_resp_valid_i),
				.ready_o(buf_ready),
				.data_o(resp_o),
				.valid_o(resp_valid_o),
				.ready_i(resp_ready_i),
				.usage_o()
			);
			// Trace: macro expansion of FF at design.sv:27447:86
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FF at design.sv:27447:174
				if (!rst_ni)
					// Trace: macro expansion of FF at design.sv:27447:262
					cnt_q <= 1'sb0;
				else
					// Trace: macro expansion of FF at design.sv:27447:434
					cnt_q <= cnt_d;
		end
		else begin : gen_no_buf
			// Trace: design.sv:27451:5
			assign mem_req_valid_o = req_valid_i;
			// Trace: design.sv:27452:5
			assign resp_valid_o = (mem_req_valid_o & mem_req_ready_i) & mem_resp_valid_i;
			// Trace: design.sv:27453:5
			assign req_ready_o = resp_ready_i & resp_valid_o;
			// Trace: design.sv:27456:5
			assign resp_o = mem_resp_i;
		end
	endgenerate
	// Trace: design.sv:27460:3
	assign mem_req_o = req_i;
	initial _sv2v_0 = 0;
endmodule
module stream_arbiter_flushable_8B6F2 (
	clk_i,
	rst_ni,
	flush_i,
	inp_data_i,
	inp_valid_i,
	inp_ready_o,
	oup_data_o,
	oup_valid_o,
	oup_ready_i
);
	// Trace: design.sv:27495:25
	// removed localparam type DATA_T
	// Trace: design.sv:27496:15
	parameter integer N_INP = -1;
	// Trace: design.sv:27497:25
	parameter ARBITER = "rr";
	// Trace: design.sv:27499:5
	input wire clk_i;
	// Trace: design.sv:27500:5
	input wire rst_ni;
	// Trace: design.sv:27501:5
	input wire flush_i;
	// Trace: design.sv:27503:5
	input wire [N_INP - 1:0] inp_data_i;
	// Trace: design.sv:27504:5
	input wire [N_INP - 1:0] inp_valid_i;
	// Trace: design.sv:27505:5
	output wire [N_INP - 1:0] inp_ready_o;
	// Trace: design.sv:27507:5
	output wire oup_data_o;
	// Trace: design.sv:27508:5
	output wire oup_valid_o;
	// Trace: design.sv:27509:5
	input wire oup_ready_i;
	// Trace: design.sv:27512:3
	generate
		if (ARBITER == "rr") begin : gen_rr_arb
			// Trace: design.sv:27513:5
			localparam [31:0] sv2v_uu_i_arbiter_NumIn = N_INP;
			localparam [31:0] sv2v_uu_i_arbiter_IdxWidth = (sv2v_uu_i_arbiter_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_arbiter_NumIn)) : 32'd1);
			// removed localparam type sv2v_uu_i_arbiter_idx_t
			// removed localparam type sv2v_uu_i_arbiter_rr_i
			localparam [sv2v_uu_i_arbiter_IdxWidth - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
			rr_arb_tree_93F52 #(
				.NumIn(N_INP),
				.ExtPrio(1'b0),
				.AxiVldRdy(1'b1),
				.LockIn(1'b1)
			) i_arbiter(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
				.req_i(inp_valid_i),
				.gnt_o(inp_ready_o),
				.data_i(inp_data_i),
				.gnt_i(oup_ready_i),
				.req_o(oup_valid_o),
				.data_o(oup_data_o),
				.idx_o()
			);
		end
		else if (ARBITER == "prio") begin : gen_prio_arb
			// Trace: design.sv:27534:5
			localparam [31:0] sv2v_uu_i_arbiter_NumIn = N_INP;
			localparam [31:0] sv2v_uu_i_arbiter_IdxWidth = (sv2v_uu_i_arbiter_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_arbiter_NumIn)) : 32'd1);
			// removed localparam type sv2v_uu_i_arbiter_idx_t
			// removed localparam type sv2v_uu_i_arbiter_rr_i
			localparam [sv2v_uu_i_arbiter_IdxWidth - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
			rr_arb_tree_93F52 #(
				.NumIn(N_INP),
				.ExtPrio(1'b1),
				.AxiVldRdy(1'b1),
				.LockIn(1'b1)
			) i_arbiter(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
				.req_i(inp_valid_i),
				.gnt_o(inp_ready_o),
				.data_i(inp_data_i),
				.gnt_i(oup_ready_i),
				.req_o(oup_valid_o),
				.data_o(oup_data_o),
				.idx_o()
			);
		end
		else begin : gen_arb_error
			// Trace: design.sv:27556:5
			$fatal(1, "Invalid value for parameter 'ARBITER'!");
		end
	endgenerate
endmodule
module stream_fifo_optimal_wrap (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	usage_o,
	data_i,
	valid_i,
	ready_o,
	data_o,
	valid_o,
	ready_i
);
	// Trace: design.sv:27572:15
	parameter [31:0] Depth = 32'd8;
	// Trace: design.sv:27574:20
	// removed localparam type type_t
	// Trace: design.sv:27576:15
	parameter [0:0] PrintInfo = 1'b0;
	// Trace: design.sv:27578:15
	parameter [31:0] AddrDepth = (Depth > 32'd1 ? $clog2(Depth) : 32'd1);
	// Trace: design.sv:27580:5
	input wire clk_i;
	// Trace: design.sv:27581:5
	input wire rst_ni;
	// Trace: design.sv:27582:5
	input wire flush_i;
	// Trace: design.sv:27583:5
	input wire testmode_i;
	// Trace: design.sv:27584:5
	output wire [AddrDepth - 1:0] usage_o;
	// Trace: design.sv:27586:5
	input wire data_i;
	// Trace: design.sv:27587:5
	input wire valid_i;
	// Trace: design.sv:27588:5
	output wire ready_o;
	// Trace: design.sv:27590:5
	output wire data_o;
	// Trace: design.sv:27591:5
	output wire valid_o;
	// Trace: design.sv:27592:5
	input wire ready_i;
	// Trace: design.sv:27600:5
	generate
		if (Depth < 32'd2) begin : gen_fatal
			// Trace: design.sv:27601:9
			initial begin
				// Trace: design.sv:27602:13
				$fatal(1, "FIFO of depth %d does not make any sense!", Depth);
			end
		end
	endgenerate
	// Trace: design.sv:27611:5
	generate
		if (Depth == 32'd2) begin : gen_spill
			if (PrintInfo) begin : gen_info
				// Trace: design.sv:27616:13
				initial begin
					// Trace: design.sv:27617:17
					$display("[%m] Instantiate spill register (of depth %d)", Depth);
				end
			end
			// Trace: design.sv:27623:9
			spill_register_flushable_D072E #(.Bypass(1'b0)) i_spill_register_flushable(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.valid_i(valid_i),
				.ready_o(ready_o),
				.data_i(data_i),
				.valid_o(valid_o),
				.ready_i(ready_i),
				.data_o(data_o)
			);
			// Trace: design.sv:27639:9
			assign usage_o = 1'sbx;
		end
	endgenerate
	// Trace: design.sv:27647:5
	generate
		if (Depth > 32'd2) begin : gen_fifo
			if (PrintInfo) begin : gen_info
				// Trace: design.sv:27652:13
				initial begin
					// Trace: design.sv:27653:17
					$info("[%m] Instantiate stream FIFO of depth %d", Depth);
				end
			end
			// Trace: design.sv:27659:9
			stream_fifo_10183 #(.DEPTH(Depth)) i_stream_fifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.testmode_i(testmode_i),
				.usage_o(usage_o),
				.data_i(data_i),
				.valid_i(valid_i),
				.ready_o(ready_o),
				.data_o(data_o),
				.valid_o(valid_o),
				.ready_i(ready_i)
			);
		end
	endgenerate
endmodule
module stream_register (
	clk_i,
	rst_ni,
	clr_i,
	testmode_i,
	valid_i,
	ready_o,
	data_i,
	valid_o,
	ready_i,
	data_o
);
	// Trace: design.sv:27694:20
	// removed localparam type T
	// Trace: design.sv:27696:5
	input wire clk_i;
	// Trace: design.sv:27697:5
	input wire rst_ni;
	// Trace: design.sv:27698:5
	input wire clr_i;
	// Trace: design.sv:27699:5
	input wire testmode_i;
	// Trace: design.sv:27701:5
	input wire valid_i;
	// Trace: design.sv:27702:5
	output wire ready_o;
	// Trace: design.sv:27703:5
	input wire data_i;
	// Trace: design.sv:27705:5
	output reg valid_o;
	// Trace: design.sv:27706:5
	input wire ready_i;
	// Trace: design.sv:27707:5
	output reg data_o;
	// Trace: design.sv:27710:5
	wire reg_ena;
	// Trace: design.sv:27711:5
	assign ready_o = ready_i | ~valid_o;
	// Trace: design.sv:27712:5
	assign reg_ena = valid_i & ready_o;
	// Trace: macro expansion of FFLARNC at design.sv:27714:291
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFLARNC at design.sv:27714:369
		if (!rst_ni)
			// Trace: macro expansion of FFLARNC at design.sv:27714:447
			valid_o <= 1'b0;
		else
			// Trace: macro expansion of FFLARNC at design.sv:27714:599
			if (clr_i)
				// Trace: macro expansion of FFLARNC at design.sv:27714:677
				valid_o <= 1'b0;
			else if (ready_o)
				// Trace: macro expansion of FFLARNC at design.sv:27714:829
				valid_o <= valid_i;
	// Trace: macro expansion of FFLARNC at design.sv:27715:291
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFLARNC at design.sv:27715:369
		if (!rst_ni)
			// Trace: macro expansion of FFLARNC at design.sv:27715:447
			data_o <= 1'sb0;
		else
			// Trace: macro expansion of FFLARNC at design.sv:27715:599
			if (clr_i)
				// Trace: macro expansion of FFLARNC at design.sv:27715:677
				data_o <= 1'sb0;
			else if (reg_ena)
				// Trace: macro expansion of FFLARNC at design.sv:27715:829
				data_o <= data_i;
endmodule
module stream_xbar_09F43_1A7A9 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	data_i,
	sel_i,
	valid_i,
	ready_o,
	data_o,
	idx_o,
	valid_o,
	ready_i
);
	// removed localparam type payload_t_DataWidth_type
	// removed localparam type payload_t_IdxWidth_type
	// removed localparam type payload_t_i_stream_xbar_sv2v_pfunc_944F6_type
	parameter [31:0] payload_t_DataWidth = 0;
	parameter [31:0] payload_t_IdxWidth = 0;
	parameter integer payload_t_i_stream_xbar_sv2v_pfunc_944F6 = 0;
	reg _sv2v_0;
	// Trace: design.sv:27735:13
	parameter [31:0] NumInp = 32'd0;
	// Trace: design.sv:27737:13
	parameter [31:0] NumOut = 32'd0;
	// Trace: design.sv:27739:13
	parameter [31:0] DataWidth = 32'd1;
	// Trace: design.sv:27741:26
	// removed localparam type payload_t
	// Trace: design.sv:27743:13
	parameter [0:0] OutSpillReg = 1'b0;
	// Trace: design.sv:27745:13
	parameter [31:0] ExtPrio = 1'b0;
	// Trace: design.sv:27748:13
	parameter [31:0] AxiVldRdy = 1'b1;
	// Trace: design.sv:27752:13
	parameter [31:0] LockIn = 1'b1;
	// Trace: design.sv:27756:13
	parameter [31:0] SelWidth = (NumOut > 32'd1 ? $unsigned($clog2(NumOut)) : 32'd1);
	// Trace: design.sv:27760:18
	// removed localparam type sel_oup_t
	// Trace: design.sv:27764:13
	parameter [31:0] IdxWidth = (NumInp > 32'd1 ? $unsigned($clog2(NumInp)) : 32'd1);
	// Trace: design.sv:27768:18
	// removed localparam type idx_inp_t
	// Trace: design.sv:27771:3
	input wire clk_i;
	// Trace: design.sv:27773:3
	input wire rst_ni;
	// Trace: design.sv:27778:3
	input wire flush_i;
	// Trace: design.sv:27781:3
	input wire [(NumOut * IdxWidth) - 1:0] rr_i;
	// Trace: design.sv:27784:3
	input wire [(NumInp * ((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth)) - 1:0] data_i;
	// Trace: design.sv:27787:3
	input wire [(NumInp * SelWidth) - 1:0] sel_i;
	// Trace: design.sv:27789:3
	input wire [NumInp - 1:0] valid_i;
	// Trace: design.sv:27791:3
	output wire [NumInp - 1:0] ready_o;
	// Trace: design.sv:27793:3
	output reg [(NumOut * ((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth)) - 1:0] data_o;
	// Trace: design.sv:27795:3
	output reg [(NumOut * IdxWidth) - 1:0] idx_o;
	// Trace: design.sv:27797:3
	output wire [NumOut - 1:0] valid_o;
	// Trace: design.sv:27799:3
	input wire [NumOut - 1:0] ready_i;
	// Trace: design.sv:27801:3
	// removed localparam type spill_data_t
	// Trace: design.sv:27806:3
	wire [(NumInp * NumOut) - 1:0] inp_valid;
	// Trace: design.sv:27807:3
	wire [(NumInp * NumOut) - 1:0] inp_ready;
	// Trace: design.sv:27809:3
	wire [((NumOut * NumInp) * ((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth)) - 1:0] out_data;
	// Trace: design.sv:27810:3
	wire [(NumOut * NumInp) - 1:0] out_valid;
	// Trace: design.sv:27811:3
	wire [(NumOut * NumInp) - 1:0] out_ready;
	// Trace: design.sv:27814:3
	genvar _gv_i_27;
	generate
		for (_gv_i_27 = 0; $unsigned(_gv_i_27) < NumInp; _gv_i_27 = _gv_i_27 + 1) begin : gen_inps
			localparam i = _gv_i_27;
			// Trace: design.sv:27815:5
			stream_demux #(.N_OUP(NumOut)) i_stream_demux(
				.inp_valid_i(valid_i[i]),
				.inp_ready_o(ready_o[i]),
				.oup_sel_i(sel_i[i * SelWidth+:SelWidth]),
				.oup_valid_o(inp_valid[i * NumOut+:NumOut]),
				.oup_ready_i(inp_ready[i * NumOut+:NumOut])
			);
			genvar _gv_j_9;
			for (_gv_j_9 = 0; $unsigned(_gv_j_9) < NumOut; _gv_j_9 = _gv_j_9 + 1) begin : gen_cross
				localparam j = _gv_j_9;
				// Trace: design.sv:27828:7
				assign out_data[((j * NumInp) + i) * ((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth)+:(payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth] = data_i[i * ((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth)+:(payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth];
				// Trace: design.sv:27830:7
				assign out_valid[(j * NumInp) + i] = inp_valid[(i * NumOut) + j];
				// Trace: design.sv:27831:7
				assign inp_ready[(i * NumOut) + j] = out_ready[(j * NumInp) + i];
			end
		end
	endgenerate
	// Trace: design.sv:27836:3
	genvar _gv_j_10;
	generate
		for (_gv_j_10 = 0; $unsigned(_gv_j_10) < NumOut; _gv_j_10 = _gv_j_10 + 1) begin : gen_outs
			localparam j = _gv_j_10;
			// Trace: design.sv:27837:5
			wire [(((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + IdxWidth) - 1:0] arb;
			// Trace: design.sv:27838:5
			wire arb_valid;
			wire arb_ready;
			// Trace: design.sv:27840:5
			rr_arb_tree_D7936_86F21 #(
				.DataType_payload_t_DataWidth(payload_t_DataWidth),
				.DataType_payload_t_IdxWidth(payload_t_IdxWidth),
				.DataType_payload_t_i_stream_xbar_sv2v_pfunc_944F6(payload_t_i_stream_xbar_sv2v_pfunc_944F6),
				.NumIn(NumInp),
				.ExtPrio(ExtPrio),
				.AxiVldRdy(AxiVldRdy),
				.LockIn(LockIn)
			) i_rr_arb_tree(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.rr_i(rr_i[j * IdxWidth+:IdxWidth]),
				.req_i(out_valid[j * NumInp+:NumInp]),
				.gnt_o(out_ready[j * NumInp+:NumInp]),
				.data_i(out_data[((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) * (j * NumInp)+:((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) * NumInp]),
				.req_o(arb_valid),
				.gnt_i(arb_ready),
				.data_o(arb[((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + (IdxWidth - 1)-:((((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + (IdxWidth - 1)) >= (IdxWidth + 0) ? ((((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + (IdxWidth - 1)) - (IdxWidth + 0)) + 1 : ((IdxWidth + 0) - (((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + (IdxWidth - 1))) + 1)]),
				.idx_o(arb[IdxWidth - 1-:IdxWidth])
			);
			// Trace: design.sv:27860:5
			wire [(((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + IdxWidth) - 1:0] spill;
			// Trace: design.sv:27862:5
			spill_register_0D540_46F20 #(
				.T_IdxWidth(IdxWidth),
				.T_payload_t_DataWidth(payload_t_DataWidth),
				.T_payload_t_IdxWidth(payload_t_IdxWidth),
				.T_payload_t_i_stream_xbar_sv2v_pfunc_944F6(payload_t_i_stream_xbar_sv2v_pfunc_944F6),
				.Bypass(!OutSpillReg)
			) i_spill_register(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.valid_i(arb_valid),
				.ready_o(arb_ready),
				.data_i(arb),
				.valid_o(valid_o[j]),
				.ready_i(ready_i[j]),
				.data_o(spill)
			);
			// Trace: design.sv:27876:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:27877:7
				data_o[j * ((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth)+:(payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth] = spill[((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + (IdxWidth - 1)-:((((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + (IdxWidth - 1)) >= (IdxWidth + 0) ? ((((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + (IdxWidth - 1)) - (IdxWidth + 0)) + 1 : ((IdxWidth + 0) - (((payload_t_i_stream_xbar_sv2v_pfunc_944F6 + payload_t_DataWidth) + payload_t_IdxWidth) + (IdxWidth - 1))) + 1)];
				// Trace: design.sv:27878:7
				idx_o[j * IdxWidth+:IdxWidth] = spill[IdxWidth - 1-:IdxWidth];
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module stream_xbar_67930_B7325 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	data_i,
	sel_i,
	valid_i,
	ready_o,
	data_o,
	idx_o,
	valid_o,
	ready_i
);
	// removed localparam type payload_t_DataWidth_type
	parameter [31:0] payload_t_DataWidth = 0;
	reg _sv2v_0;
	// Trace: design.sv:27735:13
	parameter [31:0] NumInp = 32'd0;
	// Trace: design.sv:27737:13
	parameter [31:0] NumOut = 32'd0;
	// Trace: design.sv:27739:13
	parameter [31:0] DataWidth = 32'd1;
	// Trace: design.sv:27741:26
	// removed localparam type payload_t
	// Trace: design.sv:27743:13
	parameter [0:0] OutSpillReg = 1'b0;
	// Trace: design.sv:27745:13
	parameter [31:0] ExtPrio = 1'b0;
	// Trace: design.sv:27748:13
	parameter [31:0] AxiVldRdy = 1'b1;
	// Trace: design.sv:27752:13
	parameter [31:0] LockIn = 1'b1;
	// Trace: design.sv:27756:13
	parameter [31:0] SelWidth = (NumOut > 32'd1 ? $unsigned($clog2(NumOut)) : 32'd1);
	// Trace: design.sv:27760:18
	// removed localparam type sel_oup_t
	// Trace: design.sv:27764:13
	parameter [31:0] IdxWidth = (NumInp > 32'd1 ? $unsigned($clog2(NumInp)) : 32'd1);
	// Trace: design.sv:27768:18
	// removed localparam type idx_inp_t
	// Trace: design.sv:27771:3
	input wire clk_i;
	// Trace: design.sv:27773:3
	input wire rst_ni;
	// Trace: design.sv:27778:3
	input wire flush_i;
	// Trace: design.sv:27781:3
	input wire [(NumOut * IdxWidth) - 1:0] rr_i;
	// Trace: design.sv:27784:3
	input wire [(NumInp * payload_t_DataWidth) - 1:0] data_i;
	// Trace: design.sv:27787:3
	input wire [(NumInp * SelWidth) - 1:0] sel_i;
	// Trace: design.sv:27789:3
	input wire [NumInp - 1:0] valid_i;
	// Trace: design.sv:27791:3
	output wire [NumInp - 1:0] ready_o;
	// Trace: design.sv:27793:3
	output reg [(NumOut * payload_t_DataWidth) - 1:0] data_o;
	// Trace: design.sv:27795:3
	output reg [(NumOut * IdxWidth) - 1:0] idx_o;
	// Trace: design.sv:27797:3
	output wire [NumOut - 1:0] valid_o;
	// Trace: design.sv:27799:3
	input wire [NumOut - 1:0] ready_i;
	// Trace: design.sv:27801:3
	// removed localparam type spill_data_t
	// Trace: design.sv:27806:3
	wire [(NumInp * NumOut) - 1:0] inp_valid;
	// Trace: design.sv:27807:3
	wire [(NumInp * NumOut) - 1:0] inp_ready;
	// Trace: design.sv:27809:3
	wire [((NumOut * NumInp) * payload_t_DataWidth) - 1:0] out_data;
	// Trace: design.sv:27810:3
	wire [(NumOut * NumInp) - 1:0] out_valid;
	// Trace: design.sv:27811:3
	wire [(NumOut * NumInp) - 1:0] out_ready;
	// Trace: design.sv:27814:3
	genvar _gv_i_27;
	generate
		for (_gv_i_27 = 0; $unsigned(_gv_i_27) < NumInp; _gv_i_27 = _gv_i_27 + 1) begin : gen_inps
			localparam i = _gv_i_27;
			// Trace: design.sv:27815:5
			stream_demux #(.N_OUP(NumOut)) i_stream_demux(
				.inp_valid_i(valid_i[i]),
				.inp_ready_o(ready_o[i]),
				.oup_sel_i(sel_i[i * SelWidth+:SelWidth]),
				.oup_valid_o(inp_valid[i * NumOut+:NumOut]),
				.oup_ready_i(inp_ready[i * NumOut+:NumOut])
			);
			genvar _gv_j_9;
			for (_gv_j_9 = 0; $unsigned(_gv_j_9) < NumOut; _gv_j_9 = _gv_j_9 + 1) begin : gen_cross
				localparam j = _gv_j_9;
				// Trace: design.sv:27828:7
				assign out_data[((j * NumInp) + i) * payload_t_DataWidth+:payload_t_DataWidth] = data_i[i * payload_t_DataWidth+:payload_t_DataWidth];
				// Trace: design.sv:27830:7
				assign out_valid[(j * NumInp) + i] = inp_valid[(i * NumOut) + j];
				// Trace: design.sv:27831:7
				assign inp_ready[(i * NumOut) + j] = out_ready[(j * NumInp) + i];
			end
		end
	endgenerate
	// Trace: design.sv:27836:3
	genvar _gv_j_10;
	generate
		for (_gv_j_10 = 0; $unsigned(_gv_j_10) < NumOut; _gv_j_10 = _gv_j_10 + 1) begin : gen_outs
			localparam j = _gv_j_10;
			// Trace: design.sv:27837:5
			wire [(payload_t_DataWidth + IdxWidth) - 1:0] arb;
			// Trace: design.sv:27838:5
			wire arb_valid;
			wire arb_ready;
			// Trace: design.sv:27840:5
			rr_arb_tree_0C7DB_08AEF #(
				.DataType_payload_t_DataWidth(payload_t_DataWidth),
				.NumIn(NumInp),
				.ExtPrio(ExtPrio),
				.AxiVldRdy(AxiVldRdy),
				.LockIn(LockIn)
			) i_rr_arb_tree(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.rr_i(rr_i[j * IdxWidth+:IdxWidth]),
				.req_i(out_valid[j * NumInp+:NumInp]),
				.gnt_o(out_ready[j * NumInp+:NumInp]),
				.data_i(out_data[payload_t_DataWidth * (j * NumInp)+:payload_t_DataWidth * NumInp]),
				.req_o(arb_valid),
				.gnt_i(arb_ready),
				.data_o(arb[payload_t_DataWidth + (IdxWidth - 1)-:((payload_t_DataWidth + (IdxWidth - 1)) >= (IdxWidth + 0) ? ((payload_t_DataWidth + (IdxWidth - 1)) - (IdxWidth + 0)) + 1 : ((IdxWidth + 0) - (payload_t_DataWidth + (IdxWidth - 1))) + 1)]),
				.idx_o(arb[IdxWidth - 1-:IdxWidth])
			);
			// Trace: design.sv:27860:5
			wire [(payload_t_DataWidth + IdxWidth) - 1:0] spill;
			// Trace: design.sv:27862:5
			spill_register_1C0C7_8C0C0 #(
				.T_IdxWidth(IdxWidth),
				.T_payload_t_DataWidth(payload_t_DataWidth),
				.Bypass(!OutSpillReg)
			) i_spill_register(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.valid_i(arb_valid),
				.ready_o(arb_ready),
				.data_i(arb),
				.valid_o(valid_o[j]),
				.ready_i(ready_i[j]),
				.data_o(spill)
			);
			// Trace: design.sv:27876:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:27877:7
				data_o[j * payload_t_DataWidth+:payload_t_DataWidth] = spill[payload_t_DataWidth + (IdxWidth - 1)-:((payload_t_DataWidth + (IdxWidth - 1)) >= (IdxWidth + 0) ? ((payload_t_DataWidth + (IdxWidth - 1)) - (IdxWidth + 0)) + 1 : ((IdxWidth + 0) - (payload_t_DataWidth + (IdxWidth - 1))) + 1)];
				// Trace: design.sv:27878:7
				idx_o[j * IdxWidth+:IdxWidth] = spill[IdxWidth - 1-:IdxWidth];
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module cdc_fifo_gray_clearable (
	src_rst_ni,
	src_clk_i,
	src_clear_i,
	src_clear_pending_o,
	src_data_i,
	src_valid_i,
	src_ready_o,
	dst_rst_ni,
	dst_clk_i,
	dst_clear_i,
	dst_clear_pending_o,
	dst_data_o,
	dst_valid_o,
	dst_ready_i
);
	// Trace: design.sv:28021:13
	parameter [31:0] WIDTH = 1;
	// Trace: design.sv:28023:18
	// removed localparam type T
	// Trace: design.sv:28025:13
	parameter signed [31:0] LOG_DEPTH = 3;
	// Trace: design.sv:28031:13
	parameter signed [31:0] SYNC_STAGES = 3;
	// Trace: design.sv:28032:13
	parameter signed [31:0] CLEAR_ON_ASYNC_RESET = 1;
	// Trace: design.sv:28034:3
	input wire src_rst_ni;
	// Trace: design.sv:28035:3
	input wire src_clk_i;
	// Trace: design.sv:28036:3
	input wire src_clear_i;
	// Trace: design.sv:28037:3
	output wire src_clear_pending_o;
	// Trace: design.sv:28038:3
	input wire [WIDTH - 1:0] src_data_i;
	// Trace: design.sv:28039:3
	input wire src_valid_i;
	// Trace: design.sv:28040:3
	output wire src_ready_o;
	// Trace: design.sv:28042:3
	input wire dst_rst_ni;
	// Trace: design.sv:28043:3
	input wire dst_clk_i;
	// Trace: design.sv:28044:3
	input wire dst_clear_i;
	// Trace: design.sv:28045:3
	output wire dst_clear_pending_o;
	// Trace: design.sv:28046:3
	output wire [WIDTH - 1:0] dst_data_o;
	// Trace: design.sv:28047:3
	output wire dst_valid_o;
	// Trace: design.sv:28048:3
	input wire dst_ready_i;
	// Trace: design.sv:28051:3
	wire s_src_clear_req;
	// Trace: design.sv:28052:3
	reg s_src_clear_ack_q;
	// Trace: design.sv:28053:3
	wire s_src_ready;
	// Trace: design.sv:28054:3
	wire s_src_isolate_req;
	// Trace: design.sv:28055:3
	reg s_src_isolate_ack_q;
	// Trace: design.sv:28056:3
	wire s_dst_clear_req;
	// Trace: design.sv:28057:3
	reg s_dst_clear_ack_q;
	// Trace: design.sv:28058:3
	wire s_dst_valid;
	// Trace: design.sv:28059:3
	wire s_dst_isolate_req;
	// Trace: design.sv:28060:3
	reg s_dst_isolate_ack_q;
	// Trace: design.sv:28063:3
	wire [((2 ** LOG_DEPTH) * WIDTH) - 1:0] async_data;
	// Trace: design.sv:28064:3
	wire [LOG_DEPTH:0] async_wptr;
	// Trace: design.sv:28065:3
	wire [LOG_DEPTH:0] async_rptr;
	// Trace: design.sv:28067:3
	generate
		if (CLEAR_ON_ASYNC_RESET) begin : gen_elaboration_assertion
			if (SYNC_STAGES < 3) begin : genblk1
				// Trace: design.sv:28069:7
				$error("The clearable CDC FIFO with async reset synchronization requires at least", "3 synchronizer stages for the FIFO.");
			end
		end
		else begin : gen_elaboration_assertion
			if (SYNC_STAGES < 2) begin : gen_elaboration_assertion
				// Trace: design.sv:28073:7
				$error("A minimum of 2 synchronizer stages is required for proper functionality.");
			end
		end
	endgenerate
	// Trace: design.sv:28077:3
	generate
		if ((2 * SYNC_STAGES) > (2 ** LOG_DEPTH)) begin : gen_elaboration_assertion2
			// Trace: design.sv:28078:5
			$warning("The FIFOs depth of %0d is insufficient to completely hide the latency of", " %0d SYNC_STAGES. The FIFO will stall in the case where f_src ~= f_dst. ", "It is reccomended to increase the FIFO's log depth to at least %0d.", 2 ** LOG_DEPTH, SYNC_STAGES, $clog2(2 * SYNC_STAGES));
		end
	endgenerate
	// Trace: design.sv:28086:3
	cdc_fifo_gray_src_clearable_0070C_CFA0B #(
		.T_WIDTH(WIDTH),
		.LOG_DEPTH(LOG_DEPTH),
		.SYNC_STAGES(SYNC_STAGES)
	) i_src(
		.src_rst_ni(src_rst_ni),
		.src_clk_i(src_clk_i),
		.src_clear_i(s_src_clear_req),
		.src_data_i(src_data_i),
		.src_valid_i(src_valid_i & !s_src_isolate_req),
		.src_ready_o(s_src_ready),
		.async_data_o(async_data),
		.async_wptr_o(async_wptr),
		.async_rptr_i(async_rptr)
	);
	// Trace: design.sv:28103:3
	assign src_ready_o = s_src_ready & !s_src_isolate_req;
	// Trace: design.sv:28105:3
	cdc_fifo_gray_dst_clearable_7A26D_20958 #(
		.T_WIDTH(WIDTH),
		.LOG_DEPTH(LOG_DEPTH),
		.SYNC_STAGES(SYNC_STAGES)
	) i_dst(
		.dst_rst_ni(dst_rst_ni),
		.dst_clk_i(dst_clk_i),
		.dst_clear_i(s_dst_clear_req),
		.dst_data_o(dst_data_o),
		.dst_valid_o(s_dst_valid),
		.dst_ready_i(dst_ready_i & !s_dst_isolate_req),
		.async_data_i(async_data),
		.async_wptr_i(async_wptr),
		.async_rptr_o(async_rptr)
	);
	// Trace: design.sv:28122:3
	assign dst_valid_o = s_dst_valid & !s_dst_isolate_req;
	// Trace: design.sv:28126:3
	cdc_reset_ctrlr #(.SYNC_STAGES(SYNC_STAGES - 1)) i_cdc_reset_ctrlr(
		.a_clk_i(src_clk_i),
		.a_rst_ni(src_rst_ni),
		.a_clear_i(src_clear_i),
		.a_clear_o(s_src_clear_req),
		.a_clear_ack_i(s_src_clear_ack_q),
		.a_isolate_o(s_src_isolate_req),
		.a_isolate_ack_i(s_src_isolate_ack_q),
		.b_clk_i(dst_clk_i),
		.b_rst_ni(dst_rst_ni),
		.b_clear_i(dst_clear_i),
		.b_clear_o(s_dst_clear_req),
		.b_clear_ack_i(s_dst_clear_ack_q),
		.b_isolate_o(s_dst_isolate_req),
		.b_isolate_ack_i(s_dst_isolate_ack_q)
	);
	// Trace: design.sv:28147:3
	always @(posedge src_clk_i or negedge src_rst_ni)
		// Trace: design.sv:28148:5
		if (!src_rst_ni) begin
			// Trace: design.sv:28149:7
			s_src_isolate_ack_q <= 1'b0;
			// Trace: design.sv:28150:7
			s_src_clear_ack_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:28152:7
			s_src_isolate_ack_q <= s_src_isolate_req;
			// Trace: design.sv:28153:7
			s_src_clear_ack_q <= s_src_clear_req;
		end
	// Trace: design.sv:28157:3
	always @(posedge dst_clk_i or negedge dst_rst_ni)
		// Trace: design.sv:28158:5
		if (!dst_rst_ni) begin
			// Trace: design.sv:28159:7
			s_dst_isolate_ack_q <= 1'b0;
			// Trace: design.sv:28160:7
			s_dst_clear_ack_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:28162:7
			s_dst_isolate_ack_q <= s_dst_isolate_req;
			// Trace: design.sv:28163:7
			s_dst_clear_ack_q <= s_dst_clear_req;
		end
	// Trace: design.sv:28168:3
	assign src_clear_pending_o = s_src_isolate_req;
	// Trace: design.sv:28171:3
	assign dst_clear_pending_o = s_dst_isolate_req;
endmodule
module cdc_fifo_gray_src_clearable_0070C_CFA0B (
	src_rst_ni,
	src_clk_i,
	src_clear_i,
	src_data_i,
	src_valid_i,
	src_ready_o,
	async_data_o,
	async_wptr_o,
	async_rptr_i
);
	// removed localparam type T_WIDTH_type
	parameter [31:0] T_WIDTH = 0;
	// Trace: design.sv:28187:18
	// removed localparam type T
	// Trace: design.sv:28188:13
	parameter signed [31:0] LOG_DEPTH = 3;
	// Trace: design.sv:28189:13
	parameter signed [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:28191:3
	input wire src_rst_ni;
	// Trace: design.sv:28192:3
	input wire src_clk_i;
	// Trace: design.sv:28193:3
	input wire src_clear_i;
	// Trace: design.sv:28194:3
	input wire [T_WIDTH - 1:0] src_data_i;
	// Trace: design.sv:28195:3
	input wire src_valid_i;
	// Trace: design.sv:28196:3
	output wire src_ready_o;
	// Trace: design.sv:28198:3
	output wire [((2 ** LOG_DEPTH) * T_WIDTH) - 1:0] async_data_o;
	// Trace: design.sv:28199:3
	output wire [LOG_DEPTH:0] async_wptr_o;
	// Trace: design.sv:28200:3
	input wire [LOG_DEPTH:0] async_rptr_i;
	// Trace: design.sv:28203:3
	localparam signed [31:0] PtrWidth = LOG_DEPTH + 1;
	// Trace: design.sv:28204:3
	localparam [PtrWidth - 1:0] PtrFull = 1 << LOG_DEPTH;
	// Trace: design.sv:28206:3
	reg [((2 ** LOG_DEPTH) * T_WIDTH) - 1:0] data_q;
	// Trace: design.sv:28207:3
	reg [PtrWidth - 1:0] wptr_q;
	wire [PtrWidth - 1:0] wptr_d;
	wire [PtrWidth - 1:0] wptr_bin;
	wire [PtrWidth - 1:0] wptr_next;
	wire [PtrWidth - 1:0] rptr;
	wire [PtrWidth - 1:0] rptr_bin;
	// Trace: design.sv:28210:3
	assign async_data_o = data_q;
	// Trace: design.sv:28211:3
	genvar _gv_i_28;
	generate
		for (_gv_i_28 = 0; _gv_i_28 < (2 ** LOG_DEPTH); _gv_i_28 = _gv_i_28 + 1) begin : gen_word
			localparam i = _gv_i_28;
			// Trace: macro expansion of FFLNR at design.sv:28213:78
			always @(posedge src_clk_i)
				// Trace: macro expansion of FFLNR at design.sv:28213:120
				if ((src_valid_i & src_ready_o) & (wptr_bin[LOG_DEPTH - 1:0] == i))
					// Trace: macro expansion of FFLNR at design.sv:28213:162
					data_q[i * T_WIDTH+:T_WIDTH] <= src_data_i;
		end
	endgenerate
	// Trace: design.sv:28217:3
	genvar _gv_i_29;
	generate
		for (_gv_i_29 = 0; _gv_i_29 < PtrWidth; _gv_i_29 = _gv_i_29 + 1) begin : gen_sync
			localparam i = _gv_i_29;
			// Trace: design.sv:28218:5
			sync #(.STAGES(SYNC_STAGES)) i_sync(
				.clk_i(src_clk_i),
				.rst_ni(src_rst_ni),
				.serial_i(async_rptr_i[i]),
				.serial_o(rptr[i])
			);
		end
	endgenerate
	// Trace: design.sv:28225:3
	gray_to_binary #(.N(PtrWidth)) i_rptr_g2b(
		.A(rptr),
		.Z(rptr_bin)
	);
	// Trace: design.sv:28228:3
	assign wptr_next = wptr_bin + 1;
	// Trace: design.sv:28229:3
	gray_to_binary #(.N(PtrWidth)) i_wptr_g2b(
		.A(wptr_q),
		.Z(wptr_bin)
	);
	// Trace: design.sv:28230:3
	binary_to_gray #(.N(PtrWidth)) i_wptr_b2g(
		.A(wptr_next),
		.Z(wptr_d)
	);
	// Trace: macro expansion of FFLARNC at design.sv:28231:317
	always @(posedge src_clk_i or negedge src_rst_ni)
		// Trace: macro expansion of FFLARNC at design.sv:28231:395
		if (!src_rst_ni)
			// Trace: macro expansion of FFLARNC at design.sv:28231:473
			wptr_q <= 1'sb0;
		else
			// Trace: macro expansion of FFLARNC at design.sv:28231:625
			if (src_clear_i)
				// Trace: macro expansion of FFLARNC at design.sv:28231:703
				wptr_q <= 1'sb0;
			else if (src_valid_i & src_ready_o)
				// Trace: macro expansion of FFLARNC at design.sv:28231:855
				wptr_q <= wptr_d;
	// Trace: design.sv:28232:3
	assign async_wptr_o = wptr_q;
	// Trace: design.sv:28238:3
	assign src_ready_o = (wptr_bin ^ rptr_bin) != PtrFull;
endmodule
module cdc_fifo_gray_dst_clearable_7A26D_20958 (
	dst_rst_ni,
	dst_clk_i,
	dst_clear_i,
	dst_data_o,
	dst_valid_o,
	dst_ready_i,
	async_data_i,
	async_wptr_i,
	async_rptr_o
);
	// removed localparam type T_WIDTH_type
	parameter [31:0] T_WIDTH = 0;
	// Trace: design.sv:28246:18
	// removed localparam type T
	// Trace: design.sv:28247:13
	parameter signed [31:0] LOG_DEPTH = 3;
	// Trace: design.sv:28248:13
	parameter signed [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:28250:3
	input wire dst_rst_ni;
	// Trace: design.sv:28251:3
	input wire dst_clk_i;
	// Trace: design.sv:28252:3
	input wire dst_clear_i;
	// Trace: design.sv:28253:3
	output wire [T_WIDTH - 1:0] dst_data_o;
	// Trace: design.sv:28254:3
	output wire dst_valid_o;
	// Trace: design.sv:28255:3
	input wire dst_ready_i;
	// Trace: design.sv:28257:3
	input wire [((2 ** LOG_DEPTH) * T_WIDTH) - 1:0] async_data_i;
	// Trace: design.sv:28258:3
	input wire [LOG_DEPTH:0] async_wptr_i;
	// Trace: design.sv:28259:3
	output wire [LOG_DEPTH:0] async_rptr_o;
	// Trace: design.sv:28262:3
	localparam signed [31:0] PtrWidth = LOG_DEPTH + 1;
	// Trace: design.sv:28263:3
	localparam [PtrWidth - 1:0] PtrEmpty = 1'sb0;
	// Trace: design.sv:28265:3
	wire [T_WIDTH - 1:0] dst_data;
	// Trace: design.sv:28266:3
	reg [PtrWidth - 1:0] rptr_q;
	wire [PtrWidth - 1:0] rptr_d;
	wire [PtrWidth - 1:0] rptr_bin;
	wire [PtrWidth - 1:0] rptr_next;
	wire [PtrWidth - 1:0] wptr;
	wire [PtrWidth - 1:0] wptr_bin;
	// Trace: design.sv:28267:3
	wire dst_valid;
	wire dst_ready;
	// Trace: design.sv:28269:3
	assign dst_data = async_data_i[rptr_bin[LOG_DEPTH - 1:0] * T_WIDTH+:T_WIDTH];
	// Trace: design.sv:28272:3
	assign rptr_next = rptr_bin + 1;
	// Trace: design.sv:28273:3
	gray_to_binary #(.N(PtrWidth)) i_rptr_g2b(
		.A(rptr_q),
		.Z(rptr_bin)
	);
	// Trace: design.sv:28274:3
	binary_to_gray #(.N(PtrWidth)) i_rptr_b2g(
		.A(rptr_next),
		.Z(rptr_d)
	);
	// Trace: macro expansion of FFLARNC at design.sv:28275:313
	always @(posedge dst_clk_i or negedge dst_rst_ni)
		// Trace: macro expansion of FFLARNC at design.sv:28275:391
		if (!dst_rst_ni)
			// Trace: macro expansion of FFLARNC at design.sv:28275:469
			rptr_q <= 1'sb0;
		else
			// Trace: macro expansion of FFLARNC at design.sv:28275:621
			if (dst_clear_i)
				// Trace: macro expansion of FFLARNC at design.sv:28275:699
				rptr_q <= 1'sb0;
			else if (dst_valid & dst_ready)
				// Trace: macro expansion of FFLARNC at design.sv:28275:851
				rptr_q <= rptr_d;
	// Trace: design.sv:28276:3
	assign async_rptr_o = rptr_q;
	// Trace: design.sv:28279:3
	genvar _gv_i_30;
	generate
		for (_gv_i_30 = 0; _gv_i_30 < PtrWidth; _gv_i_30 = _gv_i_30 + 1) begin : gen_sync
			localparam i = _gv_i_30;
			// Trace: design.sv:28280:5
			sync #(.STAGES(SYNC_STAGES)) i_sync(
				.clk_i(dst_clk_i),
				.rst_ni(dst_rst_ni),
				.serial_i(async_wptr_i[i]),
				.serial_o(wptr[i])
			);
		end
	endgenerate
	// Trace: design.sv:28287:3
	gray_to_binary #(.N(PtrWidth)) i_wptr_g2b(
		.A(wptr),
		.Z(wptr_bin)
	);
	// Trace: design.sv:28293:3
	assign dst_valid = (wptr_bin ^ rptr_bin) != PtrEmpty;
	// Trace: design.sv:28296:3
	spill_register_flushable_44288_566E2 #(.T_T_WIDTH(T_WIDTH)) i_spill_register(
		.clk_i(dst_clk_i),
		.rst_ni(dst_rst_ni),
		.flush_i(dst_clear_i),
		.valid_i(dst_valid & !dst_clear_i),
		.ready_o(dst_ready),
		.data_i(dst_data),
		.valid_o(dst_valid_o),
		.ready_i(dst_ready_i),
		.data_o(dst_data_o)
	);
endmodule
module cdc_2phase_clearable_88D17 (
	src_rst_ni,
	src_clk_i,
	src_clear_i,
	src_clear_pending_o,
	src_data_i,
	src_valid_i,
	src_ready_o,
	dst_rst_ni,
	dst_clk_i,
	dst_clear_i,
	dst_clear_pending_o,
	dst_data_o,
	dst_valid_o,
	dst_ready_i
);
	// Trace: design.sv:28364:18
	// removed localparam type T
	// Trace: design.sv:28365:13
	parameter [31:0] SYNC_STAGES = 3;
	// Trace: design.sv:28366:13
	parameter signed [31:0] CLEAR_ON_ASYNC_RESET = 1;
	// Trace: design.sv:28368:3
	input wire src_rst_ni;
	// Trace: design.sv:28369:3
	input wire src_clk_i;
	// Trace: design.sv:28370:3
	input wire src_clear_i;
	// Trace: design.sv:28371:3
	output wire src_clear_pending_o;
	// Trace: design.sv:28372:3
	input wire [40:0] src_data_i;
	// Trace: design.sv:28373:3
	input wire src_valid_i;
	// Trace: design.sv:28374:3
	output wire src_ready_o;
	// Trace: design.sv:28376:3
	input wire dst_rst_ni;
	// Trace: design.sv:28377:3
	input wire dst_clk_i;
	// Trace: design.sv:28378:3
	input wire dst_clear_i;
	// Trace: design.sv:28379:3
	output wire dst_clear_pending_o;
	// Trace: design.sv:28380:3
	output wire [40:0] dst_data_o;
	// Trace: design.sv:28381:3
	output wire dst_valid_o;
	// Trace: design.sv:28382:3
	input wire dst_ready_i;
	// Trace: design.sv:28384:3
	wire s_src_clear_req;
	// Trace: design.sv:28385:3
	reg s_src_clear_ack_q;
	// Trace: design.sv:28386:3
	wire s_src_ready;
	// Trace: design.sv:28387:3
	wire s_src_isolate_req;
	// Trace: design.sv:28388:3
	reg s_src_isolate_ack_q;
	// Trace: design.sv:28389:3
	wire s_dst_clear_req;
	// Trace: design.sv:28390:3
	reg s_dst_clear_ack_q;
	// Trace: design.sv:28391:3
	wire s_dst_valid;
	// Trace: design.sv:28392:3
	wire s_dst_isolate_req;
	// Trace: design.sv:28393:3
	reg s_dst_isolate_ack_q;
	// Trace: design.sv:28396:4
	wire async_req;
	// Trace: design.sv:28397:4
	wire async_ack;
	// Trace: design.sv:28398:4
	wire [40:0] async_data;
	// Trace: design.sv:28400:3
	generate
		if (CLEAR_ON_ASYNC_RESET) begin : gen_elaboration_assertion
			if (SYNC_STAGES < 3) begin : genblk1
				// Trace: design.sv:28402:7
				$error("The clearable 2-phase CDC with async reset", "synchronization requires at least 3 synchronizer stages for the FIFO.");
			end
		end
		else begin : gen_elaboration_assertion
			if (SYNC_STAGES < 2) begin : gen_elaboration_assertion
				// Trace: design.sv:28406:7
				$error("A minimum of 2 synchronizer stages is required for proper functionality.");
			end
		end
	endgenerate
	// Trace: design.sv:28412:3
	cdc_2phase_src_clearable_A5DBE #(.SYNC_STAGES(SYNC_STAGES)) i_src(
		.rst_ni(src_rst_ni),
		.clk_i(src_clk_i),
		.clear_i(s_src_clear_req),
		.data_i(src_data_i),
		.valid_i(src_valid_i & !s_src_isolate_req),
		.ready_o(s_src_ready),
		.async_req_o(async_req),
		.async_ack_i(async_ack),
		.async_data_o(async_data)
	);
	// Trace: design.sv:28427:3
	assign src_ready_o = s_src_ready & !s_src_isolate_req;
	// Trace: design.sv:28431:3
	cdc_2phase_dst_clearable_3F52F #(.SYNC_STAGES(SYNC_STAGES)) i_dst(
		.rst_ni(dst_rst_ni),
		.clk_i(dst_clk_i),
		.clear_i(s_dst_clear_req),
		.data_o(dst_data_o),
		.valid_o(s_dst_valid),
		.ready_i(dst_ready_i & !s_dst_isolate_req),
		.async_req_i(async_req),
		.async_ack_o(async_ack),
		.async_data_i(async_data)
	);
	// Trace: design.sv:28446:3
	assign dst_valid_o = s_dst_valid & !s_dst_isolate_req;
	// Trace: design.sv:28450:3
	cdc_reset_ctrlr #(.SYNC_STAGES(SYNC_STAGES - 1)) i_cdc_reset_ctrlr(
		.a_clk_i(src_clk_i),
		.a_rst_ni(src_rst_ni),
		.a_clear_i(src_clear_i),
		.a_clear_o(s_src_clear_req),
		.a_clear_ack_i(s_src_clear_ack_q),
		.a_isolate_o(s_src_isolate_req),
		.a_isolate_ack_i(s_src_isolate_ack_q),
		.b_clk_i(dst_clk_i),
		.b_rst_ni(dst_rst_ni),
		.b_clear_i(dst_clear_i),
		.b_clear_o(s_dst_clear_req),
		.b_clear_ack_i(s_dst_clear_ack_q),
		.b_isolate_o(s_dst_isolate_req),
		.b_isolate_ack_i(s_dst_isolate_ack_q)
	);
	// Trace: design.sv:28471:3
	always @(posedge src_clk_i or negedge src_rst_ni)
		// Trace: design.sv:28472:5
		if (!src_rst_ni) begin
			// Trace: design.sv:28473:7
			s_src_isolate_ack_q <= 1'b0;
			// Trace: design.sv:28474:7
			s_src_clear_ack_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:28476:7
			s_src_isolate_ack_q <= s_src_isolate_req;
			// Trace: design.sv:28477:7
			s_src_clear_ack_q <= s_src_clear_req;
		end
	// Trace: design.sv:28481:3
	always @(posedge dst_clk_i or negedge dst_rst_ni)
		// Trace: design.sv:28482:5
		if (!dst_rst_ni) begin
			// Trace: design.sv:28483:7
			s_dst_isolate_ack_q <= 1'b0;
			// Trace: design.sv:28484:7
			s_dst_clear_ack_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:28486:7
			s_dst_isolate_ack_q <= s_dst_isolate_req;
			// Trace: design.sv:28487:7
			s_dst_clear_ack_q <= s_dst_clear_req;
		end
	// Trace: design.sv:28492:3
	assign src_clear_pending_o = s_src_isolate_req;
	// Trace: design.sv:28495:3
	assign dst_clear_pending_o = s_dst_isolate_req;
endmodule
module cdc_2phase_clearable_DC602 (
	src_rst_ni,
	src_clk_i,
	src_clear_i,
	src_clear_pending_o,
	src_data_i,
	src_valid_i,
	src_ready_o,
	dst_rst_ni,
	dst_clk_i,
	dst_clear_i,
	dst_clear_pending_o,
	dst_data_o,
	dst_valid_o,
	dst_ready_i
);
	// Trace: design.sv:28364:18
	// removed localparam type T
	// Trace: design.sv:28365:13
	parameter [31:0] SYNC_STAGES = 3;
	// Trace: design.sv:28366:13
	parameter signed [31:0] CLEAR_ON_ASYNC_RESET = 1;
	// Trace: design.sv:28368:3
	input wire src_rst_ni;
	// Trace: design.sv:28369:3
	input wire src_clk_i;
	// Trace: design.sv:28370:3
	input wire src_clear_i;
	// Trace: design.sv:28371:3
	output wire src_clear_pending_o;
	// Trace: design.sv:28372:3
	input wire [33:0] src_data_i;
	// Trace: design.sv:28373:3
	input wire src_valid_i;
	// Trace: design.sv:28374:3
	output wire src_ready_o;
	// Trace: design.sv:28376:3
	input wire dst_rst_ni;
	// Trace: design.sv:28377:3
	input wire dst_clk_i;
	// Trace: design.sv:28378:3
	input wire dst_clear_i;
	// Trace: design.sv:28379:3
	output wire dst_clear_pending_o;
	// Trace: design.sv:28380:3
	output wire [33:0] dst_data_o;
	// Trace: design.sv:28381:3
	output wire dst_valid_o;
	// Trace: design.sv:28382:3
	input wire dst_ready_i;
	// Trace: design.sv:28384:3
	wire s_src_clear_req;
	// Trace: design.sv:28385:3
	reg s_src_clear_ack_q;
	// Trace: design.sv:28386:3
	wire s_src_ready;
	// Trace: design.sv:28387:3
	wire s_src_isolate_req;
	// Trace: design.sv:28388:3
	reg s_src_isolate_ack_q;
	// Trace: design.sv:28389:3
	wire s_dst_clear_req;
	// Trace: design.sv:28390:3
	reg s_dst_clear_ack_q;
	// Trace: design.sv:28391:3
	wire s_dst_valid;
	// Trace: design.sv:28392:3
	wire s_dst_isolate_req;
	// Trace: design.sv:28393:3
	reg s_dst_isolate_ack_q;
	// Trace: design.sv:28396:4
	wire async_req;
	// Trace: design.sv:28397:4
	wire async_ack;
	// Trace: design.sv:28398:4
	wire [33:0] async_data;
	// Trace: design.sv:28400:3
	generate
		if (CLEAR_ON_ASYNC_RESET) begin : gen_elaboration_assertion
			if (SYNC_STAGES < 3) begin : genblk1
				// Trace: design.sv:28402:7
				$error("The clearable 2-phase CDC with async reset", "synchronization requires at least 3 synchronizer stages for the FIFO.");
			end
		end
		else begin : gen_elaboration_assertion
			if (SYNC_STAGES < 2) begin : gen_elaboration_assertion
				// Trace: design.sv:28406:7
				$error("A minimum of 2 synchronizer stages is required for proper functionality.");
			end
		end
	endgenerate
	// Trace: design.sv:28412:3
	cdc_2phase_src_clearable_B85FB #(.SYNC_STAGES(SYNC_STAGES)) i_src(
		.rst_ni(src_rst_ni),
		.clk_i(src_clk_i),
		.clear_i(s_src_clear_req),
		.data_i(src_data_i),
		.valid_i(src_valid_i & !s_src_isolate_req),
		.ready_o(s_src_ready),
		.async_req_o(async_req),
		.async_ack_i(async_ack),
		.async_data_o(async_data)
	);
	// Trace: design.sv:28427:3
	assign src_ready_o = s_src_ready & !s_src_isolate_req;
	// Trace: design.sv:28431:3
	cdc_2phase_dst_clearable_0389A #(.SYNC_STAGES(SYNC_STAGES)) i_dst(
		.rst_ni(dst_rst_ni),
		.clk_i(dst_clk_i),
		.clear_i(s_dst_clear_req),
		.data_o(dst_data_o),
		.valid_o(s_dst_valid),
		.ready_i(dst_ready_i & !s_dst_isolate_req),
		.async_req_i(async_req),
		.async_ack_o(async_ack),
		.async_data_i(async_data)
	);
	// Trace: design.sv:28446:3
	assign dst_valid_o = s_dst_valid & !s_dst_isolate_req;
	// Trace: design.sv:28450:3
	cdc_reset_ctrlr #(.SYNC_STAGES(SYNC_STAGES - 1)) i_cdc_reset_ctrlr(
		.a_clk_i(src_clk_i),
		.a_rst_ni(src_rst_ni),
		.a_clear_i(src_clear_i),
		.a_clear_o(s_src_clear_req),
		.a_clear_ack_i(s_src_clear_ack_q),
		.a_isolate_o(s_src_isolate_req),
		.a_isolate_ack_i(s_src_isolate_ack_q),
		.b_clk_i(dst_clk_i),
		.b_rst_ni(dst_rst_ni),
		.b_clear_i(dst_clear_i),
		.b_clear_o(s_dst_clear_req),
		.b_clear_ack_i(s_dst_clear_ack_q),
		.b_isolate_o(s_dst_isolate_req),
		.b_isolate_ack_i(s_dst_isolate_ack_q)
	);
	// Trace: design.sv:28471:3
	always @(posedge src_clk_i or negedge src_rst_ni)
		// Trace: design.sv:28472:5
		if (!src_rst_ni) begin
			// Trace: design.sv:28473:7
			s_src_isolate_ack_q <= 1'b0;
			// Trace: design.sv:28474:7
			s_src_clear_ack_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:28476:7
			s_src_isolate_ack_q <= s_src_isolate_req;
			// Trace: design.sv:28477:7
			s_src_clear_ack_q <= s_src_clear_req;
		end
	// Trace: design.sv:28481:3
	always @(posedge dst_clk_i or negedge dst_rst_ni)
		// Trace: design.sv:28482:5
		if (!dst_rst_ni) begin
			// Trace: design.sv:28483:7
			s_dst_isolate_ack_q <= 1'b0;
			// Trace: design.sv:28484:7
			s_dst_clear_ack_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:28486:7
			s_dst_isolate_ack_q <= s_dst_isolate_req;
			// Trace: design.sv:28487:7
			s_dst_clear_ack_q <= s_dst_clear_req;
		end
	// Trace: design.sv:28492:3
	assign src_clear_pending_o = s_src_isolate_req;
	// Trace: design.sv:28495:3
	assign dst_clear_pending_o = s_dst_isolate_req;
endmodule
module cdc_2phase_src_clearable_A5DBE (
	rst_ni,
	clk_i,
	clear_i,
	data_i,
	valid_i,
	ready_o,
	async_req_o,
	async_ack_i,
	async_data_o
);
	reg _sv2v_0;
	// Trace: design.sv:28511:18
	// removed localparam type T
	// Trace: design.sv:28512:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:28514:3
	input wire rst_ni;
	// Trace: design.sv:28515:3
	input wire clk_i;
	// Trace: design.sv:28516:3
	input wire clear_i;
	// Trace: design.sv:28517:3
	input wire [40:0] data_i;
	// Trace: design.sv:28518:3
	input wire valid_i;
	// Trace: design.sv:28519:3
	output wire ready_o;
	// Trace: design.sv:28520:3
	output wire async_req_o;
	// Trace: design.sv:28521:3
	input wire async_ack_i;
	// Trace: design.sv:28522:3
	output wire [40:0] async_data_o;
	// Trace: design.sv:28526:3
	reg req_src_d;
	reg req_src_q;
	wire ack_synced;
	// Trace: design.sv:28528:3
	reg [40:0] data_src_d;
	reg [40:0] data_src_q;
	// Trace: design.sv:28531:3
	sync #(.STAGES(SYNC_STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(async_ack_i),
		.serial_o(ack_synced)
	);
	// Trace: design.sv:28542:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:28543:5
		data_src_d = data_src_q;
		// Trace: design.sv:28544:5
		req_src_d = req_src_q;
		// Trace: design.sv:28545:5
		if (clear_i)
			// Trace: design.sv:28546:7
			req_src_d = 1'b0;
		else if (valid_i && ready_o) begin
			// Trace: design.sv:28549:7
			req_src_d = ~req_src_q;
			// Trace: design.sv:28550:7
			data_src_d = data_i;
		end
	end
	// Trace: macro expansion of FFNR at design.sv:28554:37
	always @(posedge clk_i)
		// Trace: macro expansion of FFNR at design.sv:28554:77
		data_src_q <= data_src_d;
	// Trace: design.sv:28556:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:28557:5
		if (!rst_ni)
			// Trace: design.sv:28558:7
			req_src_q <= 0;
		else
			// Trace: design.sv:28560:7
			req_src_q <= req_src_d;
	// Trace: design.sv:28565:3
	assign ready_o = req_src_q == ack_synced;
	// Trace: design.sv:28566:3
	assign async_req_o = req_src_q;
	// Trace: design.sv:28567:3
	assign async_data_o = data_src_q;
	initial _sv2v_0 = 0;
endmodule
module cdc_2phase_src_clearable_B85FB (
	rst_ni,
	clk_i,
	clear_i,
	data_i,
	valid_i,
	ready_o,
	async_req_o,
	async_ack_i,
	async_data_o
);
	reg _sv2v_0;
	// Trace: design.sv:28511:18
	// removed localparam type T
	// Trace: design.sv:28512:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:28514:3
	input wire rst_ni;
	// Trace: design.sv:28515:3
	input wire clk_i;
	// Trace: design.sv:28516:3
	input wire clear_i;
	// Trace: design.sv:28517:3
	input wire [33:0] data_i;
	// Trace: design.sv:28518:3
	input wire valid_i;
	// Trace: design.sv:28519:3
	output wire ready_o;
	// Trace: design.sv:28520:3
	output wire async_req_o;
	// Trace: design.sv:28521:3
	input wire async_ack_i;
	// Trace: design.sv:28522:3
	output wire [33:0] async_data_o;
	// Trace: design.sv:28526:3
	reg req_src_d;
	reg req_src_q;
	wire ack_synced;
	// Trace: design.sv:28528:3
	reg [33:0] data_src_d;
	reg [33:0] data_src_q;
	// Trace: design.sv:28531:3
	sync #(.STAGES(SYNC_STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(async_ack_i),
		.serial_o(ack_synced)
	);
	// Trace: design.sv:28542:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:28543:5
		data_src_d = data_src_q;
		// Trace: design.sv:28544:5
		req_src_d = req_src_q;
		// Trace: design.sv:28545:5
		if (clear_i)
			// Trace: design.sv:28546:7
			req_src_d = 1'b0;
		else if (valid_i && ready_o) begin
			// Trace: design.sv:28549:7
			req_src_d = ~req_src_q;
			// Trace: design.sv:28550:7
			data_src_d = data_i;
		end
	end
	// Trace: macro expansion of FFNR at design.sv:28554:37
	always @(posedge clk_i)
		// Trace: macro expansion of FFNR at design.sv:28554:77
		data_src_q <= data_src_d;
	// Trace: design.sv:28556:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:28557:5
		if (!rst_ni)
			// Trace: design.sv:28558:7
			req_src_q <= 0;
		else
			// Trace: design.sv:28560:7
			req_src_q <= req_src_d;
	// Trace: design.sv:28565:3
	assign ready_o = req_src_q == ack_synced;
	// Trace: design.sv:28566:3
	assign async_req_o = req_src_q;
	// Trace: design.sv:28567:3
	assign async_data_o = data_src_q;
	initial _sv2v_0 = 0;
endmodule
module cdc_2phase_dst_clearable_0389A (
	rst_ni,
	clk_i,
	clear_i,
	data_o,
	valid_o,
	ready_i,
	async_req_i,
	async_ack_o,
	async_data_i
);
	reg _sv2v_0;
	// Trace: design.sv:28585:18
	// removed localparam type T
	// Trace: design.sv:28586:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:28588:3
	input wire rst_ni;
	// Trace: design.sv:28589:3
	input wire clk_i;
	// Trace: design.sv:28590:3
	input wire clear_i;
	// Trace: design.sv:28591:3
	output wire [33:0] data_o;
	// Trace: design.sv:28592:3
	output wire valid_o;
	// Trace: design.sv:28593:3
	input wire ready_i;
	// Trace: design.sv:28594:3
	input wire async_req_i;
	// Trace: design.sv:28595:3
	output wire async_ack_o;
	// Trace: design.sv:28596:3
	input wire [33:0] async_data_i;
	// Trace: design.sv:28601:2
	reg ack_dst_d;
	reg ack_dst_q;
	wire req_synced;
	reg req_synced_q1;
	// Trace: design.sv:28603:3
	reg [33:0] data_dst_d;
	reg [33:0] data_dst_q;
	// Trace: design.sv:28607:3
	sync #(.STAGES(SYNC_STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(async_req_i),
		.serial_o(req_synced)
	);
	// Trace: design.sv:28617:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:28618:5
		ack_dst_d = ack_dst_q;
		// Trace: design.sv:28619:5
		if (clear_i)
			// Trace: design.sv:28620:7
			ack_dst_d = 1'b0;
		else if (valid_o && ready_i)
			// Trace: design.sv:28622:7
			ack_dst_d = ~ack_dst_q;
	end
	// Trace: design.sv:28628:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:28629:5
		data_dst_d = data_dst_q;
		// Trace: design.sv:28630:5
		if ((req_synced != req_synced_q1) && !valid_o)
			// Trace: design.sv:28631:7
			data_dst_d = async_data_i;
	end
	// Trace: macro expansion of FFNR at design.sv:28635:37
	always @(posedge clk_i)
		// Trace: macro expansion of FFNR at design.sv:28635:77
		data_dst_q <= data_dst_d;
	// Trace: design.sv:28637:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:28638:5
		if (!rst_ni) begin
			// Trace: design.sv:28639:7
			ack_dst_q <= 0;
			// Trace: design.sv:28640:7
			req_synced_q1 <= 1'b0;
		end
		else begin
			// Trace: design.sv:28642:7
			ack_dst_q <= ack_dst_d;
			// Trace: design.sv:28645:7
			req_synced_q1 <= req_synced;
		end
	// Trace: design.sv:28650:3
	assign valid_o = ack_dst_q != req_synced_q1;
	// Trace: design.sv:28651:3
	assign data_o = data_dst_q;
	// Trace: design.sv:28652:3
	assign async_ack_o = ack_dst_q;
	initial _sv2v_0 = 0;
endmodule
module cdc_2phase_dst_clearable_3F52F (
	rst_ni,
	clk_i,
	clear_i,
	data_o,
	valid_o,
	ready_i,
	async_req_i,
	async_ack_o,
	async_data_i
);
	reg _sv2v_0;
	// Trace: design.sv:28585:18
	// removed localparam type T
	// Trace: design.sv:28586:13
	parameter [31:0] SYNC_STAGES = 2;
	// Trace: design.sv:28588:3
	input wire rst_ni;
	// Trace: design.sv:28589:3
	input wire clk_i;
	// Trace: design.sv:28590:3
	input wire clear_i;
	// Trace: design.sv:28591:3
	output wire [40:0] data_o;
	// Trace: design.sv:28592:3
	output wire valid_o;
	// Trace: design.sv:28593:3
	input wire ready_i;
	// Trace: design.sv:28594:3
	input wire async_req_i;
	// Trace: design.sv:28595:3
	output wire async_ack_o;
	// Trace: design.sv:28596:3
	input wire [40:0] async_data_i;
	// Trace: design.sv:28601:2
	reg ack_dst_d;
	reg ack_dst_q;
	wire req_synced;
	reg req_synced_q1;
	// Trace: design.sv:28603:3
	reg [40:0] data_dst_d;
	reg [40:0] data_dst_q;
	// Trace: design.sv:28607:3
	sync #(.STAGES(SYNC_STAGES)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(async_req_i),
		.serial_o(req_synced)
	);
	// Trace: design.sv:28617:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:28618:5
		ack_dst_d = ack_dst_q;
		// Trace: design.sv:28619:5
		if (clear_i)
			// Trace: design.sv:28620:7
			ack_dst_d = 1'b0;
		else if (valid_o && ready_i)
			// Trace: design.sv:28622:7
			ack_dst_d = ~ack_dst_q;
	end
	// Trace: design.sv:28628:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:28629:5
		data_dst_d = data_dst_q;
		// Trace: design.sv:28630:5
		if ((req_synced != req_synced_q1) && !valid_o)
			// Trace: design.sv:28631:7
			data_dst_d = async_data_i;
	end
	// Trace: macro expansion of FFNR at design.sv:28635:37
	always @(posedge clk_i)
		// Trace: macro expansion of FFNR at design.sv:28635:77
		data_dst_q <= data_dst_d;
	// Trace: design.sv:28637:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:28638:5
		if (!rst_ni) begin
			// Trace: design.sv:28639:7
			ack_dst_q <= 0;
			// Trace: design.sv:28640:7
			req_synced_q1 <= 1'b0;
		end
		else begin
			// Trace: design.sv:28642:7
			ack_dst_q <= ack_dst_d;
			// Trace: design.sv:28645:7
			req_synced_q1 <= req_synced;
		end
	// Trace: design.sv:28650:3
	assign valid_o = ack_dst_q != req_synced_q1;
	// Trace: design.sv:28651:3
	assign data_o = data_dst_q;
	// Trace: design.sv:28652:3
	assign async_ack_o = ack_dst_q;
	initial _sv2v_0 = 0;
endmodule
module mem_to_banks (
	clk_i,
	rst_ni,
	req_i,
	gnt_o,
	addr_i,
	wdata_i,
	strb_i,
	atop_i,
	we_i,
	rvalid_o,
	rdata_o,
	bank_req_o,
	bank_gnt_i,
	bank_addr_o,
	bank_wdata_o,
	bank_strb_o,
	bank_atop_o,
	bank_we_o,
	bank_rvalid_i,
	bank_rdata_i
);
	// Trace: design.sv:28672:13
	parameter [31:0] AddrWidth = 32'd0;
	// Trace: design.sv:28674:13
	parameter [31:0] DataWidth = 32'd0;
	// Trace: design.sv:28676:13
	parameter [31:0] AtopWidth = 32'd0;
	// Trace: design.sv:28678:13
	parameter [31:0] NumBanks = 32'd0;
	// Trace: design.sv:28680:13
	parameter [0:0] HideStrb = 1'b0;
	// Trace: design.sv:28682:13
	parameter [31:0] MaxTrans = 32'd1;
	// Trace: design.sv:28684:13
	parameter [31:0] FifoDepth = 32'd1;
	// Trace: design.sv:28686:19
	// removed localparam type atop_t
	// Trace: design.sv:28688:19
	// removed localparam type addr_t
	// Trace: design.sv:28690:19
	// removed localparam type inp_data_t
	// Trace: design.sv:28692:19
	// removed localparam type inp_strb_t
	// Trace: design.sv:28694:19
	// removed localparam type oup_data_t
	// Trace: design.sv:28696:19
	// removed localparam type oup_strb_t
	// Trace: design.sv:28699:3
	input wire clk_i;
	// Trace: design.sv:28701:3
	input wire rst_ni;
	// Trace: design.sv:28703:3
	input wire req_i;
	// Trace: design.sv:28705:3
	output wire gnt_o;
	// Trace: design.sv:28707:3
	input wire [AddrWidth - 1:0] addr_i;
	// Trace: design.sv:28709:3
	input wire [DataWidth - 1:0] wdata_i;
	// Trace: design.sv:28711:3
	input wire [(DataWidth / 8) - 1:0] strb_i;
	// Trace: design.sv:28713:3
	input wire [AtopWidth - 1:0] atop_i;
	// Trace: design.sv:28715:3
	input wire we_i;
	// Trace: design.sv:28717:3
	output wire rvalid_o;
	// Trace: design.sv:28719:3
	output wire [DataWidth - 1:0] rdata_o;
	// Trace: design.sv:28721:3
	output wire [NumBanks - 1:0] bank_req_o;
	// Trace: design.sv:28723:3
	input wire [NumBanks - 1:0] bank_gnt_i;
	// Trace: design.sv:28725:3
	output wire [(NumBanks * AddrWidth) - 1:0] bank_addr_o;
	// Trace: design.sv:28727:3
	output wire [(NumBanks * (DataWidth / NumBanks)) - 1:0] bank_wdata_o;
	// Trace: design.sv:28729:3
	output wire [(NumBanks * ((DataWidth / NumBanks) / 8)) - 1:0] bank_strb_o;
	// Trace: design.sv:28731:3
	output wire [(NumBanks * AtopWidth) - 1:0] bank_atop_o;
	// Trace: design.sv:28733:3
	output wire [NumBanks - 1:0] bank_we_o;
	// Trace: design.sv:28735:3
	input wire [NumBanks - 1:0] bank_rvalid_i;
	// Trace: design.sv:28737:3
	input wire [(NumBanks * (DataWidth / NumBanks)) - 1:0] bank_rdata_i;
	// Trace: design.sv:28740:3
	localparam [31:0] DataBytes = DataWidth / 8;
	// Trace: design.sv:28741:3
	localparam [31:0] BitsPerBank = DataWidth / NumBanks;
	// Trace: design.sv:28742:3
	localparam [31:0] BytesPerBank = (DataWidth / NumBanks) / 8;
	// Trace: design.sv:28744:3
	// removed localparam type req_t
	// Trace: design.sv:28752:3
	wire req_valid;
	// Trace: design.sv:28753:3
	wire [NumBanks - 1:0] req_ready;
	wire [NumBanks - 1:0] resp_valid;
	wire [NumBanks - 1:0] resp_ready;
	// Trace: design.sv:28755:3
	wire [(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (NumBanks * ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1)) - 1 : (NumBanks * (1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) - 1)):(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? 0 : (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0)] bank_req;
	wire [(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (NumBanks * ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1)) - 1 : (NumBanks * (1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) - 1)):(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? 0 : (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0)] bank_oup;
	// Trace: design.sv:28757:3
	wire [NumBanks - 1:0] bank_req_internal;
	wire [NumBanks - 1:0] bank_gnt_internal;
	wire [NumBanks - 1:0] zero_strobe;
	wire [NumBanks - 1:0] dead_response;
	// Trace: design.sv:28758:3
	wire dead_write_fifo_full;
	// Trace: design.sv:28760:3
	function automatic [AddrWidth - 1:0] align_addr;
		// Trace: design.sv:28760:40
		input reg [AddrWidth - 1:0] addr;
		// Trace: design.sv:28761:5
		align_addr = (addr >> $clog2(DataBytes)) << $clog2(DataBytes);
	endfunction
	// Trace: design.sv:28765:3
	assign req_valid = req_i & gnt_o;
	// Trace: design.sv:28766:3
	genvar _gv_i_31;
	generate
		for (_gv_i_31 = 0; $unsigned(_gv_i_31) < NumBanks; _gv_i_31 = _gv_i_31 + 1) begin : gen_reqs
			localparam i = _gv_i_31;
			// Trace: design.sv:28767:5
			assign bank_req[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))))) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))))) + ((AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) >= ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) ? ((AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1)))) + 1 : (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) - (AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))))) + 1)) - 1)-:((AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) >= ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) ? ((AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1)))) + 1 : (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) - (AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))))) + 1)] = align_addr(addr_i) + (i * BytesPerBank);
			// Trace: design.sv:28768:5
			assign bank_req[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))))) + (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) >= (((DataWidth / NumBanks) / 8) + (AtopWidth + 1)) ? (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) + 1 : ((((DataWidth / NumBanks) / 8) + (AtopWidth + 1)) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) + 1)) - 1)-:(((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) >= (((DataWidth / NumBanks) / 8) + (AtopWidth + 1)) ? (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) + 1 : ((((DataWidth / NumBanks) / 8) + (AtopWidth + 1)) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) + 1)] = wdata_i[i * BitsPerBank+:BitsPerBank];
			// Trace: design.sv:28769:5
			assign bank_req[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? ((DataWidth / NumBanks) / 8) + (AtopWidth + 0) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? ((DataWidth / NumBanks) / 8) + (AtopWidth + 0) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) + ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) >= (AtopWidth + 1) ? ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) - (AtopWidth + 1)) + 1 : ((AtopWidth + 1) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) + 1)) - 1)-:((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) >= (AtopWidth + 1) ? ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) - (AtopWidth + 1)) + 1 : ((AtopWidth + 1) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) + 1)] = strb_i[i * BytesPerBank+:BytesPerBank];
			// Trace: design.sv:28770:5
			assign bank_req[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? AtopWidth + 0 : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (AtopWidth + 0)) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? AtopWidth + 0 : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (AtopWidth + 0))) + ((AtopWidth + 0) >= 1 ? AtopWidth + 0 : 2 - (AtopWidth + 0))) - 1)-:((AtopWidth + 0) >= 1 ? AtopWidth + 0 : 2 - (AtopWidth + 0))] = atop_i;
			// Trace: design.sv:28771:5
			assign bank_req[(i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? 0 : (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0)] = we_i;
			// Trace: design.sv:28772:5
			stream_fifo_30B4A_70D5B #(
				.T_AddrWidth(AddrWidth),
				.T_AtopWidth(AtopWidth),
				.T_DataWidth(DataWidth),
				.T_NumBanks(NumBanks),
				.FALL_THROUGH(1'b1),
				.DATA_WIDTH(1 * (((((0 + AddrWidth) + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1)),
				.DEPTH(FifoDepth)
			) i_ft_reg(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(1'b0),
				.usage_o(),
				.data_i(bank_req[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? 0 : (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) + (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0)))+:(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))]),
				.valid_i(req_valid),
				.ready_o(req_ready[i]),
				.data_o(bank_oup[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? 0 : (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) + (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0)))+:(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))]),
				.valid_o(bank_req_internal[i]),
				.ready_i(bank_gnt_internal[i])
			);
			// Trace: design.sv:28790:5
			assign bank_addr_o[i * AddrWidth+:AddrWidth] = bank_oup[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))))) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))))) + ((AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) >= ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) ? ((AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1)))) + 1 : (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) - (AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))))) + 1)) - 1)-:((AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) >= ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) ? ((AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1)))) + 1 : (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) - (AddrWidth + ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))))) + 1)];
			// Trace: design.sv:28791:5
			assign bank_wdata_o[i * (DataWidth / NumBanks)+:DataWidth / NumBanks] = bank_oup[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))))) + (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) >= (((DataWidth / NumBanks) / 8) + (AtopWidth + 1)) ? (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) + 1 : ((((DataWidth / NumBanks) / 8) + (AtopWidth + 1)) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) + 1)) - 1)-:(((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) >= (((DataWidth / NumBanks) / 8) + (AtopWidth + 1)) ? (((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 1))) + 1 : ((((DataWidth / NumBanks) / 8) + (AtopWidth + 1)) - ((DataWidth / NumBanks) + (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) + 1)];
			// Trace: design.sv:28792:5
			assign bank_strb_o[i * ((DataWidth / NumBanks) / 8)+:(DataWidth / NumBanks) / 8] = bank_oup[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? ((DataWidth / NumBanks) / 8) + (AtopWidth + 0) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? ((DataWidth / NumBanks) / 8) + (AtopWidth + 0) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) + ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) >= (AtopWidth + 1) ? ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) - (AtopWidth + 1)) + 1 : ((AtopWidth + 1) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) + 1)) - 1)-:((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) >= (AtopWidth + 1) ? ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) - (AtopWidth + 1)) + 1 : ((AtopWidth + 1) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) + 1)];
			// Trace: design.sv:28793:5
			assign bank_atop_o[i * AtopWidth+:AtopWidth] = bank_oup[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? AtopWidth + 0 : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (AtopWidth + 0)) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? AtopWidth + 0 : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (AtopWidth + 0))) + ((AtopWidth + 0) >= 1 ? AtopWidth + 0 : 2 - (AtopWidth + 0))) - 1)-:((AtopWidth + 0) >= 1 ? AtopWidth + 0 : 2 - (AtopWidth + 0))];
			// Trace: design.sv:28794:5
			assign bank_we_o[i] = bank_oup[(i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? 0 : (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0)];
			// Trace: design.sv:28796:5
			assign zero_strobe[i] = bank_oup[(((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? ((DataWidth / NumBanks) / 8) + (AtopWidth + 0) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) : (((i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? ((DataWidth / NumBanks) / 8) + (AtopWidth + 0) : ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0)))) + ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) >= (AtopWidth + 1) ? ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) - (AtopWidth + 1)) + 1 : ((AtopWidth + 1) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) + 1)) - 1)-:((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) >= (AtopWidth + 1) ? ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) - (AtopWidth + 1)) + 1 : ((AtopWidth + 1) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) + 1)] == {((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) >= (AtopWidth + 1) ? ((((DataWidth / NumBanks) / 8) + (AtopWidth + 0)) - (AtopWidth + 1)) + 1 : ((AtopWidth + 1) - (((DataWidth / NumBanks) / 8) + (AtopWidth + 0))) + 1) * 1 {1'sb0}};
			if (HideStrb) begin : gen_hide_strb
				// Trace: design.sv:28799:7
				assign bank_req_o[i] = (bank_oup[(i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? 0 : (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0)] && zero_strobe[i] ? 1'b0 : bank_req_internal[i]);
				// Trace: design.sv:28800:7
				assign bank_gnt_internal[i] = (bank_oup[(i * (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 1 : 1 - ((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0))) + (((((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0) >= 0 ? 0 : (((AddrWidth + (DataWidth / NumBanks)) + ((DataWidth / NumBanks) / 8)) + AtopWidth) + 0)] && zero_strobe[i] ? 1'b1 : bank_gnt_i[i]);
			end
			else begin : gen_legacy_strb
				// Trace: design.sv:28802:7
				assign bank_req_o[i] = bank_req_internal[i];
				// Trace: design.sv:28803:7
				assign bank_gnt_internal[i] = bank_gnt_i[i];
			end
		end
	endgenerate
	// Trace: design.sv:28808:3
	assign gnt_o = (&req_ready & (&resp_ready)) & !dead_write_fifo_full;
	// Trace: design.sv:28810:3
	generate
		if (HideStrb) begin : gen_dead_write_fifo
			// Trace: design.sv:28811:5
			fifo_v3 #(
				.FALL_THROUGH(1'b1),
				.DEPTH(MaxTrans + 1),
				.DATA_WIDTH(NumBanks)
			) i_dead_write_fifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(1'b0),
				.full_o(dead_write_fifo_full),
				.empty_o(),
				.usage_o(),
				.data_i(bank_we_o & zero_strobe),
				.push_i(req_i & gnt_o),
				.data_o(dead_response),
				.pop_i(rvalid_o)
			);
		end
		else begin : gen_no_dead_write_fifo
			// Trace: design.sv:28829:5
			assign dead_response = 1'sb0;
			// Trace: design.sv:28830:5
			assign dead_write_fifo_full = 1'b0;
		end
	endgenerate
	// Trace: design.sv:28834:3
	genvar _gv_i_32;
	generate
		for (_gv_i_32 = 0; $unsigned(_gv_i_32) < NumBanks; _gv_i_32 = _gv_i_32 + 1) begin : gen_resp_regs
			localparam i = _gv_i_32;
			// Trace: design.sv:28835:5
			stream_fifo_7F5E8_FC84F #(
				.T_DataWidth(DataWidth),
				.T_NumBanks(NumBanks),
				.FALL_THROUGH(1'b1),
				.DATA_WIDTH(DataWidth / NumBanks),
				.DEPTH(FifoDepth)
			) i_ft_reg(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(1'b0),
				.usage_o(),
				.data_i(bank_rdata_i[i * (DataWidth / NumBanks)+:DataWidth / NumBanks]),
				.valid_i(bank_rvalid_i[i]),
				.ready_o(resp_ready[i]),
				.data_o(rdata_o[i * BitsPerBank+:BitsPerBank]),
				.valid_o(resp_valid[i]),
				.ready_i(rvalid_o & !dead_response[i])
			);
		end
	endgenerate
	// Trace: design.sv:28854:3
	assign rvalid_o = &(resp_valid | dead_response);
endmodule
module stream_arbiter (
	clk_i,
	rst_ni,
	inp_data_i,
	inp_valid_i,
	inp_ready_o,
	oup_data_o,
	oup_valid_o,
	oup_ready_i
);
	// Trace: design.sv:28888:25
	// removed localparam type DATA_T
	// Trace: design.sv:28889:15
	parameter integer N_INP = -1;
	// Trace: design.sv:28890:25
	parameter ARBITER = "rr";
	// Trace: design.sv:28892:5
	input wire clk_i;
	// Trace: design.sv:28893:5
	input wire rst_ni;
	// Trace: design.sv:28895:5
	input wire [N_INP - 1:0] inp_data_i;
	// Trace: design.sv:28896:5
	input wire [N_INP - 1:0] inp_valid_i;
	// Trace: design.sv:28897:5
	output wire [N_INP - 1:0] inp_ready_o;
	// Trace: design.sv:28899:5
	output wire oup_data_o;
	// Trace: design.sv:28900:5
	output wire oup_valid_o;
	// Trace: design.sv:28901:5
	input wire oup_ready_i;
	// Trace: design.sv:28904:3
	stream_arbiter_flushable_8B6F2 #(
		.N_INP(N_INP),
		.ARBITER(ARBITER)
	) i_arb(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.inp_data_i(inp_data_i),
		.inp_valid_i(inp_valid_i),
		.inp_ready_o(inp_ready_o),
		.oup_data_o(oup_data_o),
		.oup_valid_o(oup_valid_o),
		.oup_ready_i(oup_ready_i)
	);
endmodule
module stream_omega_net (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	data_i,
	sel_i,
	valid_i,
	ready_o,
	data_o,
	idx_o,
	valid_o,
	ready_i
);
	// Trace: design.sv:28940:13
	parameter [31:0] NumInp = 32'd0;
	// Trace: design.sv:28942:13
	parameter [31:0] NumOut = 32'd0;
	// Trace: design.sv:28945:13
	parameter [31:0] Radix = 32'd2;
	// Trace: design.sv:28947:13
	parameter [31:0] DataWidth = 32'd1;
	// Trace: design.sv:28949:26
	// removed localparam type payload_t
	// Trace: design.sv:28951:13
	parameter [0:0] SpillReg = 1'b0;
	// Trace: design.sv:28953:13
	parameter [31:0] ExtPrio = 1'b0;
	// Trace: design.sv:28956:13
	parameter [31:0] AxiVldRdy = 1'b1;
	// Trace: design.sv:28960:13
	parameter [31:0] LockIn = 1'b1;
	// Trace: design.sv:28964:13
	parameter [31:0] SelWidth = (NumOut > 32'd1 ? $unsigned($clog2(NumOut)) : 32'd1);
	// Trace: design.sv:28968:18
	// removed localparam type sel_oup_t
	// Trace: design.sv:28972:13
	parameter [31:0] IdxWidth = (NumInp > 32'd1 ? $unsigned($clog2(NumInp)) : 32'd1);
	// Trace: design.sv:28976:18
	// removed localparam type idx_inp_t
	// Trace: design.sv:28979:3
	input wire clk_i;
	// Trace: design.sv:28981:3
	input wire rst_ni;
	// Trace: design.sv:28986:3
	input wire flush_i;
	// Trace: design.sv:28989:3
	input wire [(NumOut * IdxWidth) - 1:0] rr_i;
	// Trace: design.sv:28992:3
	input wire [(NumInp * DataWidth) - 1:0] data_i;
	// Trace: design.sv:28995:3
	input wire [(NumInp * SelWidth) - 1:0] sel_i;
	// Trace: design.sv:28997:3
	input wire [NumInp - 1:0] valid_i;
	// Trace: design.sv:28999:3
	output wire [NumInp - 1:0] ready_o;
	// Trace: design.sv:29001:3
	output wire [(NumOut * DataWidth) - 1:0] data_o;
	// Trace: design.sv:29003:3
	output wire [(NumOut * IdxWidth) - 1:0] idx_o;
	// Trace: design.sv:29005:3
	output wire [NumOut - 1:0] valid_o;
	// Trace: design.sv:29007:3
	input wire [NumOut - 1:0] ready_i;
	// Trace: design.sv:29009:3
	function automatic integer cf_math_pkg_ceil_div;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:23:42
		input reg signed [63:0] dividend;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:23:66
		input reg signed [63:0] divisor;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:24:9
		reg signed [63:0] remainder;
		begin
			// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:42:9
			remainder = dividend;
			// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:43:9
			for (cf_math_pkg_ceil_div = 0; remainder > 0; cf_math_pkg_ceil_div = cf_math_pkg_ceil_div + 1)
				begin
					// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:44:13
					remainder = remainder - divisor;
				end
		end
	endfunction
	function automatic [DataWidth - 1:0] sv2v_cast_8536A;
		input reg [DataWidth - 1:0] inp;
		sv2v_cast_8536A = inp;
	endfunction
	function automatic [IdxWidth - 1:0] sv2v_cast_5FDFE;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_5FDFE = inp;
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	generate
		if ((NumInp <= Radix) && (NumOut <= Radix)) begin : gen_degenerate_omega_net
			// Trace: design.sv:29012:5
			stream_xbar_67930_B7325 #(
				.payload_t_DataWidth(DataWidth),
				.NumInp(NumInp),
				.NumOut(NumOut),
				.OutSpillReg(SpillReg),
				.ExtPrio(ExtPrio),
				.AxiVldRdy(AxiVldRdy),
				.LockIn(LockIn)
			) i_stream_xbar(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.rr_i(rr_i),
				.data_i(data_i),
				.sel_i(sel_i),
				.valid_i(valid_i),
				.ready_o(ready_o),
				.data_o(data_o),
				.idx_o(idx_o),
				.valid_o(valid_o),
				.ready_i(ready_i)
			);
		end
		else begin : gen_omega_net
			// Trace: design.sv:29041:5
			localparam [31:0] NumLanes = (NumOut > NumInp ? $unsigned(Radix ** cf_math_pkg_ceil_div($clog2(NumOut), $clog2(Radix))) : $unsigned(Radix ** cf_math_pkg_ceil_div($clog2(NumInp), $clog2(Radix))));
			// Trace: design.sv:29046:5
			localparam [31:0] NumLevels = $unsigned((($clog2(NumLanes) + $clog2(Radix)) - 1) / $clog2(Radix));
			// Trace: design.sv:29050:5
			localparam [31:0] NumRouters = NumLanes / Radix;
			// Trace: design.sv:29058:5
			// removed localparam type sel_dst_t
			// Trace: design.sv:29061:5
			localparam [31:0] SelW = $unsigned($clog2(Radix));
			// Trace: design.sv:29062:5
			initial begin : proc_selw
				// Trace: design.sv:29063:7
				$display("SelW is:    %0d", SelW);
				// Trace: design.sv:29064:7
				$display("SelDstW is: %0d", $clog2(NumLanes));
			end
			// Trace: design.sv:29066:5
			// removed localparam type sel_t
			// Trace: design.sv:29069:5
			// removed localparam type omega_data_t
			// Trace: design.sv:29076:5
			wire [(((NumLevels * NumRouters) * Radix) * (($clog2(NumLanes) + DataWidth) + IdxWidth)) - 1:0] inp_router_data;
			// Trace: design.sv:29077:5
			wire [((NumLevels * NumRouters) * Radix) - 1:0] inp_router_valid;
			wire [((NumLevels * NumRouters) * Radix) - 1:0] inp_router_ready;
			// Trace: design.sv:29078:5
			wire [(((NumLevels * NumRouters) * Radix) * (($clog2(NumLanes) + DataWidth) + IdxWidth)) - 1:0] out_router_data;
			// Trace: design.sv:29079:5
			wire [((NumLevels * NumRouters) * Radix) - 1:0] out_router_valid;
			wire [((NumLevels * NumRouters) * Radix) - 1:0] out_router_ready;
			genvar _gv_i_33;
			for (_gv_i_33 = 0; $unsigned(_gv_i_33) < (NumLevels - 1); _gv_i_33 = _gv_i_33 + 1) begin : gen_shuffle_levels
				localparam i = _gv_i_33;
				genvar _gv_j_11;
				for (_gv_j_11 = 0; $unsigned(_gv_j_11) < NumRouters; _gv_j_11 = _gv_j_11 + 1) begin : gen_shuffle_routers
					localparam j = _gv_j_11;
					genvar _gv_k_7;
					for (_gv_k_7 = 0; $unsigned(_gv_k_7) < Radix; _gv_k_7 = _gv_k_7 + 1) begin : gen_shuffle_radix
						localparam k = _gv_k_7;
						// Trace: design.sv:29086:11
						localparam [31:0] IdxLane = (Radix * j) + k;
						// Trace: design.sv:29088:11
						assign inp_router_data[(((((i + 1) * NumRouters) + (IdxLane % NumRouters)) * Radix) + (IdxLane / NumRouters)) * (($clog2(NumLanes) + DataWidth) + IdxWidth)+:($clog2(NumLanes) + DataWidth) + IdxWidth] = out_router_data[((((i * NumRouters) + j) * Radix) + k) * (($clog2(NumLanes) + DataWidth) + IdxWidth)+:($clog2(NumLanes) + DataWidth) + IdxWidth];
						// Trace: design.sv:29091:11
						assign inp_router_valid[((((i + 1) * NumRouters) + (IdxLane % NumRouters)) * Radix) + (IdxLane / NumRouters)] = out_router_valid[(((i * NumRouters) + j) * Radix) + k];
						// Trace: design.sv:29094:11
						assign out_router_ready[(((i * NumRouters) + j) * Radix) + k] = inp_router_ready[((((i + 1) * NumRouters) + (IdxLane % NumRouters)) * Radix) + (IdxLane / NumRouters)];
						if (i == 0) begin : gen_shuffle_inp
							if ((NumLanes - IdxLane) <= NumInp) begin : gen_inp_ports
								// Trace: design.sv:29103:15
								localparam [31:0] IdxInp = (NumLanes - IdxLane) - 32'd1;
								// Trace: design.sv:29104:15
								function automatic [$clog2(NumLanes) - 1:0] sv2v_cast_51149;
									input reg [$clog2(NumLanes) - 1:0] inp;
									sv2v_cast_51149 = inp;
								endfunction
								assign inp_router_data[(((0 + (IdxLane % NumRouters)) * Radix) + (IdxLane / NumRouters)) * (($clog2(NumLanes) + DataWidth) + IdxWidth)+:($clog2(NumLanes) + DataWidth) + IdxWidth] = {sv2v_cast_51149(sel_i[IdxInp * SelWidth+:SelWidth]), sv2v_cast_8536A(data_i[IdxInp * DataWidth+:DataWidth]), sv2v_cast_5FDFE(IdxInp)};
								// Trace: design.sv:29110:15
								assign inp_router_valid[((0 + (IdxLane % NumRouters)) * Radix) + (IdxLane / NumRouters)] = valid_i[IdxInp];
								// Trace: design.sv:29111:15
								assign ready_o[IdxInp] = inp_router_ready[((0 + (IdxLane % NumRouters)) * Radix) + (IdxLane / NumRouters)];
							end
							else begin : gen_tie_off
								// Trace: design.sv:29114:15
								function automatic [$clog2(NumLanes) - 1:0] sv2v_cast_51149;
									input reg [$clog2(NumLanes) - 1:0] inp;
									sv2v_cast_51149 = inp;
								endfunction
								assign inp_router_data[(((0 + (IdxLane % NumRouters)) * Radix) + (IdxLane / NumRouters)) * (($clog2(NumLanes) + DataWidth) + IdxWidth)+:($clog2(NumLanes) + DataWidth) + IdxWidth] = {sv2v_cast_51149(1'sb0), sv2v_cast_8536A(1'sb0), sv2v_cast_5FDFE(1'sb0)};
								// Trace: design.sv:29115:15
								assign inp_router_valid[((0 + (IdxLane % NumRouters)) * Radix) + (IdxLane / NumRouters)] = 1'b0;
							end
						end
					end
				end
			end
			genvar _gv_i_34;
			for (_gv_i_34 = 0; $unsigned(_gv_i_34) < NumLevels; _gv_i_34 = _gv_i_34 + 1) begin : gen_router_levels
				localparam i = _gv_i_34;
				genvar _gv_j_12;
				for (_gv_j_12 = 0; $unsigned(_gv_j_12) < NumRouters; _gv_j_12 = _gv_j_12 + 1) begin : gen_routers
					localparam j = _gv_j_12;
					// Trace: design.sv:29125:9
					wire [(Radix * SelW) - 1:0] sel_router;
					genvar _gv_k_8;
					for (_gv_k_8 = 0; $unsigned(_gv_k_8) < Radix; _gv_k_8 = _gv_k_8 + 1) begin : gen_router_sel
						localparam k = _gv_k_8;
						// Trace: design.sv:29132:11
						assign sel_router[k * SelW+:SelW] = inp_router_data[(((((i * NumRouters) + j) * Radix) + k) * (($clog2(NumLanes) + DataWidth) + IdxWidth)) + (($clog2(NumLanes) + (DataWidth + (IdxWidth - 1))) - (($clog2(NumLanes) - 1) - (SelW * ((NumLevels - i) - 1))))+:SelW];
					end
					// Trace: design.sv:29135:9
					localparam integer i_stream_xbar_sv2v_pfunc_944F6 = $clog2(NumLanes);
					localparam [31:0] sv2v_uu_i_stream_xbar_NumInp = Radix;
					localparam [31:0] sv2v_uu_i_stream_xbar_IdxWidth = (sv2v_uu_i_stream_xbar_NumInp > 32'd1 ? $unsigned($clog2(sv2v_uu_i_stream_xbar_NumInp)) : 32'd1);
					localparam [31:0] sv2v_uu_i_stream_xbar_NumOut = Radix;
					// removed localparam type sv2v_uu_i_stream_xbar_rr_i
					localparam [(Radix * sv2v_cast_32((Radix > 32'd1 ? $unsigned($clog2(Radix)) : 32'd1))) - 1:0] sv2v_uu_i_stream_xbar_ext_rr_i_0 = 1'sb0;
					stream_xbar_09F43_1A7A9 #(
						.payload_t_DataWidth(DataWidth),
						.payload_t_IdxWidth(IdxWidth),
						.payload_t_i_stream_xbar_sv2v_pfunc_944F6(i_stream_xbar_sv2v_pfunc_944F6),
						.NumInp(Radix),
						.NumOut(Radix),
						.OutSpillReg(SpillReg),
						.ExtPrio(1'b0),
						.AxiVldRdy(AxiVldRdy),
						.LockIn(LockIn)
					) i_stream_xbar(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.flush_i(flush_i),
						.rr_i(sv2v_uu_i_stream_xbar_ext_rr_i_0),
						.data_i(inp_router_data[(($clog2(NumLanes) + DataWidth) + IdxWidth) * (((i * NumRouters) + j) * Radix)+:(($clog2(NumLanes) + DataWidth) + IdxWidth) * Radix]),
						.sel_i(sel_router),
						.valid_i(inp_router_valid[((i * NumRouters) + j) * Radix+:Radix]),
						.ready_o(inp_router_ready[((i * NumRouters) + j) * Radix+:Radix]),
						.data_o(out_router_data[(($clog2(NumLanes) + DataWidth) + IdxWidth) * (((i * NumRouters) + j) * Radix)+:(($clog2(NumLanes) + DataWidth) + IdxWidth) * Radix]),
						.idx_o(),
						.valid_o(out_router_valid[((i * NumRouters) + j) * Radix+:Radix]),
						.ready_i(out_router_ready[((i * NumRouters) + j) * Radix+:Radix])
					);
				end
			end
			genvar _gv_i_35;
			for (_gv_i_35 = 0; $unsigned(_gv_i_35) < NumLanes; _gv_i_35 = _gv_i_35 + 1) begin : gen_outputs
				localparam i = _gv_i_35;
				if (i < NumOut) begin : gen_connect
					// Trace: design.sv:29163:9
					assign data_o[i * DataWidth+:DataWidth] = out_router_data[((((((NumLevels - 1) * NumRouters) + (i / Radix)) * Radix) + (i % Radix)) * (($clog2(NumLanes) + DataWidth) + IdxWidth)) + (DataWidth + (IdxWidth - 1))-:((DataWidth + (IdxWidth - 1)) >= (IdxWidth + 0) ? ((DataWidth + (IdxWidth - 1)) - (IdxWidth + 0)) + 1 : ((IdxWidth + 0) - (DataWidth + (IdxWidth - 1))) + 1)];
					// Trace: design.sv:29164:9
					assign idx_o[i * IdxWidth+:IdxWidth] = out_router_data[((((((NumLevels - 1) * NumRouters) + (i / Radix)) * Radix) + (i % Radix)) * (($clog2(NumLanes) + DataWidth) + IdxWidth)) + (IdxWidth - 1)-:IdxWidth];
					// Trace: design.sv:29165:9
					assign valid_o[i] = out_router_valid[((((NumLevels - 1) * NumRouters) + (i / Radix)) * Radix) + (i % Radix)];
					// Trace: design.sv:29166:9
					assign out_router_ready[((((NumLevels - 1) * NumRouters) + (i / Radix)) * Radix) + (i % Radix)] = ready_i[i];
				end
				else begin : gen_tie_off
					// Trace: design.sv:29168:9
					assign out_router_ready[((((NumLevels - 1) * NumRouters) + (i / Radix)) * Radix) + (i % Radix)] = 1'b0;
				end
			end
			// Trace: design.sv:29172:5
			initial begin : proc_debug_print
				// Trace: design.sv:29173:7
				$display("NumInp:     %0d", NumInp);
				// Trace: design.sv:29174:7
				$display("NumOut:     %0d", NumOut);
				// Trace: design.sv:29175:7
				$display("Radix:      %0d", Radix);
				// Trace: design.sv:29176:7
				$display("NumLanes:   %0d", NumLanes);
				// Trace: design.sv:29177:7
				$display("NumLevels:  %0d", NumLevels);
				// Trace: design.sv:29178:7
				$display("NumRouters: %0d", NumRouters);
			end
		end
	endgenerate
endmodule
module clock_divider_counter (
	clk,
	rstn,
	test_mode,
	clk_div,
	clk_div_valid,
	clk_out
);
	reg _sv2v_0;
	// Trace: design.sv:29266:15
	parameter BYPASS_INIT = 1;
	// Trace: design.sv:29267:15
	parameter DIV_INIT = 'hff;
	// Trace: design.sv:29270:5
	input wire clk;
	// Trace: design.sv:29271:5
	input wire rstn;
	// Trace: design.sv:29272:5
	input wire test_mode;
	// Trace: design.sv:29273:5
	input wire [7:0] clk_div;
	// Trace: design.sv:29274:5
	input wire clk_div_valid;
	// Trace: design.sv:29275:5
	output wire clk_out;
	// Trace: design.sv:29278:5
	reg [7:0] counter;
	// Trace: design.sv:29279:5
	reg [7:0] counter_next;
	// Trace: design.sv:29280:5
	reg [7:0] clk_cnt;
	// Trace: design.sv:29281:5
	reg en1;
	// Trace: design.sv:29282:5
	reg en2;
	// Trace: design.sv:29284:5
	reg is_odd;
	// Trace: design.sv:29286:5
	reg div1;
	// Trace: design.sv:29287:5
	reg div2;
	// Trace: design.sv:29288:5
	wire div2_neg_sync;
	// Trace: design.sv:29290:5
	wire [7:0] clk_cnt_odd;
	// Trace: design.sv:29291:5
	wire [7:0] clk_cnt_odd_incr;
	// Trace: design.sv:29292:5
	wire [7:0] clk_cnt_even;
	// Trace: design.sv:29293:5
	wire [7:0] clk_cnt_en2;
	// Trace: design.sv:29295:5
	reg bypass;
	// Trace: design.sv:29297:5
	wire clk_out_gen;
	// Trace: design.sv:29298:5
	reg clk_div_valid_reg;
	// Trace: design.sv:29300:5
	wire clk_inv_test;
	// Trace: design.sv:29301:5
	wire clk_inv;
	// Trace: design.sv:29305:5
	assign clk_cnt_odd = clk_div - 8'h01;
	// Trace: design.sv:29306:5
	assign clk_cnt_even = (clk_div == 8'h02 ? 8'h00 : {1'b0, clk_div[7:1]} - 8'h01);
	// Trace: design.sv:29307:5
	assign clk_cnt_en2 = {1'b0, clk_cnt[7:1]} + 8'h01;
	// Trace: design.sv:29309:5
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:29311:9
		if (counter == 'h0)
			// Trace: design.sv:29312:13
			en1 = 1'b1;
		else
			// Trace: design.sv:29314:13
			en1 = 1'b0;
		if (clk_div_valid)
			// Trace: design.sv:29317:13
			counter_next = 'h0;
		else if (counter == clk_cnt)
			// Trace: design.sv:29319:17
			counter_next = 'h0;
		else
			// Trace: design.sv:29321:17
			counter_next = counter + 1;
		if (clk_div_valid)
			// Trace: design.sv:29324:13
			en2 = 1'b0;
		else if (counter == clk_cnt_en2)
			// Trace: design.sv:29326:17
			en2 = 1'b1;
		else
			// Trace: design.sv:29328:17
			en2 = 1'b0;
	end
	// Trace: design.sv:29331:4
	always @(posedge clk or negedge rstn)
		// Trace: design.sv:29333:9
		if (~rstn) begin
			// Trace: design.sv:29335:14
			counter <= 'h0;
			// Trace: design.sv:29336:14
			div1 <= 1'b0;
			// Trace: design.sv:29337:14
			bypass <= BYPASS_INIT;
			// Trace: design.sv:29338:14
			clk_cnt <= DIV_INIT;
			// Trace: design.sv:29339:14
			is_odd <= 1'b0;
			// Trace: design.sv:29340:14
			clk_div_valid_reg <= 1'b0;
		end
		else begin
			// Trace: design.sv:29344:15
			if (!bypass)
				// Trace: design.sv:29345:19
				counter <= counter_next;
			// Trace: design.sv:29347:15
			clk_div_valid_reg <= clk_div_valid;
			if (clk_div_valid) begin
				// Trace: design.sv:29350:17
				if ((clk_div == 8'h00) || (clk_div == 8'h01)) begin
					// Trace: design.sv:29352:23
					bypass <= 1'b1;
					// Trace: design.sv:29353:23
					clk_cnt <= 'h0;
					// Trace: design.sv:29354:23
					is_odd <= 1'b0;
				end
				else begin
					// Trace: design.sv:29358:23
					bypass <= 1'b0;
					// Trace: design.sv:29359:23
					if (clk_div[0]) begin
						// Trace: design.sv:29361:27
						is_odd <= 1'b1;
						// Trace: design.sv:29362:27
						clk_cnt <= clk_cnt_odd;
					end
					else begin
						// Trace: design.sv:29366:27
						is_odd <= 1'b0;
						// Trace: design.sv:29367:27
						clk_cnt <= clk_cnt_even;
					end
				end
				// Trace: design.sv:29370:17
				div1 <= 1'b0;
			end
			else
				// Trace: design.sv:29374:17
				if (en1 && !bypass)
					// Trace: design.sv:29375:19
					div1 <= ~div1;
		end
	// Trace: design.sv:29380:5
	pulp_clock_inverter clk_inv_i(
		.clk_i(clk),
		.clk_o(clk_inv)
	);
	// Trace: design.sv:29396:4
	assign clk_inv_test = clk_inv;
	// Trace: design.sv:29402:5
	always @(posedge clk_inv_test or negedge rstn)
		// Trace: design.sv:29404:9
		if (!rstn)
			// Trace: design.sv:29406:13
			div2 <= 1'b0;
		else
			// Trace: design.sv:29410:13
			if (clk_div_valid_reg)
				// Trace: design.sv:29411:17
				div2 <= 1'b0;
			else if ((en2 && is_odd) && !bypass)
				// Trace: design.sv:29413:21
				div2 <= ~div2;
	// Trace: design.sv:29417:5
	pulp_clock_xor2 clock_xor_i(
		.clk_o(clk_out_gen),
		.clk0_i(div1),
		.clk1_i(div2)
	);
	// Trace: design.sv:29424:5
	pulp_clock_mux2 clk_mux_i(
		.clk0_i(clk_out_gen),
		.clk1_i(clk),
		.clk_sel_i(bypass || test_mode),
		.clk_o(clk_out)
	);
	initial _sv2v_0 = 0;
endmodule
module clk_div (
	clk_i,
	rst_ni,
	testmode_i,
	en_i,
	clk_o
);
	// Trace: design.sv:29446:15
	parameter [31:0] RATIO = 4;
	// Trace: design.sv:29447:15
	parameter [0:0] SHOW_WARNING = 1'b1;
	// Trace: design.sv:29449:5
	input wire clk_i;
	// Trace: design.sv:29450:5
	input wire rst_ni;
	// Trace: design.sv:29451:5
	input wire testmode_i;
	// Trace: design.sv:29452:5
	input wire en_i;
	// Trace: design.sv:29453:5
	output wire clk_o;
	// Trace: design.sv:29455:5
	reg [RATIO - 1:0] counter_q;
	// Trace: design.sv:29456:5
	reg clk_q;
	// Trace: design.sv:29458:5
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:29459:9
		if (~rst_ni) begin
			// Trace: design.sv:29460:13
			clk_q <= 1'b0;
			// Trace: design.sv:29461:13
			counter_q <= 1'sb0;
		end
		else begin
			// Trace: design.sv:29463:13
			clk_q <= 1'b0;
			// Trace: design.sv:29464:13
			if (en_i) begin
				begin
					// Trace: design.sv:29465:17
					if (counter_q == (RATIO[RATIO - 1:0] - 1))
						// Trace: design.sv:29466:21
						clk_q <= 1'b1;
					else
						// Trace: design.sv:29468:21
						counter_q <= counter_q + 1;
				end
			end
		end
	// Trace: design.sv:29474:5
	assign clk_o = (testmode_i ? clk_i : clk_q);
	// Trace: design.sv:29476:3
	generate
		if (SHOW_WARNING) begin : gen_elab_warning
			// Trace: design.sv:29477:5
			$warning("This clock divider is deprecated and not reccomended since  ", "the generated output clock has a very unbalanced duty cycle  ", "(1/RATIO). For new designs we reccomend using the at-runtime ", "configurable clk_int_div module which always generates 50%%  ", "duty cycle clock. If you don't need at runtime configuration ", "support, you can instantiate clk_int_div as follows to       ", "obtain a module with roughly the same behavior (except for   ", "the 50 %% duty cycle):\n                                     ", "\n                                                           ", "  clk_int_div #(\n                                           ", "    .DIV_VALUE_WIDTH($clog2(RATIO+1)),\n                     ", "    .DEFAULT_DIV_VALUE(RATIO)\n                              ", "  ) i_clk_int_div(\n                                         ", "    .clk_i,\n                                                ", "    .rst_ni,\n                                               ", "    .test_mode_en_i(testmode_i),\n                           ", "    .en_i,\n                                                 ", "    .div_i('1), // Ignored, used default value\n             ", "    .div_valid_i(1'b0),\n                                    ", "    .div_ready_o(),\n                                        ", "    .clk_o\n                                                 ", "  );                                                         ", "\n                                                           ", "If you know what your are doing and want to disable this     ", "warning message, you can disable it by overriding the new    ", "optional clk_div parameter SHOW_WARNING to 1'b0.");
		end
	endgenerate
endmodule
module find_first_one (
	in_i,
	first_one_o,
	no_ones_o
);
	// Trace: design.sv:29525:15
	parameter signed [31:0] WIDTH = -1;
	// Trace: design.sv:29526:15
	parameter signed [31:0] FLIP = 0;
	// Trace: design.sv:29528:5
	input wire [WIDTH - 1:0] in_i;
	// Trace: design.sv:29529:5
	output wire [$clog2(WIDTH) - 1:0] first_one_o;
	// Trace: design.sv:29530:5
	output wire no_ones_o;
	// Trace: design.sv:29533:5
	localparam signed [31:0] NUM_LEVELS = $clog2(WIDTH);
	// Trace: design.sv:29536:5
	initial begin
		// Trace: design.sv:29537:9
		assert (WIDTH >= 0) ;
	end
	// Trace: design.sv:29541:5
	wire [(WIDTH * NUM_LEVELS) - 1:0] index_lut;
	// Trace: design.sv:29542:5
	wire [(2 ** NUM_LEVELS) - 1:0] sel_nodes;
	// Trace: design.sv:29543:5
	wire [((2 ** NUM_LEVELS) * NUM_LEVELS) - 1:0] index_nodes;
	// Trace: design.sv:29545:5
	wire [WIDTH - 1:0] in_tmp;
	// Trace: design.sv:29547:5
	genvar _gv_i_36;
	generate
		for (_gv_i_36 = 0; _gv_i_36 < WIDTH; _gv_i_36 = _gv_i_36 + 1) begin : genblk1
			localparam i = _gv_i_36;
			// Trace: design.sv:29548:9
			assign in_tmp[i] = (FLIP ? in_i[(WIDTH - 1) - i] : in_i[i]);
		end
	endgenerate
	// Trace: design.sv:29551:5
	genvar _gv_j_13;
	generate
		for (_gv_j_13 = 0; _gv_j_13 < WIDTH; _gv_j_13 = _gv_j_13 + 1) begin : genblk2
			localparam j = _gv_j_13;
			// Trace: design.sv:29552:9
			assign index_lut[j * NUM_LEVELS+:NUM_LEVELS] = j;
		end
	endgenerate
	// Trace: design.sv:29555:5
	genvar _gv_level_4;
	generate
		for (_gv_level_4 = 0; _gv_level_4 < NUM_LEVELS; _gv_level_4 = _gv_level_4 + 1) begin : genblk3
			localparam level = _gv_level_4;
			if (level < (NUM_LEVELS - 1)) begin : genblk1
				genvar _gv_l_6;
				for (_gv_l_6 = 0; _gv_l_6 < (2 ** level); _gv_l_6 = _gv_l_6 + 1) begin : genblk1
					localparam l = _gv_l_6;
					// Trace: design.sv:29559:17
					assign sel_nodes[((2 ** level) - 1) + l] = sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] | sel_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) + 1];
					// Trace: design.sv:29560:17
					assign index_nodes[(((2 ** level) - 1) + l) * NUM_LEVELS+:NUM_LEVELS] = (sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] == 1'b1 ? index_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) * NUM_LEVELS+:NUM_LEVELS] : index_nodes[((((2 ** (level + 1)) - 1) + (l * 2)) + 1) * NUM_LEVELS+:NUM_LEVELS]);
				end
			end
			if (level == (NUM_LEVELS - 1)) begin : genblk2
				genvar _gv_k_9;
				for (_gv_k_9 = 0; _gv_k_9 < (2 ** level); _gv_k_9 = _gv_k_9 + 1) begin : genblk1
					localparam k = _gv_k_9;
					if ((k * 2) < (WIDTH - 1)) begin : genblk1
						// Trace: design.sv:29569:21
						assign sel_nodes[((2 ** level) - 1) + k] = in_tmp[k * 2] | in_tmp[(k * 2) + 1];
						// Trace: design.sv:29570:21
						assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = (in_tmp[k * 2] == 1'b1 ? index_lut[(k * 2) * NUM_LEVELS+:NUM_LEVELS] : index_lut[((k * 2) + 1) * NUM_LEVELS+:NUM_LEVELS]);
					end
					if ((k * 2) == (WIDTH - 1)) begin : genblk2
						// Trace: design.sv:29574:21
						assign sel_nodes[((2 ** level) - 1) + k] = in_tmp[k * 2];
						// Trace: design.sv:29575:21
						assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = index_lut[(k * 2) * NUM_LEVELS+:NUM_LEVELS];
					end
					if ((k * 2) > (WIDTH - 1)) begin : genblk3
						// Trace: design.sv:29579:21
						assign sel_nodes[((2 ** level) - 1) + k] = 1'b0;
						// Trace: design.sv:29580:21
						assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = 1'sb0;
					end
				end
			end
		end
	endgenerate
	// Trace: design.sv:29586:5
	assign first_one_o = (NUM_LEVELS > 0 ? index_nodes[0+:NUM_LEVELS] : {$clog2(WIDTH) {1'sb0}});
	// Trace: design.sv:29587:5
	assign no_ones_o = (NUM_LEVELS > 0 ? ~sel_nodes[0] : 1'b1);
endmodule
module generic_LFSR_8bit (
	data_OH_o,
	data_BIN_o,
	enable_i,
	clk,
	rst_n
);
	reg _sv2v_0;
	// Trace: design.sv:29604:15
	parameter OH_WIDTH = 4;
	// Trace: design.sv:29605:15
	parameter BIN_WIDTH = $clog2(OH_WIDTH);
	// Trace: design.sv:29606:15
	parameter SEED = 8'b00000000;
	// Trace: design.sv:29609:5
	output reg [OH_WIDTH - 1:0] data_OH_o;
	// Trace: design.sv:29610:5
	output wire [BIN_WIDTH - 1:0] data_BIN_o;
	// Trace: design.sv:29611:5
	input wire enable_i;
	// Trace: design.sv:29612:5
	input wire clk;
	// Trace: design.sv:29613:5
	input wire rst_n;
	// Trace: design.sv:29616:4
	reg [7:0] out;
	// Trace: design.sv:29617:4
	wire linear_feedback;
	// Trace: design.sv:29618:4
	wire [BIN_WIDTH - 1:0] temp_ref_way;
	// Trace: design.sv:29622:4
	assign linear_feedback = !(((out[7] ^ out[3]) ^ out[2]) ^ out[1]);
	// Trace: design.sv:29624:4
	assign data_BIN_o = temp_ref_way;
	// Trace: design.sv:29626:4
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:29628:2
		if (rst_n == 1'b0)
			// Trace: design.sv:29630:7
			out <= SEED;
		else if (enable_i)
			// Trace: design.sv:29634:14
			out <= {out[6], out[5], out[4], out[3], out[2], out[1], out[0], linear_feedback};
	// Trace: design.sv:29638:4
	generate
		if (OH_WIDTH == 2) begin : genblk1
			// Trace: design.sv:29641:2
			assign temp_ref_way = out[1];
		end
		else begin : genblk1
			// Trace: design.sv:29643:2
			assign temp_ref_way = out[BIN_WIDTH:1];
		end
	endgenerate
	// Trace: design.sv:29647:4
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:29649:2
		data_OH_o = 1'sb0;
		// Trace: design.sv:29650:2
		data_OH_o[temp_ref_way] = 1'b1;
	end
	initial _sv2v_0 = 0;
endmodule
module generic_fifo (
	clk,
	rst_n,
	data_i,
	valid_i,
	grant_o,
	data_o,
	valid_o,
	grant_i,
	test_mode_i
);
	reg _sv2v_0;
	// Trace: design.sv:29693:14
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:29694:14
	parameter [31:0] DATA_DEPTH = 8;
	// Trace: design.sv:29697:4
	input wire clk;
	// Trace: design.sv:29698:4
	input wire rst_n;
	// Trace: design.sv:29700:4
	input wire [DATA_WIDTH - 1:0] data_i;
	// Trace: design.sv:29701:4
	input wire valid_i;
	// Trace: design.sv:29702:4
	output reg grant_o;
	// Trace: design.sv:29704:4
	output wire [DATA_WIDTH - 1:0] data_o;
	// Trace: design.sv:29705:4
	output reg valid_o;
	// Trace: design.sv:29706:4
	input wire grant_i;
	// Trace: design.sv:29708:4
	input wire test_mode_i;
	// Trace: design.sv:29713:4
	localparam [31:0] ADDR_DEPTH = $clog2(DATA_DEPTH);
	// Trace: design.sv:29714:4
	reg [1:0] CS;
	reg [1:0] NS;
	// Trace: design.sv:29717:4
	reg gate_clock;
	// Trace: design.sv:29718:4
	wire clk_gated;
	// Trace: design.sv:29720:4
	reg [ADDR_DEPTH - 1:0] Pop_Pointer_CS;
	reg [ADDR_DEPTH - 1:0] Pop_Pointer_NS;
	// Trace: design.sv:29721:4
	reg [ADDR_DEPTH - 1:0] Push_Pointer_CS;
	reg [ADDR_DEPTH - 1:0] Push_Pointer_NS;
	// Trace: design.sv:29722:4
	reg [DATA_WIDTH - 1:0] FIFO_REGISTERS [DATA_DEPTH - 1:0];
	// Trace: design.sv:29723:4
	reg [31:0] i;
	// Trace: design.sv:29727:4
	initial begin : parameter_check
		// Trace: design.sv:29728:7
		integer param_err_flg;
		// Trace: design.sv:29729:7
		param_err_flg = 0;
		// Trace: design.sv:29731:7
		if (DATA_WIDTH < 1) begin
			// Trace: design.sv:29732:10
			param_err_flg = 1;
			// Trace: design.sv:29733:10
			$display("ERROR: %m :\n  Invalid value (%d) for parameter DATA_WIDTH (legal range: greater than 1)", DATA_WIDTH);
		end
		if (DATA_DEPTH < 1) begin
			// Trace: design.sv:29737:10
			param_err_flg = 1;
			// Trace: design.sv:29738:10
			$display("ERROR: %m :\n  Invalid value (%d) for parameter DATA_DEPTH (legal range: greater than 1)", DATA_DEPTH);
		end
	end
	// Trace: design.sv:29744:4
	cluster_clock_gating cg_cell(
		.clk_i(clk),
		.en_i(~gate_clock),
		.test_en_i(test_mode_i),
		.clk_o(clk_gated)
	);
	// Trace: design.sv:29756:4
	always @(posedge clk or negedge rst_n)
		// Trace: design.sv:29758:8
		if (rst_n == 1'b0) begin
			// Trace: design.sv:29760:16
			CS <= 2'd0;
			// Trace: design.sv:29761:16
			Pop_Pointer_CS <= {ADDR_DEPTH {1'b0}};
			// Trace: design.sv:29762:16
			Push_Pointer_CS <= {ADDR_DEPTH {1'b0}};
		end
		else begin
			// Trace: design.sv:29766:16
			CS <= NS;
			// Trace: design.sv:29767:16
			Pop_Pointer_CS <= Pop_Pointer_NS;
			// Trace: design.sv:29768:16
			Push_Pointer_CS <= Push_Pointer_NS;
		end
	// Trace: design.sv:29774:4
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:29776:7
		gate_clock = 1'b0;
		// Trace: design.sv:29778:7
		case (CS)
			2'd0: begin
				// Trace: design.sv:29782:11
				grant_o = 1'b1;
				// Trace: design.sv:29783:11
				valid_o = 1'b0;
				// Trace: design.sv:29785:11
				case (valid_i)
					1'b0: begin
						// Trace: design.sv:29788:19
						NS = 2'd0;
						// Trace: design.sv:29789:19
						Push_Pointer_NS = Push_Pointer_CS;
						// Trace: design.sv:29790:19
						Pop_Pointer_NS = Pop_Pointer_CS;
						// Trace: design.sv:29791:19
						gate_clock = 1'b1;
					end
					1'b1: begin
						// Trace: design.sv:29796:19
						NS = 2'd2;
						// Trace: design.sv:29797:19
						Push_Pointer_NS = Push_Pointer_CS + 1'b1;
						// Trace: design.sv:29798:19
						Pop_Pointer_NS = Pop_Pointer_CS;
					end
				endcase
			end
			2'd2: begin
				// Trace: design.sv:29806:11
				grant_o = 1'b1;
				// Trace: design.sv:29807:11
				valid_o = 1'b1;
				// Trace: design.sv:29809:11
				case ({valid_i, grant_i})
					2'b01: begin
						// Trace: design.sv:29813:19
						gate_clock = 1'b1;
						// Trace: design.sv:29815:19
						if ((Pop_Pointer_CS == (Push_Pointer_CS - 1)) || ((Pop_Pointer_CS == (DATA_DEPTH - 1)) && (Push_Pointer_CS == 0)))
							// Trace: design.sv:29816:27
							NS = 2'd0;
						else
							// Trace: design.sv:29818:27
							NS = 2'd2;
						// Trace: design.sv:29820:19
						Push_Pointer_NS = Push_Pointer_CS;
						if (Pop_Pointer_CS == (DATA_DEPTH - 1))
							// Trace: design.sv:29823:27
							Pop_Pointer_NS = 0;
						else
							// Trace: design.sv:29825:27
							Pop_Pointer_NS = Pop_Pointer_CS + 1'b1;
					end
					2'b00: begin
						// Trace: design.sv:29830:19
						gate_clock = 1'b1;
						// Trace: design.sv:29831:19
						NS = 2'd2;
						// Trace: design.sv:29832:19
						Push_Pointer_NS = Push_Pointer_CS;
						// Trace: design.sv:29833:19
						Pop_Pointer_NS = Pop_Pointer_CS;
					end
					2'b11: begin
						// Trace: design.sv:29838:19
						NS = 2'd2;
						// Trace: design.sv:29840:19
						if (Push_Pointer_CS == (DATA_DEPTH - 1))
							// Trace: design.sv:29841:27
							Push_Pointer_NS = 0;
						else
							// Trace: design.sv:29843:27
							Push_Pointer_NS = Push_Pointer_CS + 1'b1;
						if (Pop_Pointer_CS == (DATA_DEPTH - 1))
							// Trace: design.sv:29846:27
							Pop_Pointer_NS = 0;
						else
							// Trace: design.sv:29848:27
							Pop_Pointer_NS = Pop_Pointer_CS + 1'b1;
					end
					2'b10: begin
						// Trace: design.sv:29853:19
						if ((Push_Pointer_CS == (Pop_Pointer_CS - 1)) || ((Push_Pointer_CS == (DATA_DEPTH - 1)) && (Pop_Pointer_CS == 0)))
							// Trace: design.sv:29854:27
							NS = 2'd1;
						else
							// Trace: design.sv:29856:27
							NS = 2'd2;
						if (Push_Pointer_CS == (DATA_DEPTH - 1))
							// Trace: design.sv:29859:27
							Push_Pointer_NS = 0;
						else
							// Trace: design.sv:29861:27
							Push_Pointer_NS = Push_Pointer_CS + 1'b1;
						// Trace: design.sv:29863:19
						Pop_Pointer_NS = Pop_Pointer_CS;
					end
				endcase
			end
			2'd1: begin
				// Trace: design.sv:29871:11
				grant_o = 1'b0;
				// Trace: design.sv:29872:11
				valid_o = 1'b1;
				// Trace: design.sv:29873:11
				gate_clock = 1'b1;
				// Trace: design.sv:29875:11
				case (grant_i)
					1'b1: begin
						// Trace: design.sv:29878:19
						NS = 2'd2;
						// Trace: design.sv:29880:19
						Push_Pointer_NS = Push_Pointer_CS;
						// Trace: design.sv:29882:19
						if (Pop_Pointer_CS == (DATA_DEPTH - 1))
							// Trace: design.sv:29883:27
							Pop_Pointer_NS = 0;
						else
							// Trace: design.sv:29885:27
							Pop_Pointer_NS = Pop_Pointer_CS + 1'b1;
					end
					1'b0: begin
						// Trace: design.sv:29890:19
						NS = 2'd1;
						// Trace: design.sv:29891:19
						Push_Pointer_NS = Push_Pointer_CS;
						// Trace: design.sv:29892:19
						Pop_Pointer_NS = Pop_Pointer_CS;
					end
				endcase
			end
			default: begin
				// Trace: design.sv:29900:11
				gate_clock = 1'b1;
				// Trace: design.sv:29901:11
				grant_o = 1'b0;
				// Trace: design.sv:29902:11
				valid_o = 1'b0;
				// Trace: design.sv:29903:11
				NS = 2'd0;
				// Trace: design.sv:29904:11
				Pop_Pointer_NS = 0;
				// Trace: design.sv:29905:11
				Push_Pointer_NS = 0;
			end
		endcase
	end
	// Trace: design.sv:29911:4
	always @(posedge clk_gated or negedge rst_n)
		// Trace: design.sv:29913:7
		if (rst_n == 1'b0)
			// Trace: design.sv:29915:7
			for (i = 0; i < DATA_DEPTH; i = i + 1)
				begin
					// Trace: design.sv:29916:10
					FIFO_REGISTERS[i] <= {DATA_WIDTH {1'b0}};
				end
		else
			// Trace: design.sv:29920:10
			if ((grant_o == 1'b1) && (valid_i == 1'b1))
				// Trace: design.sv:29921:13
				FIFO_REGISTERS[Push_Pointer_CS] <= data_i;
	// Trace: design.sv:29925:4
	assign data_o = FIFO_REGISTERS[Pop_Pointer_CS];
	initial _sv2v_0 = 0;
endmodule
module prioarbiter (
	clk_i,
	rst_ni,
	flush_i,
	en_i,
	req_i,
	ack_o,
	vld_o,
	idx_o
);
	// Trace: design.sv:29946:13
	parameter [31:0] NUM_REQ = 13;
	// Trace: design.sv:29947:13
	parameter [31:0] LOCK_IN = 0;
	// Trace: design.sv:29949:3
	input wire clk_i;
	// Trace: design.sv:29950:3
	input wire rst_ni;
	// Trace: design.sv:29952:3
	input wire flush_i;
	// Trace: design.sv:29953:3
	input wire en_i;
	// Trace: design.sv:29954:3
	input wire [NUM_REQ - 1:0] req_i;
	// Trace: design.sv:29956:3
	output wire [NUM_REQ - 1:0] ack_o;
	// Trace: design.sv:29957:3
	output wire vld_o;
	// Trace: design.sv:29958:3
	output wire [$clog2(NUM_REQ) - 1:0] idx_o;
	// Trace: design.sv:29961:3
	localparam SEL_WIDTH = $clog2(NUM_REQ);
	// Trace: design.sv:29963:3
	wire [SEL_WIDTH - 1:0] arb_sel_lock_d;
	reg [SEL_WIDTH - 1:0] arb_sel_lock_q;
	// Trace: design.sv:29964:3
	wire lock_d;
	reg lock_q;
	// Trace: design.sv:29966:3
	wire [$clog2(NUM_REQ) - 1:0] idx;
	// Trace: design.sv:29969:3
	assign vld_o = |req_i & en_i;
	// Trace: design.sv:29970:3
	assign idx_o = (lock_q ? arb_sel_lock_q : idx);
	// Trace: design.sv:29974:3
	assign ack_o[0] = (req_i[0] ? en_i : 1'b0);
	// Trace: design.sv:29976:3
	genvar _gv_i_37;
	generate
		for (_gv_i_37 = 1; _gv_i_37 < NUM_REQ; _gv_i_37 = _gv_i_37 + 1) begin : gen_arb_req_ports
			localparam i = _gv_i_37;
			// Trace: design.sv:29978:7
			assign ack_o[i] = (req_i[i] & ~(|ack_o[i - 1:0]) ? en_i : 1'b0);
		end
	endgenerate
	// Trace: design.sv:29981:3
	onehot_to_bin #(.ONEHOT_WIDTH(NUM_REQ)) i_onehot_to_bin(
		.onehot(ack_o),
		.bin(idx)
	);
	// Trace: design.sv:29988:3
	generate
		if (LOCK_IN) begin : gen_lock_in
			// Trace: design.sv:29990:5
			assign lock_d = |req_i & ~en_i;
			// Trace: design.sv:29991:5
			assign arb_sel_lock_d = idx_o;
		end
		else begin : genblk2
			// Trace: design.sv:29994:5
			assign lock_d = 1'sb0;
			// Trace: design.sv:29995:5
			assign arb_sel_lock_d = 1'sb0;
		end
	endgenerate
	// Trace: design.sv:29998:3
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:29999:5
		if (!rst_ni) begin
			// Trace: design.sv:30000:7
			lock_q <= 1'b0;
			// Trace: design.sv:30001:7
			arb_sel_lock_q <= 1'sb0;
		end
		else
			// Trace: design.sv:30003:7
			if (flush_i) begin
				// Trace: design.sv:30004:9
				lock_q <= 1'b0;
				// Trace: design.sv:30005:9
				arb_sel_lock_q <= 1'sb0;
			end
			else begin
				// Trace: design.sv:30007:9
				lock_q <= lock_d;
				// Trace: design.sv:30008:9
				arb_sel_lock_q <= arb_sel_lock_d;
			end
	end
endmodule
module pulp_sync (
	clk_i,
	rstn_i,
	serial_i,
	serial_o
);
	// Trace: design.sv:30031:15
	parameter STAGES = 2;
	// Trace: design.sv:30034:5
	input wire clk_i;
	// Trace: design.sv:30035:5
	input wire rstn_i;
	// Trace: design.sv:30036:5
	input wire serial_i;
	// Trace: design.sv:30037:5
	output wire serial_o;
	// Trace: design.sv:30040:4
	reg [STAGES - 1:0] r_reg;
	// Trace: design.sv:30042:4
	always @(posedge clk_i or negedge rstn_i)
		// Trace: design.sv:30044:2
		if (!rstn_i)
			// Trace: design.sv:30045:11
			r_reg <= 'h0;
		else
			// Trace: design.sv:30047:11
			r_reg <= {r_reg[STAGES - 2:0], serial_i};
	// Trace: design.sv:30050:4
	assign serial_o = r_reg[STAGES - 1];
endmodule
module pulp_sync_wedge (
	clk_i,
	rstn_i,
	en_i,
	serial_i,
	r_edge_o,
	f_edge_o,
	serial_o
);
	// Trace: design.sv:30066:15
	parameter [31:0] STAGES = 2;
	// Trace: design.sv:30068:5
	input wire clk_i;
	// Trace: design.sv:30069:5
	input wire rstn_i;
	// Trace: design.sv:30070:5
	input wire en_i;
	// Trace: design.sv:30071:5
	input wire serial_i;
	// Trace: design.sv:30072:5
	output wire r_edge_o;
	// Trace: design.sv:30073:5
	output wire f_edge_o;
	// Trace: design.sv:30074:5
	output wire serial_o;
	// Trace: design.sv:30076:5
	wire clk;
	// Trace: design.sv:30077:5
	wire serial;
	reg serial_q;
	// Trace: design.sv:30079:5
	assign serial_o = serial_q;
	// Trace: design.sv:30080:5
	assign f_edge_o = ~serial & serial_q;
	// Trace: design.sv:30081:5
	assign r_edge_o = serial & ~serial_q;
	// Trace: design.sv:30083:5
	pulp_sync #(.STAGES(STAGES)) i_pulp_sync(
		.clk_i(clk_i),
		.rstn_i(rstn_i),
		.serial_i(serial_i),
		.serial_o(serial)
	);
	// Trace: design.sv:30092:5
	pulp_clock_gating i_pulp_clock_gating(
		.clk_i(clk_i),
		.en_i(en_i),
		.test_en_i(1'b0),
		.clk_o(clk)
	);
	// Trace: design.sv:30099:5
	always @(posedge clk or negedge rstn_i)
		// Trace: design.sv:30100:9
		if (!rstn_i)
			// Trace: design.sv:30101:13
			serial_q <= 1'b0;
		else
			// Trace: design.sv:30103:13
			serial_q <= serial;
endmodule
module rrarbiter (
	clk_i,
	rst_ni,
	flush_i,
	en_i,
	req_i,
	ack_o,
	vld_o,
	idx_o
);
	// Trace: design.sv:30132:13
	parameter [31:0] NUM_REQ = 64;
	// Trace: design.sv:30133:13
	parameter [0:0] LOCK_IN = 1'b0;
	// Trace: design.sv:30135:3
	input wire clk_i;
	// Trace: design.sv:30136:3
	input wire rst_ni;
	// Trace: design.sv:30138:3
	input wire flush_i;
	// Trace: design.sv:30139:3
	input wire en_i;
	// Trace: design.sv:30140:3
	input wire [NUM_REQ - 1:0] req_i;
	// Trace: design.sv:30142:3
	output wire [NUM_REQ - 1:0] ack_o;
	// Trace: design.sv:30143:3
	output wire vld_o;
	// Trace: design.sv:30144:3
	output wire [$clog2(NUM_REQ) - 1:0] idx_o;
	// Trace: design.sv:30147:3
	wire req;
	// Trace: design.sv:30148:3
	assign vld_o = |req_i & en_i;
	// Trace: design.sv:30150:3
	localparam [31:0] sv2v_uu_i_rr_arb_tree_NumIn = NUM_REQ;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_IdxWidth = (sv2v_uu_i_rr_arb_tree_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_rr_arb_tree_NumIn)) : 32'd1);
	// removed localparam type sv2v_uu_i_rr_arb_tree_idx_t
	// removed localparam type sv2v_uu_i_rr_arb_tree_rr_i
	localparam [sv2v_uu_i_rr_arb_tree_IdxWidth - 1:0] sv2v_uu_i_rr_arb_tree_ext_rr_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_DataWidth = 1;
	// removed localparam type sv2v_uu_i_rr_arb_tree_DataType
	// removed localparam type sv2v_uu_i_rr_arb_tree_data_i
	localparam [(sv2v_uu_i_rr_arb_tree_NumIn * sv2v_uu_i_rr_arb_tree_DataWidth) - 1:0] sv2v_uu_i_rr_arb_tree_ext_data_i_0 = 1'sb0;
	rr_arb_tree #(
		.NumIn(NUM_REQ),
		.DataWidth(1),
		.LockIn(LOCK_IN)
	) i_rr_arb_tree(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_rr_arb_tree_ext_rr_i_0),
		.req_i(req_i),
		.gnt_o(ack_o),
		.data_i(sv2v_uu_i_rr_arb_tree_ext_data_i_0),
		.gnt_i(en_i & req),
		.req_o(req),
		.data_o(),
		.idx_o(idx_o)
	);
endmodule
module clock_divider (
	clk_i,
	rstn_i,
	test_mode_i,
	clk_gate_async_i,
	clk_div_data_i,
	clk_div_valid_i,
	clk_div_ack_o,
	clk_o
);
	reg _sv2v_0;
	// Trace: design.sv:30213:15
	parameter DIV_INIT = 0;
	// Trace: design.sv:30214:15
	parameter BYPASS_INIT = 1;
	// Trace: design.sv:30217:5
	input wire clk_i;
	// Trace: design.sv:30218:5
	input wire rstn_i;
	// Trace: design.sv:30219:5
	input wire test_mode_i;
	// Trace: design.sv:30220:5
	input wire clk_gate_async_i;
	// Trace: design.sv:30221:5
	input wire [7:0] clk_div_data_i;
	// Trace: design.sv:30222:5
	input wire clk_div_valid_i;
	// Trace: design.sv:30223:5
	output wire clk_div_ack_o;
	// Trace: design.sv:30224:5
	output wire clk_o;
	// Trace: design.sv:30227:4
	reg [1:0] state;
	reg [1:0] state_next;
	// Trace: design.sv:30229:4
	wire s_clk_out;
	// Trace: design.sv:30230:4
	reg s_clock_enable;
	// Trace: design.sv:30231:4
	wire s_clock_enable_gate;
	// Trace: design.sv:30232:4
	reg s_clk_div_valid;
	// Trace: design.sv:30234:4
	reg [7:0] reg_clk_div;
	// Trace: design.sv:30235:4
	wire s_clk_div_valid_sync;
	// Trace: design.sv:30237:4
	wire s_rstn_sync;
	// Trace: design.sv:30239:4
	reg [1:0] reg_ext_gate_sync;
	// Trace: design.sv:30241:5
	assign s_clock_enable_gate = s_clock_enable & reg_ext_gate_sync;
	// Trace: design.sv:30244:5
	rstgen i_rst_gen(
		.clk_i(clk_i),
		.rst_ni(rstn_i),
		.test_mode_i(test_mode_i),
		.rst_no(s_rstn_sync),
		.init_no()
	);
	// Trace: design.sv:30263:5
	pulp_sync_wedge i_edge_prop(
		.clk_i(clk_i),
		.rstn_i(s_rstn_sync),
		.en_i(1'b1),
		.serial_i(clk_div_valid_i),
		.serial_o(clk_div_ack_o),
		.r_edge_o(s_clk_div_valid_sync),
		.f_edge_o()
	);
	// Trace: design.sv:30274:5
	clock_divider_counter #(
		.BYPASS_INIT(BYPASS_INIT),
		.DIV_INIT(DIV_INIT)
	) i_clkdiv_cnt(
		.clk(clk_i),
		.rstn(s_rstn_sync),
		.test_mode(test_mode_i),
		.clk_div(reg_clk_div),
		.clk_div_valid(s_clk_div_valid),
		.clk_out(s_clk_out)
	);
	// Trace: design.sv:30289:5
	pulp_clock_gating i_clk_gate(
		.clk_i(s_clk_out),
		.en_i(s_clock_enable_gate),
		.test_en_i(test_mode_i),
		.clk_o(clk_o)
	);
	// Trace: design.sv:30297:5
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:30299:9
		case (state)
			2'd0: begin
				// Trace: design.sv:30302:13
				s_clock_enable = 1'b1;
				// Trace: design.sv:30303:13
				s_clk_div_valid = 1'b0;
				// Trace: design.sv:30304:13
				if (s_clk_div_valid_sync)
					// Trace: design.sv:30305:17
					state_next = 2'd1;
				else
					// Trace: design.sv:30307:17
					state_next = 2'd0;
			end
			2'd1: begin
				// Trace: design.sv:30312:13
				s_clock_enable = 1'b0;
				// Trace: design.sv:30313:13
				s_clk_div_valid = 1'b1;
				// Trace: design.sv:30314:13
				state_next = 2'd2;
			end
			2'd2: begin
				// Trace: design.sv:30319:13
				s_clock_enable = 1'b0;
				// Trace: design.sv:30320:13
				s_clk_div_valid = 1'b0;
				// Trace: design.sv:30321:13
				state_next = 2'd3;
			end
			2'd3: begin
				// Trace: design.sv:30326:13
				s_clock_enable = 1'b0;
				// Trace: design.sv:30327:13
				s_clk_div_valid = 1'b0;
				// Trace: design.sv:30328:13
				state_next = 2'd0;
			end
		endcase
	end
	// Trace: design.sv:30333:5
	always @(posedge clk_i or negedge s_rstn_sync)
		// Trace: design.sv:30335:9
		if (!s_rstn_sync)
			// Trace: design.sv:30336:13
			state <= 2'd0;
		else
			// Trace: design.sv:30338:13
			state <= state_next;
	// Trace: design.sv:30342:5
	always @(posedge clk_i or negedge s_rstn_sync)
		// Trace: design.sv:30344:9
		if (!s_rstn_sync)
			// Trace: design.sv:30345:13
			reg_clk_div <= 1'sb0;
		else if (s_clk_div_valid_sync)
			// Trace: design.sv:30347:19
			reg_clk_div <= clk_div_data_i;
	// Trace: design.sv:30351:5
	always @(posedge clk_i or negedge s_rstn_sync)
		// Trace: design.sv:30353:9
		if (!s_rstn_sync)
			// Trace: design.sv:30354:13
			reg_ext_gate_sync <= 2'b00;
		else
			// Trace: design.sv:30356:13
			reg_ext_gate_sync <= {clk_gate_async_i, reg_ext_gate_sync[1]};
	initial _sv2v_0 = 0;
endmodule
module fifo_v2_264A2 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	alm_full_o,
	alm_empty_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	// Trace: design.sv:30373:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:30374:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:30375:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:30376:15
	parameter [31:0] ALM_EMPTY_TH = 1;
	// Trace: design.sv:30377:15
	parameter [31:0] ALM_FULL_TH = 1;
	// Trace: design.sv:30378:20
	// removed localparam type dtype
	// Trace: design.sv:30380:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:30382:5
	input wire clk_i;
	// Trace: design.sv:30383:5
	input wire rst_ni;
	// Trace: design.sv:30384:5
	input wire flush_i;
	// Trace: design.sv:30385:5
	input wire testmode_i;
	// Trace: design.sv:30387:5
	output wire full_o;
	// Trace: design.sv:30388:5
	output wire empty_o;
	// Trace: design.sv:30389:5
	output wire alm_full_o;
	// Trace: design.sv:30390:5
	output wire alm_empty_o;
	// Trace: design.sv:30392:5
	input wire [31:0] data_i;
	// Trace: design.sv:30393:5
	input wire push_i;
	// Trace: design.sv:30395:5
	output wire [31:0] data_o;
	// Trace: design.sv:30396:5
	input wire pop_i;
	// Trace: design.sv:30399:5
	wire [ADDR_DEPTH - 1:0] usage;
	// Trace: design.sv:30402:5
	generate
		if (DEPTH == 0) begin : genblk1
			// Trace: design.sv:30403:9
			assign alm_full_o = 1'b0;
			// Trace: design.sv:30404:9
			assign alm_empty_o = 1'b0;
		end
		else begin : genblk1
			// Trace: design.sv:30406:9
			assign alm_full_o = usage >= ALM_FULL_TH[ADDR_DEPTH - 1:0];
			// Trace: design.sv:30407:9
			assign alm_empty_o = usage <= ALM_EMPTY_TH[ADDR_DEPTH - 1:0];
		end
	endgenerate
	// Trace: design.sv:30410:5
	fifo_v3_4D453 #(
		.FALL_THROUGH(FALL_THROUGH),
		.DATA_WIDTH(DATA_WIDTH),
		.DEPTH(DEPTH)
	) i_fifo_v3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.testmode_i(testmode_i),
		.full_o(full_o),
		.empty_o(empty_o),
		.usage_o(usage),
		.data_i(data_i),
		.push_i(push_i),
		.data_o(data_o),
		.pop_i(pop_i)
	);
endmodule
module fifo_v2_2D55D_D5824 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	alm_full_o,
	alm_empty_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	// removed localparam type dtype_DATA_WIDTH_type
	parameter [31:0] dtype_DATA_WIDTH = 0;
	// Trace: design.sv:30373:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:30374:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:30375:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:30376:15
	parameter [31:0] ALM_EMPTY_TH = 1;
	// Trace: design.sv:30377:15
	parameter [31:0] ALM_FULL_TH = 1;
	// Trace: design.sv:30378:20
	// removed localparam type dtype
	// Trace: design.sv:30380:15
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: design.sv:30382:5
	input wire clk_i;
	// Trace: design.sv:30383:5
	input wire rst_ni;
	// Trace: design.sv:30384:5
	input wire flush_i;
	// Trace: design.sv:30385:5
	input wire testmode_i;
	// Trace: design.sv:30387:5
	output wire full_o;
	// Trace: design.sv:30388:5
	output wire empty_o;
	// Trace: design.sv:30389:5
	output wire alm_full_o;
	// Trace: design.sv:30390:5
	output wire alm_empty_o;
	// Trace: design.sv:30392:5
	input wire [dtype_DATA_WIDTH - 1:0] data_i;
	// Trace: design.sv:30393:5
	input wire push_i;
	// Trace: design.sv:30395:5
	output wire [dtype_DATA_WIDTH - 1:0] data_o;
	// Trace: design.sv:30396:5
	input wire pop_i;
	// Trace: design.sv:30399:5
	wire [ADDR_DEPTH - 1:0] usage;
	// Trace: design.sv:30402:5
	generate
		if (DEPTH == 0) begin : genblk1
			// Trace: design.sv:30403:9
			assign alm_full_o = 1'b0;
			// Trace: design.sv:30404:9
			assign alm_empty_o = 1'b0;
		end
		else begin : genblk1
			// Trace: design.sv:30406:9
			assign alm_full_o = usage >= ALM_FULL_TH[ADDR_DEPTH - 1:0];
			// Trace: design.sv:30407:9
			assign alm_empty_o = usage <= ALM_EMPTY_TH[ADDR_DEPTH - 1:0];
		end
	endgenerate
	// Trace: design.sv:30410:5
	fifo_v3_19420_E888C #(
		.dtype_dtype_DATA_WIDTH(dtype_DATA_WIDTH),
		.FALL_THROUGH(FALL_THROUGH),
		.DATA_WIDTH(DATA_WIDTH),
		.DEPTH(DEPTH)
	) i_fifo_v3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.testmode_i(testmode_i),
		.full_o(full_o),
		.empty_o(empty_o),
		.usage_o(usage),
		.data_i(data_i),
		.push_i(push_i),
		.data_o(data_o),
		.pop_i(pop_i)
	);
endmodule
module fifo (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	threshold_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	// Trace: design.sv:30453:15
	parameter [0:0] FALL_THROUGH = 1'b0;
	// Trace: design.sv:30454:15
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:30455:15
	parameter [31:0] DEPTH = 8;
	// Trace: design.sv:30456:15
	parameter [31:0] THRESHOLD = 1;
	// Trace: design.sv:30457:20
	// removed localparam type dtype
	// Trace: design.sv:30459:5
	input wire clk_i;
	// Trace: design.sv:30460:5
	input wire rst_ni;
	// Trace: design.sv:30461:5
	input wire flush_i;
	// Trace: design.sv:30462:5
	input wire testmode_i;
	// Trace: design.sv:30464:5
	output wire full_o;
	// Trace: design.sv:30465:5
	output wire empty_o;
	// Trace: design.sv:30466:5
	output wire threshold_o;
	// Trace: design.sv:30468:5
	input wire [DATA_WIDTH - 1:0] data_i;
	// Trace: design.sv:30469:5
	input wire push_i;
	// Trace: design.sv:30471:5
	output wire [DATA_WIDTH - 1:0] data_o;
	// Trace: design.sv:30472:5
	input wire pop_i;
	// Trace: design.sv:30474:5
	fifo_v2_2D55D_D5824 #(
		.dtype_DATA_WIDTH(DATA_WIDTH),
		.FALL_THROUGH(FALL_THROUGH),
		.DATA_WIDTH(DATA_WIDTH),
		.DEPTH(DEPTH),
		.ALM_FULL_TH(THRESHOLD)
	) impl(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.testmode_i(testmode_i),
		.full_o(full_o),
		.empty_o(empty_o),
		.alm_full_o(threshold_o),
		.alm_empty_o(),
		.data_i(data_i),
		.push_i(push_i),
		.data_o(data_o),
		.pop_i(pop_i)
	);
endmodule
module edge_propagator_ack (
	clk_tx_i,
	rstn_tx_i,
	edge_i,
	ack_tx_o,
	clk_rx_i,
	rstn_rx_i,
	edge_o
);
	// Trace: design.sv:30509:3
	input wire clk_tx_i;
	// Trace: design.sv:30510:3
	input wire rstn_tx_i;
	// Trace: design.sv:30511:3
	input wire edge_i;
	// Trace: design.sv:30512:3
	output wire ack_tx_o;
	// Trace: design.sv:30513:3
	input wire clk_rx_i;
	// Trace: design.sv:30514:3
	input wire rstn_rx_i;
	// Trace: design.sv:30515:3
	output wire edge_o;
	// Trace: design.sv:30518:3
	reg [1:0] sync_a;
	// Trace: design.sv:30519:3
	wire sync_b;
	// Trace: design.sv:30521:3
	reg r_input_reg;
	// Trace: design.sv:30522:3
	wire s_input_reg_next;
	// Trace: design.sv:30524:3
	assign ack_tx_o = sync_a[0];
	// Trace: design.sv:30526:3
	assign s_input_reg_next = edge_i | (r_input_reg & ~sync_a[0]);
	// Trace: design.sv:30528:3
	always @(negedge rstn_tx_i or posedge clk_tx_i)
		// Trace: design.sv:30529:5
		if (~rstn_tx_i) begin
			// Trace: design.sv:30530:7
			r_input_reg <= 1'b0;
			// Trace: design.sv:30531:7
			sync_a <= 2'b00;
		end
		else begin
			// Trace: design.sv:30533:7
			r_input_reg <= s_input_reg_next;
			// Trace: design.sv:30534:7
			sync_a <= {sync_b, sync_a[1]};
		end
	// Trace: design.sv:30538:3
	pulp_sync_wedge u_sync_clkb(
		.clk_i(clk_rx_i),
		.rstn_i(rstn_rx_i),
		.en_i(1'b1),
		.serial_i(r_input_reg),
		.r_edge_o(edge_o),
		.f_edge_o(),
		.serial_o(sync_b)
	);
endmodule
module edge_propagator (
	clk_tx_i,
	rstn_tx_i,
	edge_i,
	clk_rx_i,
	rstn_rx_i,
	edge_o
);
	// Trace: design.sv:30562:3
	input wire clk_tx_i;
	// Trace: design.sv:30563:3
	input wire rstn_tx_i;
	// Trace: design.sv:30564:3
	input wire edge_i;
	// Trace: design.sv:30565:3
	input wire clk_rx_i;
	// Trace: design.sv:30566:3
	input wire rstn_rx_i;
	// Trace: design.sv:30567:3
	output wire edge_o;
	// Trace: design.sv:30570:3
	edge_propagator_ack i_edge_propagator_ack(
		.clk_tx_i(clk_tx_i),
		.rstn_tx_i(rstn_tx_i),
		.edge_i(edge_i),
		.ack_tx_o(),
		.clk_rx_i(clk_rx_i),
		.rstn_rx_i(rstn_rx_i),
		.edge_o(edge_o)
	);
endmodule
module edge_propagator_rx (
	clk_i,
	rstn_i,
	valid_i,
	ack_o,
	valid_o
);
	// Trace: design.sv:30594:5
	input wire clk_i;
	// Trace: design.sv:30595:5
	input wire rstn_i;
	// Trace: design.sv:30596:5
	input wire valid_i;
	// Trace: design.sv:30597:5
	output wire ack_o;
	// Trace: design.sv:30598:5
	output wire valid_o;
	// Trace: design.sv:30601:5
	pulp_sync_wedge i_sync_clkb(
		.clk_i(clk_i),
		.rstn_i(rstn_i),
		.en_i(1'b1),
		.serial_i(valid_i),
		.r_edge_o(valid_o),
		.f_edge_o(),
		.serial_o(ack_o)
	);
endmodule
// removed interface: REG_BUS
module periph_to_reg_35129 (
	clk_i,
	rst_ni,
	req_i,
	add_i,
	wen_i,
	wdata_i,
	be_i,
	id_i,
	gnt_o,
	r_rdata_o,
	r_opc_o,
	r_id_o,
	r_valid_o,
	reg_req_o,
	reg_rsp_i
);
	reg _sv2v_0;
	// Trace: design.sv:30668:13
	parameter [31:0] AW = 32;
	// Trace: design.sv:30669:13
	parameter [31:0] DW = 32;
	// Trace: design.sv:30670:13
	parameter [31:0] BW = 8;
	// Trace: design.sv:30671:13
	parameter [31:0] IW = 0;
	// Trace: design.sv:30672:26
	// removed localparam type req_t
	// Trace: design.sv:30673:26
	// removed localparam type rsp_t
	// Trace: design.sv:30675:3
	input wire clk_i;
	// Trace: design.sv:30676:3
	input wire rst_ni;
	// Trace: design.sv:30678:3
	input wire req_i;
	// Trace: design.sv:30679:3
	input wire [AW - 1:0] add_i;
	// Trace: design.sv:30680:3
	input wire wen_i;
	// Trace: design.sv:30681:3
	input wire [DW - 1:0] wdata_i;
	// Trace: design.sv:30682:3
	input wire [(DW / BW) - 1:0] be_i;
	// Trace: design.sv:30683:3
	input wire [IW - 1:0] id_i;
	// Trace: design.sv:30684:3
	output wire gnt_o;
	// Trace: design.sv:30685:3
	output wire [DW - 1:0] r_rdata_o;
	// Trace: design.sv:30686:3
	output wire r_opc_o;
	// Trace: design.sv:30687:3
	output wire [IW - 1:0] r_id_o;
	// Trace: design.sv:30688:3
	output wire r_valid_o;
	// Trace: design.sv:30690:3
	output wire [69:0] reg_req_o;
	// Trace: design.sv:30691:3
	input wire [33:0] reg_rsp_i;
	// Trace: design.sv:30694:3
	reg [IW - 1:0] r_id_d;
	reg [IW - 1:0] r_id_q;
	// Trace: design.sv:30695:3
	reg r_opc_d;
	reg r_opc_q;
	// Trace: design.sv:30696:3
	reg r_valid_d;
	reg r_valid_q;
	// Trace: design.sv:30697:3
	reg [DW - 1:0] r_rdata_d;
	reg [DW - 1:0] r_rdata_q;
	// Trace: design.sv:30699:3
	always @(*) begin : proc_logic
		if (_sv2v_0)
			;
		// Trace: design.sv:30700:5
		r_id_d = id_i;
		// Trace: design.sv:30701:5
		r_opc_d = reg_rsp_i[33];
		// Trace: design.sv:30702:5
		r_valid_d = gnt_o;
		// Trace: design.sv:30703:5
		r_rdata_d = reg_rsp_i[31-:32];
	end
	// Trace: design.sv:30706:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_seq
		// Trace: design.sv:30707:5
		if (!rst_ni) begin
			// Trace: design.sv:30708:7
			r_id_q <= 1'sb0;
			// Trace: design.sv:30709:7
			r_opc_q <= 1'sb0;
			// Trace: design.sv:30710:7
			r_valid_q <= 1'sb0;
			// Trace: design.sv:30711:7
			r_rdata_q <= 1'sb0;
		end
		else begin
			// Trace: design.sv:30713:7
			r_id_q <= r_id_d;
			// Trace: design.sv:30714:7
			r_opc_q <= r_opc_d;
			// Trace: design.sv:30715:7
			r_valid_q <= r_valid_d;
			// Trace: design.sv:30716:7
			r_rdata_q <= r_rdata_d;
		end
	end
	// Trace: design.sv:30720:3
	assign reg_req_o[63-:32] = add_i;
	// Trace: design.sv:30721:3
	assign reg_req_o[68] = ~wen_i;
	// Trace: design.sv:30722:3
	assign reg_req_o[31-:32] = wdata_i;
	// Trace: design.sv:30723:3
	assign reg_req_o[67-:4] = be_i;
	// Trace: design.sv:30724:3
	assign reg_req_o[69] = req_i;
	// Trace: design.sv:30726:3
	assign gnt_o = req_i & reg_rsp_i[32];
	// Trace: design.sv:30728:3
	assign r_rdata_o = r_rdata_q;
	// Trace: design.sv:30729:3
	assign r_opc_o = r_opc_q;
	// Trace: design.sv:30730:3
	assign r_id_o = r_id_q;
	// Trace: design.sv:30731:3
	assign r_valid_o = r_valid_q;
	initial _sv2v_0 = 0;
endmodule
module reg_demux_64ED6 (
	clk_i,
	rst_ni,
	in_select_i,
	in_req_i,
	in_rsp_o,
	out_req_o,
	out_rsp_i
);
	reg _sv2v_0;
	// Trace: design.sv:30773:13
	parameter [31:0] NoPorts = 32'd0;
	// Trace: design.sv:30774:18
	// removed localparam type req_t
	// Trace: design.sv:30775:18
	// removed localparam type rsp_t
	// Trace: design.sv:30777:13
	parameter [31:0] SelectWidth = (NoPorts > 32'd1 ? $clog2(NoPorts) : 32'd1);
	// Trace: design.sv:30778:26
	// removed localparam type select_t
	// Trace: design.sv:30780:3
	input wire clk_i;
	// Trace: design.sv:30781:3
	input wire rst_ni;
	// Trace: design.sv:30782:3
	input wire [SelectWidth - 1:0] in_select_i;
	// Trace: design.sv:30783:3
	input wire [69:0] in_req_i;
	// Trace: design.sv:30784:3
	output reg [33:0] in_rsp_o;
	// Trace: design.sv:30785:3
	output reg [(NoPorts * 70) - 1:0] out_req_o;
	// Trace: design.sv:30786:3
	input wire [(NoPorts * 34) - 1:0] out_rsp_i;
	// Trace: design.sv:30789:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:30790:5
		out_req_o = 1'sb0;
		// Trace: design.sv:30791:5
		in_rsp_o = 1'sb0;
		// Trace: design.sv:30792:5
		out_req_o[in_select_i * 70+:70] = in_req_i;
		// Trace: design.sv:30793:5
		in_rsp_o = out_rsp_i[in_select_i * 34+:34];
	end
	initial _sv2v_0 = 0;
endmodule
module reg_to_tlul_223C2_EF763 (
	tl_o,
	tl_i,
	reg_req_i,
	reg_rsp_o
);
	// removed localparam type tl_a_user_t_tlul_pkg_DataIntgWidth_type
	// removed localparam type tl_a_user_t_tlul_pkg_H2DCmdIntgWidth_type
	parameter signed [31:0] tl_a_user_t_tlul_pkg_DataIntgWidth = 0;
	parameter signed [31:0] tl_a_user_t_tlul_pkg_H2DCmdIntgWidth = 0;
	// removed localparam type tl_d2h_t_tlul_pkg_D2HRspIntgWidth_type
	// removed localparam type tl_d2h_t_tlul_pkg_DataIntgWidth_type
	// removed localparam type tl_d2h_t_top_pkg_TL_AIW_type
	// removed localparam type tl_d2h_t_top_pkg_TL_DIW_type
	// removed localparam type tl_d2h_t_top_pkg_TL_DW_type
	// removed localparam type tl_d2h_t_top_pkg_TL_SZW_type
	parameter signed [31:0] tl_d2h_t_tlul_pkg_D2HRspIntgWidth = 0;
	parameter signed [31:0] tl_d2h_t_tlul_pkg_DataIntgWidth = 0;
	parameter signed [31:0] tl_d2h_t_top_pkg_TL_AIW = 0;
	parameter signed [31:0] tl_d2h_t_top_pkg_TL_DIW = 0;
	parameter signed [31:0] tl_d2h_t_top_pkg_TL_DW = 0;
	parameter signed [31:0] tl_d2h_t_top_pkg_TL_SZW = 0;
	// removed localparam type tl_h2d_t_tlul_pkg_DataIntgWidth_type
	// removed localparam type tl_h2d_t_tlul_pkg_H2DCmdIntgWidth_type
	// removed localparam type tl_h2d_t_top_pkg_TL_AIW_type
	// removed localparam type tl_h2d_t_top_pkg_TL_AW_type
	// removed localparam type tl_h2d_t_top_pkg_TL_DBW_type
	// removed localparam type tl_h2d_t_top_pkg_TL_DW_type
	// removed localparam type tl_h2d_t_top_pkg_TL_SZW_type
	parameter signed [31:0] tl_h2d_t_tlul_pkg_DataIntgWidth = 0;
	parameter signed [31:0] tl_h2d_t_tlul_pkg_H2DCmdIntgWidth = 0;
	parameter signed [31:0] tl_h2d_t_top_pkg_TL_AIW = 0;
	parameter signed [31:0] tl_h2d_t_top_pkg_TL_AW = 0;
	parameter signed [31:0] tl_h2d_t_top_pkg_TL_DBW = 0;
	parameter signed [31:0] tl_h2d_t_top_pkg_TL_DW = 0;
	parameter signed [31:0] tl_h2d_t_top_pkg_TL_SZW = 0;
	// Trace: design.sv:30806:18
	// removed localparam type req_t
	// Trace: design.sv:30807:18
	// removed localparam type rsp_t
	// Trace: design.sv:30808:18
	// removed localparam type tl_h2d_t
	// Trace: design.sv:30809:18
	// removed localparam type tl_d2h_t
	// Trace: design.sv:30811:18
	// removed localparam type tl_a_user_t
	// Trace: design.sv:30812:18
	// removed localparam type tl_a_op_e
	// Trace: design.sv:30813:13
	parameter [((7 + tl_a_user_t_tlul_pkg_H2DCmdIntgWidth) + tl_a_user_t_tlul_pkg_DataIntgWidth) - 1:0] TL_A_USER_DEFAULT = 1'sb0;
	// Trace: design.sv:30814:13
	parameter [2:0] PutFullData = 1'sb0;
	// Trace: design.sv:30815:13
	parameter [2:0] Get = 1'sb0;
	// Trace: design.sv:30818:5
	output wire [((((((7 + tl_h2d_t_top_pkg_TL_SZW) + tl_h2d_t_top_pkg_TL_AIW) + tl_h2d_t_top_pkg_TL_AW) + tl_h2d_t_top_pkg_TL_DBW) + tl_h2d_t_top_pkg_TL_DW) + ((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth)) + 0:0] tl_o;
	// Trace: design.sv:30819:5
	input wire [(((((7 + tl_d2h_t_top_pkg_TL_SZW) + tl_d2h_t_top_pkg_TL_AIW) + tl_d2h_t_top_pkg_TL_DIW) + tl_d2h_t_top_pkg_TL_DW) + (tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth)) + 1:0] tl_i;
	// Trace: design.sv:30822:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:30823:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:30827:3
	assign tl_o[7 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))))] = reg_req_i[69] & tl_i[0];
	// Trace: design.sv:30828:3
	assign tl_o[6 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))))-:((6 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))))) >= (3 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))))))) ? ((6 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))))) - (3 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)))))))) + 1 : ((3 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))))))) - (6 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))))))) + 1)] = (reg_req_i[68] ? PutFullData : Get);
	// Trace: design.sv:30829:3
	assign tl_o[3 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))))-:((3 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))))) >= (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)))))) ? ((3 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))))) - (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))))))) + 1 : ((tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))))))) + 1)] = 1'sb0;
	// Trace: design.sv:30830:3
	assign tl_o[tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))))-:((tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))))) >= (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))))) ? ((tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))))) - (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)))))) + 1 : ((tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))))) - (tl_h2d_t_top_pkg_TL_SZW + (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))))) + 1)] = 'h2;
	// Trace: design.sv:30831:3
	assign tl_o[tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))-:((tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))) >= (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)))) ? ((tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))) - (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))))) + 1 : ((tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)))) - (tl_h2d_t_top_pkg_TL_AIW + (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))))) + 1)] = 1'sb0;
	// Trace: design.sv:30832:3
	assign tl_o[tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))-:((tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))) >= (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))) ? ((tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))) - (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)))) + 1 : ((tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))) - (tl_h2d_t_top_pkg_TL_AW + (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))))) + 1)] = reg_req_i[63-:32];
	// Trace: design.sv:30833:3
	assign tl_o[tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))-:((tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))) >= (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)) ? ((tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))) - (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1))) + 1 : ((tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)) - (tl_h2d_t_top_pkg_TL_DBW + (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)))) + 1)] = reg_req_i[67-:4];
	// Trace: design.sv:30834:3
	assign tl_o[tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)-:((tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)) >= (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1) ? ((tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0)) - (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1)) + 1 : ((((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 1) - (tl_h2d_t_top_pkg_TL_DW + (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))) + 1)] = reg_req_i[31-:32];
	// Trace: design.sv:30835:3
	assign tl_o[((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0-:((((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0) >= 1 ? ((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0 : 2 - (((7 + tl_h2d_t_tlul_pkg_H2DCmdIntgWidth) + tl_h2d_t_tlul_pkg_DataIntgWidth) + 0))] = TL_A_USER_DEFAULT;
	// Trace: design.sv:30836:3
	assign tl_o[0] = 1'b1;
	// Trace: design.sv:30838:3
	assign reg_rsp_o[32] = tl_i[7 + (tl_d2h_t_top_pkg_TL_SZW + (tl_d2h_t_top_pkg_TL_AIW + (tl_d2h_t_top_pkg_TL_DIW + (tl_d2h_t_top_pkg_TL_DW + ((tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth) + 1)))))] & tl_o[0];
	// Trace: design.sv:30839:3
	assign reg_rsp_o[31-:32] = tl_i[tl_d2h_t_top_pkg_TL_DW + ((tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth) + 1)-:((tl_d2h_t_top_pkg_TL_DW + ((tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth) + 1)) >= ((tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth) + 2) ? ((tl_d2h_t_top_pkg_TL_DW + ((tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth) + 1)) - ((tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth) + 2) - (tl_d2h_t_top_pkg_TL_DW + ((tl_d2h_t_tlul_pkg_D2HRspIntgWidth + tl_d2h_t_tlul_pkg_DataIntgWidth) + 1))) + 1)];
	// Trace: design.sv:30840:3
	assign reg_rsp_o[33] = tl_i[1];
endmodule
// removed package "dm"
// removed package "addr_map_rule_pkg"
// removed package "obi_pkg"
// removed package "reg_pkg"
// removed package "core_v_mini_mcu_pkg"
// removed package "power_manager_reg_pkg"
module rv_plic_gateway (
	clk_i,
	rst_ni,
	src_i,
	le_i,
	claim_i,
	complete_i,
	ip_o
);
	reg _sv2v_0;
	// Trace: design.sv:32127:13
	parameter signed [31:0] N_SOURCE = 32;
	// Trace: design.sv:32129:3
	input clk_i;
	// Trace: design.sv:32130:3
	input rst_ni;
	// Trace: design.sv:32132:3
	input [N_SOURCE - 1:0] src_i;
	// Trace: design.sv:32133:3
	input [N_SOURCE - 1:0] le_i;
	// Trace: design.sv:32135:3
	input [N_SOURCE - 1:0] claim_i;
	// Trace: design.sv:32136:3
	input [N_SOURCE - 1:0] complete_i;
	// Trace: design.sv:32138:3
	output reg [N_SOURCE - 1:0] ip_o;
	// Trace: design.sv:32141:3
	reg [N_SOURCE - 1:0] ia;
	// Trace: design.sv:32143:3
	reg [N_SOURCE - 1:0] set;
	// Trace: design.sv:32144:3
	reg [N_SOURCE - 1:0] src_q;
	// Trace: design.sv:32146:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:32147:5
		if (!rst_ni)
			// Trace: design.sv:32147:18
			src_q <= 1'sb0;
		else
			// Trace: design.sv:32148:18
			src_q <= src_i;
	// Trace: design.sv:32151:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:32152:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:32152:10
			reg signed [31:0] i;
			// Trace: design.sv:32152:10
			for (i = 0; i < N_SOURCE; i = i + 1)
				begin
					// Trace: design.sv:32153:7
					set[i] = (le_i[i] ? src_i[i] & ~src_q[i] : src_i[i]);
				end
		end
	end
	// Trace: design.sv:32161:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:32162:5
		if (!rst_ni)
			// Trace: design.sv:32163:7
			ip_o <= 1'sb0;
		else
			// Trace: design.sv:32165:7
			ip_o <= (ip_o | ((set & ~ia) & ~ip_o)) & ~(ip_o & claim_i);
	// Trace: design.sv:32173:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:32174:5
		if (!rst_ni)
			// Trace: design.sv:32175:7
			ia <= 1'sb0;
		else
			// Trace: design.sv:32177:7
			ia <= (ia | (set & ~ia)) & ~((ia & complete_i) & ~ip_o);
	initial _sv2v_0 = 0;
endmodule
module rv_plic_target (
	clk_i,
	rst_ni,
	ip_i,
	ie_i,
	prio_i,
	threshold_i,
	irq_o,
	irq_id_o
);
	// Trace: design.sv:32199:13
	parameter signed [31:0] N_SOURCE = 32;
	// Trace: design.sv:32200:13
	parameter signed [31:0] MAX_PRIO = 7;
	// Trace: design.sv:32203:14
	localparam signed [31:0] SrcWidth = 6;
	// Trace: design.sv:32204:14
	localparam signed [31:0] PrioWidth = $clog2(MAX_PRIO + 1);
	// Trace: design.sv:32206:3
	input clk_i;
	// Trace: design.sv:32207:3
	input rst_ni;
	// Trace: design.sv:32209:3
	input [N_SOURCE - 1:0] ip_i;
	// Trace: design.sv:32210:3
	input [N_SOURCE - 1:0] ie_i;
	// Trace: design.sv:32212:3
	input [(N_SOURCE * PrioWidth) - 1:0] prio_i;
	// Trace: design.sv:32213:3
	input [PrioWidth - 1:0] threshold_i;
	// Trace: design.sv:32215:3
	output wire irq_o;
	// Trace: design.sv:32216:3
	output wire [5:0] irq_id_o;
	// Trace: design.sv:32224:3
	localparam signed [31:0] NumLevels = $clog2(N_SOURCE);
	// Trace: design.sv:32225:3
	wire [(2 ** (NumLevels + 1)) - 2:0] is_tree;
	// Trace: design.sv:32226:3
	wire [(((2 ** (NumLevels + 1)) - 2) >= 0 ? (((2 ** (NumLevels + 1)) - 1) * SrcWidth) - 1 : ((3 - (2 ** (NumLevels + 1))) * SrcWidth) + ((((2 ** (NumLevels + 1)) - 2) * SrcWidth) - 1)):(((2 ** (NumLevels + 1)) - 2) >= 0 ? 0 : ((2 ** (NumLevels + 1)) - 2) * SrcWidth)] id_tree;
	// Trace: design.sv:32227:3
	wire [(((2 ** (NumLevels + 1)) - 2) >= 0 ? (((2 ** (NumLevels + 1)) - 1) * PrioWidth) - 1 : ((3 - (2 ** (NumLevels + 1))) * PrioWidth) + ((((2 ** (NumLevels + 1)) - 2) * PrioWidth) - 1)):(((2 ** (NumLevels + 1)) - 2) >= 0 ? 0 : ((2 ** (NumLevels + 1)) - 2) * PrioWidth)] max_tree;
	// Trace: design.sv:32229:3
	genvar _gv_level_5;
	generate
		for (_gv_level_5 = 0; _gv_level_5 < (NumLevels + 1); _gv_level_5 = _gv_level_5 + 1) begin : gen_tree
			localparam level = _gv_level_5;
			// Trace: design.sv:32241:5
			localparam signed [31:0] Base0 = (2 ** level) - 1;
			// Trace: design.sv:32242:5
			localparam signed [31:0] Base1 = (2 ** (level + 1)) - 1;
			genvar _gv_offset_1;
			for (_gv_offset_1 = 0; _gv_offset_1 < (2 ** level); _gv_offset_1 = _gv_offset_1 + 1) begin : gen_level
				localparam offset = _gv_offset_1;
				// Trace: design.sv:32245:7
				localparam signed [31:0] Pa = Base0 + offset;
				// Trace: design.sv:32246:7
				localparam signed [31:0] C0 = Base1 + (2 * offset);
				// Trace: design.sv:32247:7
				localparam signed [31:0] C1 = (Base1 + (2 * offset)) + 1;
				if (level == NumLevels) begin : gen_leafs
					if (offset < N_SOURCE) begin : gen_assign
						// Trace: design.sv:32253:11
						assign is_tree[Pa] = ip_i[offset] & ie_i[offset];
						// Trace: design.sv:32254:11
						assign id_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? Pa : ((2 ** (NumLevels + 1)) - 2) - Pa) * SrcWidth+:SrcWidth] = offset;
						// Trace: design.sv:32255:11
						assign max_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? Pa : ((2 ** (NumLevels + 1)) - 2) - Pa) * PrioWidth+:PrioWidth] = prio_i[((N_SOURCE - 1) - offset) * PrioWidth+:PrioWidth];
					end
					else begin : gen_tie_off
						// Trace: design.sv:32257:11
						assign is_tree[Pa] = 1'sb0;
						// Trace: design.sv:32258:11
						assign id_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? Pa : ((2 ** (NumLevels + 1)) - 2) - Pa) * SrcWidth+:SrcWidth] = 1'sb0;
						// Trace: design.sv:32259:11
						assign max_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? Pa : ((2 ** (NumLevels + 1)) - 2) - Pa) * PrioWidth+:PrioWidth] = 1'sb0;
					end
				end
				else begin : gen_nodes
					// Trace: design.sv:32277:9
					wire sel;
					// Trace: design.sv:32280:9
					assign sel = (~is_tree[C0] & is_tree[C1]) | ((is_tree[C0] & is_tree[C1]) & (max_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? C1 : ((2 ** (NumLevels + 1)) - 2) - C1) * PrioWidth+:PrioWidth] > max_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? C0 : ((2 ** (NumLevels + 1)) - 2) - C0) * PrioWidth+:PrioWidth]));
					// Trace: design.sv:32283:9
					assign is_tree[Pa] = (sel & is_tree[C1]) | (~sel & is_tree[C0]);
					// Trace: design.sv:32285:9
					assign id_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? Pa : ((2 ** (NumLevels + 1)) - 2) - Pa) * SrcWidth+:SrcWidth] = ({SrcWidth {sel}} & id_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? C1 : ((2 ** (NumLevels + 1)) - 2) - C1) * SrcWidth+:SrcWidth]) | ({SrcWidth {~sel}} & id_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? C0 : ((2 ** (NumLevels + 1)) - 2) - C0) * SrcWidth+:SrcWidth]);
					// Trace: design.sv:32287:9
					assign max_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? Pa : ((2 ** (NumLevels + 1)) - 2) - Pa) * PrioWidth+:PrioWidth] = ({PrioWidth {sel}} & max_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? C1 : ((2 ** (NumLevels + 1)) - 2) - C1) * PrioWidth+:PrioWidth]) | ({PrioWidth {~sel}} & max_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? C0 : ((2 ** (NumLevels + 1)) - 2) - C0) * PrioWidth+:PrioWidth]);
				end
			end
		end
	endgenerate
	// Trace: design.sv:32293:3
	wire irq_d;
	reg irq_q;
	// Trace: design.sv:32294:3
	wire [5:0] irq_id_d;
	reg [5:0] irq_id_q;
	// Trace: design.sv:32297:3
	assign irq_d = (max_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? 0 : (2 ** (NumLevels + 1)) - 2) * PrioWidth+:PrioWidth] > threshold_i ? is_tree[0] : 1'b0);
	// Trace: design.sv:32298:3
	assign irq_id_d = (is_tree[0] ? id_tree[(((2 ** (NumLevels + 1)) - 2) >= 0 ? 0 : (2 ** (NumLevels + 1)) - 2) * SrcWidth+:SrcWidth] : {6 {1'sb0}});
	// Trace: design.sv:32300:3
	always @(posedge clk_i or negedge rst_ni) begin : gen_regs
		// Trace: design.sv:32301:5
		if (!rst_ni) begin
			// Trace: design.sv:32302:7
			irq_q <= 1'b0;
			// Trace: design.sv:32303:7
			irq_id_q <= 1'sb0;
		end
		else begin
			// Trace: design.sv:32305:7
			irq_q <= irq_d;
			// Trace: design.sv:32306:7
			irq_id_q <= irq_id_d;
		end
	end
	// Trace: design.sv:32310:3
	assign irq_o = irq_q;
	// Trace: design.sv:32311:3
	assign irq_id_o = irq_id_q;
endmodule
module prim_arbiter_ppc (
	clk_i,
	rst_ni,
	req_i,
	data_i,
	gnt_o,
	idx_o,
	valid_o,
	data_o,
	ready_i
);
	reg _sv2v_0;
	// Trace: design.sv:32343:13
	parameter [31:0] N = 8;
	// Trace: design.sv:32344:13
	parameter [31:0] DW = 32;
	// Trace: design.sv:32348:13
	parameter [0:0] EnDataPort = 1;
	// Trace: design.sv:32351:13
	parameter [0:0] EnReqStabA = 1;
	// Trace: design.sv:32354:14
	localparam signed [31:0] IdxW = $clog2(N);
	// Trace: design.sv:32356:3
	input clk_i;
	// Trace: design.sv:32357:3
	input rst_ni;
	// Trace: design.sv:32359:3
	input [N - 1:0] req_i;
	// Trace: design.sv:32360:3
	input [(N * DW) - 1:0] data_i;
	// Trace: design.sv:32361:3
	output wire [N - 1:0] gnt_o;
	// Trace: design.sv:32362:3
	output reg [IdxW - 1:0] idx_o;
	// Trace: design.sv:32364:3
	output wire valid_o;
	// Trace: design.sv:32365:3
	output reg [DW - 1:0] data_o;
	// Trace: design.sv:32366:3
	input ready_i;
	// Trace: design.sv:32372:3
	generate
		if (N == 1) begin : gen_degenerate_case
			// Trace: design.sv:32374:5
			assign valid_o = req_i[0];
			// Trace: design.sv:32375:5
			wire [DW:1] sv2v_tmp_9E8F4;
			assign sv2v_tmp_9E8F4 = data_i[(N - 1) * DW+:DW];
			always @(*) data_o = sv2v_tmp_9E8F4;
			// Trace: design.sv:32376:5
			assign gnt_o[0] = valid_o & ready_i;
			// Trace: design.sv:32377:5
			wire [IdxW:1] sv2v_tmp_8C7A7;
			assign sv2v_tmp_8C7A7 = 1'sb0;
			always @(*) idx_o = sv2v_tmp_8C7A7;
		end
		else begin : gen_normal_case
			// Trace: design.sv:32381:5
			wire [N - 1:0] masked_req;
			// Trace: design.sv:32382:5
			reg [N - 1:0] ppc_out;
			// Trace: design.sv:32383:5
			wire [N - 1:0] arb_req;
			// Trace: design.sv:32384:5
			reg [N - 1:0] mask;
			wire [N - 1:0] mask_next;
			// Trace: design.sv:32385:5
			wire [N - 1:0] winner;
			// Trace: design.sv:32387:5
			assign masked_req = mask & req_i;
			// Trace: design.sv:32388:5
			assign arb_req = (|masked_req ? masked_req : req_i);
			// Trace: design.sv:32393:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:32394:7
				ppc_out[0] = arb_req[0];
				// Trace: design.sv:32395:7
				begin : sv2v_autoblock_1
					// Trace: design.sv:32395:12
					reg signed [31:0] i;
					// Trace: design.sv:32395:12
					for (i = 1; i < N; i = i + 1)
						begin
							// Trace: design.sv:32396:9
							ppc_out[i] = ppc_out[i - 1] | arb_req[i];
						end
				end
			end
			// Trace: design.sv:32401:5
			assign winner = ppc_out ^ {ppc_out[N - 2:0], 1'b0};
			// Trace: design.sv:32402:5
			assign gnt_o = (ready_i ? winner : {N {1'sb0}});
			// Trace: design.sv:32404:5
			assign valid_o = |req_i;
			// Trace: design.sv:32406:5
			assign mask_next = {ppc_out[N - 2:0], 1'b0};
			// Trace: design.sv:32407:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:32408:7
				if (!rst_ni)
					// Trace: design.sv:32409:9
					mask <= 1'sb0;
				else if (valid_o && ready_i)
					// Trace: design.sv:32412:9
					mask <= mask_next;
				else if (valid_o && !ready_i)
					// Trace: design.sv:32415:9
					mask <= ppc_out;
			if (EnDataPort == 1) begin : gen_datapath
				// Trace: design.sv:32420:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:32421:9
					data_o = 1'sb0;
					// Trace: design.sv:32422:9
					begin : sv2v_autoblock_2
						// Trace: design.sv:32422:14
						reg signed [31:0] i;
						// Trace: design.sv:32422:14
						for (i = 0; i < N; i = i + 1)
							begin
								// Trace: design.sv:32423:11
								if (winner[i])
									// Trace: design.sv:32424:13
									data_o = data_i[((N - 1) - i) * DW+:DW];
							end
					end
				end
			end
			else begin : gen_nodatapath
				// Trace: design.sv:32429:7
				wire [DW:1] sv2v_tmp_116D0;
				assign sv2v_tmp_116D0 = 1'sb1;
				always @(*) data_o = sv2v_tmp_116D0;
				// Trace: design.sv:32431:7
				wire [(N * DW) - 1:0] unused_data;
				// Trace: design.sv:32432:7
				assign unused_data = data_i;
			end
			// Trace: design.sv:32435:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:32436:7
				idx_o = 1'sb0;
				// Trace: design.sv:32437:7
				begin : sv2v_autoblock_3
					// Trace: design.sv:32437:12
					reg [31:0] i;
					// Trace: design.sv:32437:12
					for (i = 0; i < N; i = i + 1)
						begin
							// Trace: design.sv:32438:9
							if (winner[i])
								// Trace: design.sv:32439:11
								idx_o = i[IdxW - 1:0];
						end
				end
			end
		end
	endgenerate
	// Trace: design.sv:32477:1
	// Trace: design.sv:32482:1
	initial _sv2v_0 = 0;
endmodule
module prim_arbiter_tree (
	clk_i,
	rst_ni,
	req_i,
	data_i,
	gnt_o,
	idx_o,
	valid_o,
	data_o,
	ready_i
);
	reg _sv2v_0;
	// Trace: design.sv:32576:13
	parameter signed [31:0] N = 8;
	// Trace: design.sv:32577:13
	parameter signed [31:0] DW = 32;
	// Trace: design.sv:32581:13
	parameter [0:0] EnDataPort = 1;
	// Trace: design.sv:32584:13
	parameter [0:0] EnReqStabA = 1;
	// Trace: design.sv:32587:14
	localparam signed [31:0] IdxW = $clog2(N);
	// Trace: design.sv:32589:3
	input clk_i;
	// Trace: design.sv:32590:3
	input rst_ni;
	// Trace: design.sv:32592:3
	input [N - 1:0] req_i;
	// Trace: design.sv:32593:3
	input [(N * DW) - 1:0] data_i;
	// Trace: design.sv:32594:3
	output wire [N - 1:0] gnt_o;
	// Trace: design.sv:32595:3
	output wire [IdxW - 1:0] idx_o;
	// Trace: design.sv:32597:3
	output wire valid_o;
	// Trace: design.sv:32598:3
	output wire [DW - 1:0] data_o;
	// Trace: design.sv:32599:3
	input ready_i;
	// Trace: design.sv:32605:3
	generate
		if (N == 1) begin : gen_degenerate_case
			// Trace: design.sv:32607:5
			assign valid_o = req_i[0];
			// Trace: design.sv:32608:5
			assign data_o = data_i[(N - 1) * DW+:DW];
			// Trace: design.sv:32609:5
			assign gnt_o[0] = valid_o & ready_i;
			// Trace: design.sv:32610:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_normal_case
			// Trace: design.sv:32616:5
			reg [(2 ** (IdxW + 1)) - 2:0] req_tree;
			// Trace: design.sv:32617:5
			reg [(2 ** (IdxW + 1)) - 2:0] prio_tree;
			// Trace: design.sv:32618:5
			reg [(2 ** (IdxW + 1)) - 2:0] sel_tree;
			// Trace: design.sv:32619:5
			reg [(2 ** (IdxW + 1)) - 2:0] mask_tree;
			// Trace: design.sv:32620:5
			reg [(((2 ** (IdxW + 1)) - 2) >= 0 ? (((2 ** (IdxW + 1)) - 1) * IdxW) - 1 : ((3 - (2 ** (IdxW + 1))) * IdxW) + ((((2 ** (IdxW + 1)) - 2) * IdxW) - 1)):(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : ((2 ** (IdxW + 1)) - 2) * IdxW)] idx_tree;
			// Trace: design.sv:32621:5
			reg [(((2 ** (IdxW + 1)) - 2) >= 0 ? (((2 ** (IdxW + 1)) - 1) * DW) - 1 : ((3 - (2 ** (IdxW + 1))) * DW) + ((((2 ** (IdxW + 1)) - 2) * DW) - 1)):(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : ((2 ** (IdxW + 1)) - 2) * DW)] data_tree;
			// Trace: design.sv:32622:5
			wire [N - 1:0] prio_mask_d;
			reg [N - 1:0] prio_mask_q;
			genvar _gv_level_6;
			for (_gv_level_6 = 0; _gv_level_6 < (IdxW + 1); _gv_level_6 = _gv_level_6 + 1) begin : gen_tree
				localparam level = _gv_level_6;
				// Trace: design.sv:32636:7
				localparam signed [31:0] Base0 = (2 ** level) - 1;
				// Trace: design.sv:32637:7
				localparam signed [31:0] Base1 = (2 ** (level + 1)) - 1;
				genvar _gv_offset_2;
				for (_gv_offset_2 = 0; _gv_offset_2 < (2 ** level); _gv_offset_2 = _gv_offset_2 + 1) begin : gen_level
					localparam offset = _gv_offset_2;
					// Trace: design.sv:32640:9
					localparam signed [31:0] Pa = Base0 + offset;
					// Trace: design.sv:32641:9
					localparam signed [31:0] C0 = Base1 + (2 * offset);
					// Trace: design.sv:32642:9
					localparam signed [31:0] C1 = (Base1 + (2 * offset)) + 1;
					if (level == IdxW) begin : gen_leafs
						if (offset < N) begin : gen_assign
							// Trace: design.sv:32650:13
							wire [1:1] sv2v_tmp_82807;
							assign sv2v_tmp_82807 = req_i[offset];
							always @(*) req_tree[Pa] = sv2v_tmp_82807;
							// Trace: design.sv:32656:13
							wire [1:1] sv2v_tmp_AA8F6;
							assign sv2v_tmp_AA8F6 = req_i[offset] & prio_mask_q[offset];
							always @(*) prio_tree[Pa] = sv2v_tmp_AA8F6;
							// Trace: design.sv:32658:13
							wire [IdxW * 1:1] sv2v_tmp_C9844;
							assign sv2v_tmp_C9844 = offset;
							always @(*) idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = sv2v_tmp_C9844;
							// Trace: design.sv:32660:13
							wire [DW * 1:1] sv2v_tmp_8A2B0;
							assign sv2v_tmp_8A2B0 = data_i[((N - 1) - offset) * DW+:DW];
							always @(*) data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = sv2v_tmp_8A2B0;
							// Trace: design.sv:32664:13
							assign gnt_o[offset] = (req_i[offset] & sel_tree[Pa]) & ready_i;
							// Trace: design.sv:32666:13
							assign prio_mask_d[offset] = (|req_i ? mask_tree[Pa] | (sel_tree[Pa] & ~ready_i) : prio_mask_q[offset]);
						end
						else begin : gen_tie_off
							// Trace: design.sv:32671:13
							wire [1:1] sv2v_tmp_DB8B3;
							assign sv2v_tmp_DB8B3 = 1'sb0;
							always @(*) req_tree[Pa] = sv2v_tmp_DB8B3;
							// Trace: design.sv:32672:13
							wire [1:1] sv2v_tmp_DFAC0;
							assign sv2v_tmp_DFAC0 = 1'sb0;
							always @(*) prio_tree[Pa] = sv2v_tmp_DFAC0;
							// Trace: design.sv:32673:13
							wire [IdxW * 1:1] sv2v_tmp_0FC8D;
							assign sv2v_tmp_0FC8D = 1'sb0;
							always @(*) idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = sv2v_tmp_0FC8D;
							// Trace: design.sv:32674:13
							wire [DW * 1:1] sv2v_tmp_8B097;
							assign sv2v_tmp_8B097 = 1'sb0;
							always @(*) data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = sv2v_tmp_8B097;
							// Trace: design.sv:32675:13
							wire unused_sigs;
							// Trace: design.sv:32676:13
							assign unused_sigs = ^{mask_tree[Pa], sel_tree[Pa]};
						end
					end
					else begin : gen_nodes
						// Trace: design.sv:32682:11
						reg sel;
						// Trace: design.sv:32683:11
						always @(*) begin : p_node
							if (_sv2v_0)
								;
							// Trace: design.sv:32686:13
							sel = ~req_tree[C0] | (~prio_tree[C0] & prio_tree[C1]);
							// Trace: design.sv:32688:13
							req_tree[Pa] = req_tree[C0] | req_tree[C1];
							// Trace: design.sv:32689:13
							prio_tree[Pa] = prio_tree[C1] | prio_tree[C0];
							// Trace: design.sv:32691:13
							idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = (sel ? idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C1 : ((2 ** (IdxW + 1)) - 2) - C1) * IdxW+:IdxW] : idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C0 : ((2 ** (IdxW + 1)) - 2) - C0) * IdxW+:IdxW]);
							// Trace: design.sv:32692:13
							data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = (sel ? data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C1 : ((2 ** (IdxW + 1)) - 2) - C1) * DW+:DW] : data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C0 : ((2 ** (IdxW + 1)) - 2) - C0) * DW+:DW]);
							// Trace: design.sv:32696:13
							sel_tree[C0] = sel_tree[Pa] & ~sel;
							// Trace: design.sv:32697:13
							sel_tree[C1] = sel_tree[Pa] & sel;
							// Trace: design.sv:32699:13
							mask_tree[C0] = mask_tree[Pa];
							// Trace: design.sv:32700:13
							mask_tree[C1] = mask_tree[Pa] | sel_tree[C0];
						end
					end
				end
			end
			if (EnDataPort) begin : gen_data_port
				// Trace: design.sv:32708:7
				assign data_o = data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * DW+:DW];
			end
			else begin : gen_no_dataport
				// Trace: design.sv:32710:7
				wire [DW - 1:0] unused_data;
				// Trace: design.sv:32711:7
				assign unused_data = data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * DW+:DW];
				// Trace: design.sv:32712:7
				assign data_o = 1'sb1;
			end
			// Trace: design.sv:32716:5
			wire unused_prio_tree;
			// Trace: design.sv:32717:5
			assign unused_prio_tree = prio_tree[0];
			// Trace: design.sv:32719:5
			assign idx_o = idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * IdxW+:IdxW];
			// Trace: design.sv:32720:5
			assign valid_o = req_tree[0];
			// Trace: design.sv:32723:5
			wire [1:1] sv2v_tmp_726FA;
			assign sv2v_tmp_726FA = 1'b1;
			always @(*) sel_tree[0] = sv2v_tmp_726FA;
			// Trace: design.sv:32725:5
			wire [1:1] sv2v_tmp_EA1F4;
			assign sv2v_tmp_EA1F4 = 1'b0;
			always @(*) mask_tree[0] = sv2v_tmp_EA1F4;
			// Trace: design.sv:32727:5
			always @(posedge clk_i or negedge rst_ni) begin : p_mask_reg
				// Trace: design.sv:32728:7
				if (!rst_ni)
					// Trace: design.sv:32729:9
					prio_mask_q <= 1'sb0;
				else
					// Trace: design.sv:32731:9
					prio_mask_q <= prio_mask_d;
			end
		end
	endgenerate
	// Trace: design.sv:32768:1
	// Trace: design.sv:32773:1
	initial _sv2v_0 = 0;
endmodule
module prim_arbiter_fixed (
	clk_i,
	rst_ni,
	req_i,
	data_i,
	gnt_o,
	idx_o,
	valid_o,
	data_o,
	ready_i
);
	reg _sv2v_0;
	// Trace: design.sv:32848:13
	parameter signed [31:0] N = 8;
	// Trace: design.sv:32849:13
	parameter signed [31:0] DW = 32;
	// Trace: design.sv:32853:13
	parameter [0:0] EnDataPort = 1;
	// Trace: design.sv:32856:14
	localparam signed [31:0] IdxW = $clog2(N);
	// Trace: design.sv:32859:3
	input clk_i;
	// Trace: design.sv:32860:3
	input rst_ni;
	// Trace: design.sv:32862:3
	input [N - 1:0] req_i;
	// Trace: design.sv:32863:3
	input [(N * DW) - 1:0] data_i;
	// Trace: design.sv:32864:3
	output wire [N - 1:0] gnt_o;
	// Trace: design.sv:32865:3
	output wire [IdxW - 1:0] idx_o;
	// Trace: design.sv:32867:3
	output wire valid_o;
	// Trace: design.sv:32868:3
	output wire [DW - 1:0] data_o;
	// Trace: design.sv:32869:3
	input ready_i;
	// Trace: design.sv:32875:3
	generate
		if (N == 1) begin : gen_degenerate_case
			// Trace: design.sv:32877:5
			assign valid_o = req_i[0];
			// Trace: design.sv:32878:5
			assign data_o = data_i[(N - 1) * DW+:DW];
			// Trace: design.sv:32879:5
			assign gnt_o[0] = valid_o & ready_i;
			// Trace: design.sv:32880:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_normal_case
			// Trace: design.sv:32886:5
			reg [(2 ** (IdxW + 1)) - 2:0] req_tree;
			// Trace: design.sv:32887:5
			reg [(2 ** (IdxW + 1)) - 2:0] gnt_tree;
			// Trace: design.sv:32888:5
			reg [(((2 ** (IdxW + 1)) - 2) >= 0 ? (((2 ** (IdxW + 1)) - 1) * IdxW) - 1 : ((3 - (2 ** (IdxW + 1))) * IdxW) + ((((2 ** (IdxW + 1)) - 2) * IdxW) - 1)):(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : ((2 ** (IdxW + 1)) - 2) * IdxW)] idx_tree;
			// Trace: design.sv:32889:5
			reg [(((2 ** (IdxW + 1)) - 2) >= 0 ? (((2 ** (IdxW + 1)) - 1) * DW) - 1 : ((3 - (2 ** (IdxW + 1))) * DW) + ((((2 ** (IdxW + 1)) - 2) * DW) - 1)):(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : ((2 ** (IdxW + 1)) - 2) * DW)] data_tree;
			genvar _gv_level_7;
			for (_gv_level_7 = 0; _gv_level_7 < (IdxW + 1); _gv_level_7 = _gv_level_7 + 1) begin : gen_tree
				localparam level = _gv_level_7;
				// Trace: design.sv:32903:7
				localparam signed [31:0] Base0 = (2 ** level) - 1;
				// Trace: design.sv:32904:7
				localparam signed [31:0] Base1 = (2 ** (level + 1)) - 1;
				genvar _gv_offset_3;
				for (_gv_offset_3 = 0; _gv_offset_3 < (2 ** level); _gv_offset_3 = _gv_offset_3 + 1) begin : gen_level
					localparam offset = _gv_offset_3;
					// Trace: design.sv:32907:9
					localparam signed [31:0] Pa = Base0 + offset;
					// Trace: design.sv:32908:9
					localparam signed [31:0] C0 = Base1 + (2 * offset);
					// Trace: design.sv:32909:9
					localparam signed [31:0] C1 = (Base1 + (2 * offset)) + 1;
					if (level == IdxW) begin : gen_leafs
						if (offset < N) begin : gen_assign
							// Trace: design.sv:32916:13
							wire [1:1] sv2v_tmp_82807;
							assign sv2v_tmp_82807 = req_i[offset];
							always @(*) req_tree[Pa] = sv2v_tmp_82807;
							// Trace: design.sv:32917:13
							wire [IdxW * 1:1] sv2v_tmp_82340;
							assign sv2v_tmp_82340 = offset;
							always @(*) idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = sv2v_tmp_82340;
							// Trace: design.sv:32918:13
							wire [DW * 1:1] sv2v_tmp_462FB;
							assign sv2v_tmp_462FB = data_i[((N - 1) - offset) * DW+:DW];
							always @(*) data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = sv2v_tmp_462FB;
							// Trace: design.sv:32920:13
							assign gnt_o[offset] = gnt_tree[Pa];
						end
						else begin : gen_tie_off
							// Trace: design.sv:32924:13
							wire [1:1] sv2v_tmp_DB8B3;
							assign sv2v_tmp_DB8B3 = 1'sb0;
							always @(*) req_tree[Pa] = sv2v_tmp_DB8B3;
							// Trace: design.sv:32925:13
							wire [IdxW * 1:1] sv2v_tmp_55789;
							assign sv2v_tmp_55789 = 1'sb0;
							always @(*) idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = sv2v_tmp_55789;
							// Trace: design.sv:32926:13
							wire [DW * 1:1] sv2v_tmp_DC98B;
							assign sv2v_tmp_DC98B = 1'sb0;
							always @(*) data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = sv2v_tmp_DC98B;
							// Trace: design.sv:32927:13
							wire unused_sigs;
							// Trace: design.sv:32928:13
							assign unused_sigs = gnt_tree[Pa];
						end
					end
					else begin : gen_nodes
						// Trace: design.sv:32933:11
						reg sel;
						// Trace: design.sv:32934:11
						always @(*) begin : p_node
							if (_sv2v_0)
								;
							// Trace: design.sv:32936:13
							sel = ~req_tree[C0];
							// Trace: design.sv:32938:13
							req_tree[Pa] = req_tree[C0] | req_tree[C1];
							// Trace: design.sv:32940:13
							idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = (sel ? idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C1 : ((2 ** (IdxW + 1)) - 2) - C1) * IdxW+:IdxW] : idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C0 : ((2 ** (IdxW + 1)) - 2) - C0) * IdxW+:IdxW]);
							// Trace: design.sv:32941:13
							data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = (sel ? data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C1 : ((2 ** (IdxW + 1)) - 2) - C1) * DW+:DW] : data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C0 : ((2 ** (IdxW + 1)) - 2) - C0) * DW+:DW]);
							// Trace: design.sv:32943:13
							gnt_tree[C0] = gnt_tree[Pa] & ~sel;
							// Trace: design.sv:32944:13
							gnt_tree[C1] = gnt_tree[Pa] & sel;
						end
					end
				end
			end
			if (EnDataPort) begin : gen_data_port
				// Trace: design.sv:32952:7
				assign data_o = data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * DW+:DW];
			end
			else begin : gen_no_dataport
				// Trace: design.sv:32954:7
				wire [DW - 1:0] unused_data;
				// Trace: design.sv:32955:7
				assign unused_data = data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * DW+:DW];
				// Trace: design.sv:32956:7
				assign data_o = 1'sb1;
			end
			// Trace: design.sv:32959:5
			assign idx_o = idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * IdxW+:IdxW];
			// Trace: design.sv:32960:5
			assign valid_o = req_tree[0];
			// Trace: design.sv:32963:5
			wire [1:1] sv2v_tmp_F03B8;
			assign sv2v_tmp_F03B8 = valid_o & ready_i;
			always @(*) gnt_tree[0] = sv2v_tmp_F03B8;
		end
	endgenerate
	// Trace: design.sv:32996:1
	initial _sv2v_0 = 0;
endmodule
module prim_subst_perm (
	data_i,
	key_i,
	data_o
);
	reg _sv2v_0;
	// Trace: design.sv:33014:13
	parameter signed [31:0] DataWidth = 64;
	// Trace: design.sv:33015:13
	parameter signed [31:0] NumRounds = 31;
	// Trace: design.sv:33016:13
	parameter [0:0] Decrypt = 0;
	// Trace: design.sv:33018:3
	input [DataWidth - 1:0] data_i;
	// Trace: design.sv:33019:3
	input [DataWidth - 1:0] key_i;
	// Trace: design.sv:33020:3
	output wire [DataWidth - 1:0] data_o;
	// Trace: design.sv:33033:3
	reg [(NumRounds >= 0 ? ((NumRounds + 1) * DataWidth) - 1 : ((1 - NumRounds) * DataWidth) + ((NumRounds * DataWidth) - 1)):(NumRounds >= 0 ? 0 : NumRounds * DataWidth)] data_state;
	// Trace: design.sv:33036:3
	wire [DataWidth * 1:1] sv2v_tmp_BB140;
	assign sv2v_tmp_BB140 = data_i;
	always @(*) data_state[(NumRounds >= 0 ? 0 : NumRounds) * DataWidth+:DataWidth] = sv2v_tmp_BB140;
	// Trace: design.sv:33038:3
	genvar _gv_r_2;
	localparam [63:0] prim_cipher_pkg_PRESENT_SBOX4 = 64'h21748fe3da09b65c;
	localparam [63:0] prim_cipher_pkg_PRESENT_SBOX4_INV = 64'ha970364bd21c8fe5;
	generate
		for (_gv_r_2 = 0; _gv_r_2 < NumRounds; _gv_r_2 = _gv_r_2 + 1) begin : gen_round
			localparam r = _gv_r_2;
			// Trace: design.sv:33039:5
			reg [DataWidth - 1:0] data_state_sbox;
			reg [DataWidth - 1:0] data_state_flipped;
			if (Decrypt) begin : gen_dec
				// Trace: design.sv:33043:7
				always @(*) begin : p_dec
					if (_sv2v_0)
						;
					// Trace: design.sv:33044:9
					data_state_sbox = data_state[(NumRounds >= 0 ? r : NumRounds - r) * DataWidth+:DataWidth] ^ key_i;
					// Trace: design.sv:33046:9
					data_state_flipped = data_state_sbox;
					// Trace: design.sv:33047:9
					begin : sv2v_autoblock_1
						// Trace: design.sv:33047:14
						reg signed [31:0] k;
						// Trace: design.sv:33047:14
						for (k = 0; k < (DataWidth / 2); k = k + 1)
							begin
								// Trace: design.sv:33048:11
								data_state_flipped[k * 2] = data_state_sbox[k];
								// Trace: design.sv:33049:11
								data_state_flipped[(k * 2) + 1] = data_state_sbox[k + (DataWidth / 2)];
							end
					end
					begin : sv2v_autoblock_2
						// Trace: design.sv:33052:14
						reg signed [31:0] k;
						// Trace: design.sv:33052:14
						for (k = 0; k < DataWidth; k = k + 1)
							begin
								// Trace: design.sv:33053:11
								data_state_sbox[(DataWidth - 1) - k] = data_state_flipped[k];
							end
					end
					begin : sv2v_autoblock_3
						// Trace: design.sv:33056:14
						reg signed [31:0] k;
						// Trace: design.sv:33056:14
						for (k = 0; k < (DataWidth / 4); k = k + 1)
							begin
								// Trace: design.sv:33057:11
								data_state_sbox[k * 4+:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[data_state_sbox[k * 4+:4] * 4+:4];
							end
					end
					// Trace: design.sv:33059:9
					data_state[(NumRounds >= 0 ? r + 1 : NumRounds - (r + 1)) * DataWidth+:DataWidth] = data_state_sbox;
				end
			end
			else begin : gen_enc
				// Trace: design.sv:33064:7
				always @(*) begin : p_enc
					if (_sv2v_0)
						;
					// Trace: design.sv:33065:9
					data_state_sbox = data_state[(NumRounds >= 0 ? r : NumRounds - r) * DataWidth+:DataWidth] ^ key_i;
					// Trace: design.sv:33069:9
					begin : sv2v_autoblock_4
						// Trace: design.sv:33069:14
						reg signed [31:0] k;
						// Trace: design.sv:33069:14
						for (k = 0; k < (DataWidth / 4); k = k + 1)
							begin
								// Trace: design.sv:33070:11
								data_state_sbox[k * 4+:4] = prim_cipher_pkg_PRESENT_SBOX4[data_state_sbox[k * 4+:4] * 4+:4];
							end
					end
					begin : sv2v_autoblock_5
						// Trace: design.sv:33073:14
						reg signed [31:0] k;
						// Trace: design.sv:33073:14
						for (k = 0; k < DataWidth; k = k + 1)
							begin
								// Trace: design.sv:33074:11
								data_state_flipped[(DataWidth - 1) - k] = data_state_sbox[k];
							end
					end
					// Trace: design.sv:33079:9
					data_state_sbox = data_state_flipped;
					begin : sv2v_autoblock_6
						// Trace: design.sv:33080:14
						reg signed [31:0] k;
						// Trace: design.sv:33080:14
						for (k = 0; k < (DataWidth / 2); k = k + 1)
							begin
								// Trace: design.sv:33081:11
								data_state_sbox[k] = data_state_flipped[k * 2];
								// Trace: design.sv:33082:11
								data_state_sbox[k + (DataWidth / 2)] = data_state_flipped[(k * 2) + 1];
							end
					end
					// Trace: design.sv:33084:9
					data_state[(NumRounds >= 0 ? r + 1 : NumRounds - (r + 1)) * DataWidth+:DataWidth] = data_state_sbox;
				end
			end
		end
	endgenerate
	// Trace: design.sv:33091:3
	assign data_o = data_state[(NumRounds >= 0 ? NumRounds : NumRounds - NumRounds) * DataWidth+:DataWidth] ^ key_i;
	initial _sv2v_0 = 0;
endmodule
module prim_present (
	data_i,
	key_i,
	idx_i,
	data_o,
	key_o,
	idx_o
);
	// Trace: design.sv:33119:13
	parameter signed [31:0] DataWidth = 64;
	// Trace: design.sv:33120:13
	parameter signed [31:0] KeyWidth = 128;
	// Trace: design.sv:33122:13
	parameter signed [31:0] NumRounds = 31;
	// Trace: design.sv:33128:13
	parameter signed [31:0] NumPhysRounds = NumRounds;
	// Trace: design.sv:33131:13
	parameter [0:0] Decrypt = 0;
	// Trace: design.sv:33133:3
	input [DataWidth - 1:0] data_i;
	// Trace: design.sv:33134:3
	input [KeyWidth - 1:0] key_i;
	// Trace: design.sv:33137:3
	input [4:0] idx_i;
	// Trace: design.sv:33138:3
	output wire [DataWidth - 1:0] data_o;
	// Trace: design.sv:33139:3
	output wire [KeyWidth - 1:0] key_o;
	// Trace: design.sv:33143:3
	output wire [4:0] idx_o;
	// Trace: design.sv:33150:3
	wire [(NumPhysRounds >= 0 ? ((NumPhysRounds + 1) * DataWidth) - 1 : ((1 - NumPhysRounds) * DataWidth) + ((NumPhysRounds * DataWidth) - 1)):(NumPhysRounds >= 0 ? 0 : NumPhysRounds * DataWidth)] data_state;
	// Trace: design.sv:33151:3
	wire [(NumPhysRounds >= 0 ? ((NumPhysRounds + 1) * KeyWidth) - 1 : ((1 - NumPhysRounds) * KeyWidth) + ((NumPhysRounds * KeyWidth) - 1)):(NumPhysRounds >= 0 ? 0 : NumPhysRounds * KeyWidth)] round_key;
	// Trace: design.sv:33152:3
	wire [(NumPhysRounds >= 0 ? ((NumPhysRounds + 1) * 5) - 1 : ((1 - NumPhysRounds) * 5) + ((NumPhysRounds * 5) - 1)):(NumPhysRounds >= 0 ? 0 : NumPhysRounds * 5)] round_idx;
	// Trace: design.sv:33155:3
	assign data_state[(NumPhysRounds >= 0 ? 0 : NumPhysRounds) * DataWidth+:DataWidth] = data_i;
	// Trace: design.sv:33156:3
	assign round_key[(NumPhysRounds >= 0 ? 0 : NumPhysRounds) * KeyWidth+:KeyWidth] = key_i;
	// Trace: design.sv:33157:3
	assign round_idx[(NumPhysRounds >= 0 ? 0 : NumPhysRounds) * 5+:5] = idx_i;
	// Trace: design.sv:33159:3
	genvar _gv_k_10;
	localparam [159:0] prim_cipher_pkg_PRESENT_PERM32 = 160'hfdde7f59c6ed5a5e5184dcd63d4942cc521c4100;
	localparam [159:0] prim_cipher_pkg_PRESENT_PERM32_INV = 160'hfeef37ace3f6ad2728c2ee6b16a4a1e629062080;
	localparam [383:0] prim_cipher_pkg_PRESENT_PERM64 = 384'hfef7cffae78ef6d74df2c70ceeb6cbeaa68ae69649e28608de75c7da6586d65545d24504ce34c3ca2482c61441c20400;
	localparam [383:0] prim_cipher_pkg_PRESENT_PERM64_INV = 384'hffbdf3beb9e37db5d33cb1c3fbadb2baa9a279a59238a182f79d71b69961759551349141f38d30b28920718510308100;
	localparam [63:0] prim_cipher_pkg_PRESENT_SBOX4 = 64'h21748fe3da09b65c;
	localparam [63:0] prim_cipher_pkg_PRESENT_SBOX4_INV = 64'ha970364bd21c8fe5;
	function automatic [31:0] prim_cipher_pkg_perm_32bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:379:46
		input reg [31:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:379:69
		input reg [159:0] perm;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:380:5
		reg [31:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:382:5
			begin : sv2v_autoblock_1
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:382:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:382:10
				for (k = 0; k < 32; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:383:7
						state_out[perm[k * 5+:5]] = state_in[k];
					end
			end
			prim_cipher_pkg_perm_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_perm_64bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:388:46
		input reg [63:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:388:69
		input reg [383:0] perm;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:389:5
		reg [63:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:391:5
			begin : sv2v_autoblock_2
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:391:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:391:10
				for (k = 0; k < 64; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:392:7
						state_out[perm[k * 6+:6]] = state_in[k];
					end
			end
			prim_cipher_pkg_perm_64bit = state_out;
		end
	endfunction
	function automatic [127:0] prim_cipher_pkg_present_inv_update_key128;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:271:62
		input reg [127:0] key_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:272:62
		input reg [4:0] round_idx;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:273:5
		reg [127:0] key_out;
		begin
			key_out = key_in;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:275:5
			key_out[66:62] = key_out[66:62] ^ round_idx;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:277:5
			key_out[123-:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[key_out[123-:4] * 4+:4];
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:279:5
			key_out[127-:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[key_out[127-:4] * 4+:4];
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:281:5
			key_out = {key_out[60:0], key_out[127:61]};
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:282:5
			prim_cipher_pkg_present_inv_update_key128 = key_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_present_inv_update_key64;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:247:60
		input reg [63:0] key_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:248:60
		input reg [4:0] round_idx;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:249:5
		reg [63:0] key_out;
		begin
			key_out = key_in;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:251:5
			key_out[19:15] = key_out[19:15] ^ round_idx;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:253:5
			key_out[63-:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[key_out[63-:4] * 4+:4];
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:255:5
			key_out = {key_out[60:0], key_out[63:61]};
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:256:5
			prim_cipher_pkg_present_inv_update_key64 = key_out;
		end
	endfunction
	function automatic [79:0] prim_cipher_pkg_present_inv_update_key80;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:259:60
		input reg [79:0] key_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:260:60
		input reg [4:0] round_idx;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:261:5
		reg [79:0] key_out;
		begin
			key_out = key_in;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:263:5
			key_out[19:15] = key_out[19:15] ^ round_idx;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:265:5
			key_out[79-:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[key_out[79-:4] * 4+:4];
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:267:5
			key_out = {key_out[60:0], key_out[79:61]};
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:268:5
			prim_cipher_pkg_present_inv_update_key80 = key_out;
		end
	endfunction
	function automatic [127:0] prim_cipher_pkg_present_update_key128;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:231:58
		input reg [127:0] key_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:232:58
		input reg [4:0] round_idx;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:233:5
		reg [127:0] key_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:235:5
			key_out = {key_in[66:0], key_in[127:67]};
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:237:5
			key_out[127-:4] = prim_cipher_pkg_PRESENT_SBOX4[key_out[127-:4] * 4+:4];
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:239:5
			key_out[123-:4] = prim_cipher_pkg_PRESENT_SBOX4[key_out[123-:4] * 4+:4];
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:241:5
			key_out[66:62] = key_out[66:62] ^ round_idx;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:242:5
			prim_cipher_pkg_present_update_key128 = key_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_present_update_key64;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:207:56
		input reg [63:0] key_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:208:56
		input reg [4:0] round_idx;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:209:5
		reg [63:0] key_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:211:5
			key_out = {key_in[2:0], key_in[63:3]};
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:213:5
			key_out[63-:4] = prim_cipher_pkg_PRESENT_SBOX4[key_out[63-:4] * 4+:4];
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:215:5
			key_out[19:15] = key_out[19:15] ^ round_idx;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:216:5
			prim_cipher_pkg_present_update_key64 = key_out;
		end
	endfunction
	function automatic [79:0] prim_cipher_pkg_present_update_key80;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:219:56
		input reg [79:0] key_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:220:56
		input reg [4:0] round_idx;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:221:5
		reg [79:0] key_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:223:5
			key_out = {key_in[18:0], key_in[79:19]};
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:225:5
			key_out[79-:4] = prim_cipher_pkg_PRESENT_SBOX4[key_out[79-:4] * 4+:4];
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:227:5
			key_out[19:15] = key_out[19:15] ^ round_idx;
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:228:5
			prim_cipher_pkg_present_update_key80 = key_out;
		end
	endfunction
	function automatic [7:0] prim_cipher_pkg_sbox4_8bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:325:45
		input reg [7:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:325:67
		input reg [63:0] sbox4;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:326:5
		reg [7:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:5
			begin : sv2v_autoblock_3
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:10
				for (k = 0; k < 2; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:329:7
						state_out[k * 4+:4] = sbox4[state_in[k * 4+:4] * 4+:4];
					end
			end
			prim_cipher_pkg_sbox4_8bit = state_out;
		end
	endfunction
	function automatic [31:0] prim_cipher_pkg_sbox4_32bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:343:47
		input reg [31:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:343:70
		input reg [63:0] sbox4;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:344:5
		reg [31:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:5
			begin : sv2v_autoblock_4
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:10
				for (k = 0; k < 4; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:347:7
						state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
					end
			end
			prim_cipher_pkg_sbox4_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_sbox4_64bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:352:47
		input reg [63:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:352:70
		input reg [63:0] sbox4;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:353:5
		reg [63:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:355:5
			begin : sv2v_autoblock_5
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:355:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:355:10
				for (k = 0; k < 8; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:356:7
						state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
					end
			end
			prim_cipher_pkg_sbox4_64bit = state_out;
		end
	endfunction
	generate
		for (_gv_k_10 = 0; _gv_k_10 < NumPhysRounds; _gv_k_10 = _gv_k_10 + 1) begin : gen_round
			localparam k = _gv_k_10;
			// Trace: design.sv:33160:5
			wire [DataWidth - 1:0] data_state_xor;
			wire [DataWidth - 1:0] data_state_sbox;
			// Trace: design.sv:33162:5
			assign data_state_xor = data_state[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * DataWidth+:DataWidth] ^ round_key[((NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth) + ((KeyWidth - 1) >= (KeyWidth - DataWidth) ? KeyWidth - 1 : ((KeyWidth - 1) + ((KeyWidth - 1) >= (KeyWidth - DataWidth) ? ((KeyWidth - 1) - (KeyWidth - DataWidth)) + 1 : ((KeyWidth - DataWidth) - (KeyWidth - 1)) + 1)) - 1)-:((KeyWidth - 1) >= (KeyWidth - DataWidth) ? ((KeyWidth - 1) - (KeyWidth - DataWidth)) + 1 : ((KeyWidth - DataWidth) - (KeyWidth - 1)) + 1)];
			if (Decrypt) begin : gen_dec
				// Trace: design.sv:33167:7
				assign round_idx[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * 5+:5] = round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5] - 1'b1;
				if (DataWidth == 64) begin : gen_d64
					// Trace: design.sv:33170:9
					assign data_state_sbox = prim_cipher_pkg_perm_64bit(data_state_xor, prim_cipher_pkg_PRESENT_PERM64_INV);
					// Trace: design.sv:33172:9
					assign data_state[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_64bit(data_state_sbox, prim_cipher_pkg_PRESENT_SBOX4_INV);
				end
				else begin : gen_d32
					// Trace: design.sv:33176:9
					assign data_state_sbox = prim_cipher_pkg_perm_32bit(data_state_xor, prim_cipher_pkg_PRESENT_PERM32_INV);
					// Trace: design.sv:33178:9
					assign data_state[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_32bit(data_state_sbox, prim_cipher_pkg_PRESENT_SBOX4_INV);
				end
				if (KeyWidth == 128) begin : gen_k128
					// Trace: design.sv:33184:9
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_inv_update_key128(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
				else if (KeyWidth == 80) begin : gen_k80
					// Trace: design.sv:33188:9
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_inv_update_key80(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
				else begin : gen_k64
					// Trace: design.sv:33192:9
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_inv_update_key64(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
			end
			else begin : gen_enc
				// Trace: design.sv:33199:7
				assign round_idx[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * 5+:5] = round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5] + 1'b1;
				if (DataWidth == 64) begin : gen_d64
					// Trace: design.sv:33202:9
					assign data_state_sbox = prim_cipher_pkg_sbox4_64bit(data_state_xor, prim_cipher_pkg_PRESENT_SBOX4);
					// Trace: design.sv:33204:9
					assign data_state[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_perm_64bit(data_state_sbox, prim_cipher_pkg_PRESENT_PERM64);
				end
				else begin : gen_d32
					// Trace: design.sv:33208:9
					assign data_state_sbox = prim_cipher_pkg_sbox4_32bit(data_state_xor, prim_cipher_pkg_PRESENT_SBOX4);
					// Trace: design.sv:33210:9
					assign data_state[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_perm_32bit(data_state_sbox, prim_cipher_pkg_PRESENT_PERM32);
				end
				if (KeyWidth == 128) begin : gen_k128
					// Trace: design.sv:33216:9
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_update_key128(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
				else if (KeyWidth == 80) begin : gen_k80
					// Trace: design.sv:33219:9
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_update_key80(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
				else begin : gen_k64
					// Trace: design.sv:33222:9
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_update_key64(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
			end
		end
	endgenerate
	// Trace: design.sv:33231:3
	localparam signed [31:0] LastRoundIdx = ((Decrypt != 0) || (NumRounds == 31) ? 0 : NumRounds + 1);
	// Trace: design.sv:33232:3
	assign data_o = (idx_o == LastRoundIdx ? data_state[(NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * DataWidth+:DataWidth] ^ round_key[((NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * KeyWidth) + ((KeyWidth - 1) >= (KeyWidth - DataWidth) ? KeyWidth - 1 : ((KeyWidth - 1) + ((KeyWidth - 1) >= (KeyWidth - DataWidth) ? ((KeyWidth - 1) - (KeyWidth - DataWidth)) + 1 : ((KeyWidth - DataWidth) - (KeyWidth - 1)) + 1)) - 1)-:((KeyWidth - 1) >= (KeyWidth - DataWidth) ? ((KeyWidth - 1) - (KeyWidth - DataWidth)) + 1 : ((KeyWidth - DataWidth) - (KeyWidth - 1)) + 1)] : data_state[(NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * DataWidth+:DataWidth]);
	// Trace: design.sv:33237:3
	assign key_o = round_key[(NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * KeyWidth+:KeyWidth];
	// Trace: design.sv:33238:3
	assign idx_o = round_idx[(NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * 5+:5];
endmodule
module prim_prince (
	clk_i,
	rst_ni,
	valid_i,
	data_i,
	key_i,
	dec_i,
	valid_o,
	data_o
);
	reg _sv2v_0;
	// Trace: design.sv:33278:13
	parameter signed [31:0] DataWidth = 64;
	// Trace: design.sv:33279:13
	parameter signed [31:0] KeyWidth = 128;
	// Trace: design.sv:33281:13
	parameter signed [31:0] NumRoundsHalf = 5;
	// Trace: design.sv:33284:13
	parameter [0:0] UseOldKeySched = 1'b0;
	// Trace: design.sv:33286:13
	parameter [0:0] HalfwayDataReg = 1'b0;
	// Trace: design.sv:33288:13
	parameter [0:0] HalfwayKeyReg = 1'b0;
	// Trace: design.sv:33290:3
	input clk_i;
	// Trace: design.sv:33291:3
	input rst_ni;
	// Trace: design.sv:33293:3
	input valid_i;
	// Trace: design.sv:33294:3
	input [DataWidth - 1:0] data_i;
	// Trace: design.sv:33295:3
	input [KeyWidth - 1:0] key_i;
	// Trace: design.sv:33296:3
	input dec_i;
	// Trace: design.sv:33297:3
	output wire valid_o;
	// Trace: design.sv:33298:3
	output reg [DataWidth - 1:0] data_o;
	// Trace: design.sv:33305:3
	reg [DataWidth - 1:0] k0;
	reg [DataWidth - 1:0] k0_prime_d;
	reg [DataWidth - 1:0] k1_d;
	reg [DataWidth - 1:0] k0_new_d;
	reg [DataWidth - 1:0] k0_prime_q;
	reg [DataWidth - 1:0] k1_q;
	reg [DataWidth - 1:0] k0_new_q;
	// Trace: design.sv:33306:3
	localparam [63:0] prim_cipher_pkg_PRINCE_ALPHA_CONST = 64'hc0ac29b7c97c50dd;
	always @(*) begin : p_key_expansion
		if (_sv2v_0)
			;
		// Trace: design.sv:33307:5
		k0 = key_i[(2 * DataWidth) - 1:DataWidth];
		// Trace: design.sv:33308:5
		k0_prime_d = {k0[0], k0[DataWidth - 1:2], k0[DataWidth - 1] ^ k0[1]};
		// Trace: design.sv:33309:5
		k1_d = key_i[DataWidth - 1:0];
		// Trace: design.sv:33312:5
		if (dec_i) begin
			// Trace: design.sv:33313:7
			k0 = k0_prime_d;
			// Trace: design.sv:33314:7
			k0_prime_d = key_i[(2 * DataWidth) - 1:DataWidth];
			// Trace: design.sv:33315:7
			k1_d = k1_d ^ prim_cipher_pkg_PRINCE_ALPHA_CONST[DataWidth - 1:0];
		end
	end
	// Trace: design.sv:33319:3
	generate
		if (UseOldKeySched) begin : gen_legacy_keyschedule
			// Trace: design.sv:33321:5
			wire [DataWidth:1] sv2v_tmp_003C5;
			assign sv2v_tmp_003C5 = k1_d;
			always @(*) k0_new_d = sv2v_tmp_003C5;
		end
		else begin : gen_new_keyschedule
			// Trace: design.sv:33325:5
			always @(*) begin : p_new_keyschedule_k0_alpha
				if (_sv2v_0)
					;
				// Trace: design.sv:33326:7
				k0_new_d = key_i[(2 * DataWidth) - 1:DataWidth];
				// Trace: design.sv:33328:7
				if (dec_i)
					// Trace: design.sv:33329:9
					k0_new_d = k0_new_d ^ prim_cipher_pkg_PRINCE_ALPHA_CONST[DataWidth - 1:0];
			end
		end
	endgenerate
	// Trace: design.sv:33334:3
	generate
		if (HalfwayKeyReg) begin : gen_key_reg
			// Trace: design.sv:33335:5
			always @(posedge clk_i or negedge rst_ni) begin : p_key_reg
				// Trace: design.sv:33336:7
				if (!rst_ni) begin
					// Trace: design.sv:33337:9
					k1_q <= 1'sb0;
					// Trace: design.sv:33338:9
					k0_prime_q <= 1'sb0;
					// Trace: design.sv:33339:9
					k0_new_q <= 1'sb0;
				end
				else
					// Trace: design.sv:33341:9
					if (valid_i) begin
						// Trace: design.sv:33342:11
						k1_q <= k1_d;
						// Trace: design.sv:33343:11
						k0_prime_q <= k0_prime_d;
						// Trace: design.sv:33344:11
						k0_new_q <= k0_new_d;
					end
			end
		end
		else begin : gen_no_key_reg
			// Trace: design.sv:33350:5
			wire [DataWidth:1] sv2v_tmp_6E066;
			assign sv2v_tmp_6E066 = k1_d;
			always @(*) k1_q = sv2v_tmp_6E066;
			// Trace: design.sv:33351:5
			wire [DataWidth:1] sv2v_tmp_BD8CA;
			assign sv2v_tmp_BD8CA = k0_prime_d;
			always @(*) k0_prime_q = sv2v_tmp_BD8CA;
			// Trace: design.sv:33352:5
			wire [DataWidth:1] sv2v_tmp_A995E;
			assign sv2v_tmp_A995E = k0_new_d;
			always @(*) k0_new_q = sv2v_tmp_A995E;
		end
	endgenerate
	// Trace: design.sv:33367:3
	reg [(((NumRoundsHalf * 2) + 1) >= 0 ? (((NumRoundsHalf * 2) + 2) * DataWidth) - 1 : ((1 - ((NumRoundsHalf * 2) + 1)) * DataWidth) + ((((NumRoundsHalf * 2) + 1) * DataWidth) - 1)):(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : ((NumRoundsHalf * 2) + 1) * DataWidth)] data_state;
	// Trace: design.sv:33370:3
	localparam [767:0] prim_cipher_pkg_PRINCE_ROUND_CONST = 768'hc0ac29b7c97c50ddd3b5a399ca0c239964a51195e0e3610dc882d32f25323c5485840851f1ac43aa7ef84f78fd955cb1be5466cf34e90c6c452821e638d01377082efa98ec4e6c89a4093822299f31d013198a2e037073440000000000000000;
	always @(*) begin : p_pre_round_xor
		if (_sv2v_0)
			;
		// Trace: design.sv:33371:5
		data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] = data_i ^ k0;
		// Trace: design.sv:33372:5
		data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] ^ k1_d;
		// Trace: design.sv:33373:5
		data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] ^ prim_cipher_pkg_PRINCE_ROUND_CONST[DataWidth - 1-:DataWidth];
	end
	// Trace: design.sv:33377:3
	genvar _gv_k_11;
	localparam [63:0] prim_cipher_pkg_PRINCE_SBOX4 = 64'h4d5e087619ca23fb;
	localparam [63:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS64 = 64'hfa50b61c72d83e94;
	localparam [15:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0 = 16'h7bde;
	localparam [15:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1 = 16'hbde7;
	localparam [15:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2 = 16'hde7b;
	localparam [15:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3 = 16'he7bd;
	function automatic [3:0] prim_cipher_pkg_prince_nibble_red16;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:89:54
		input reg [15:0] vect;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:90:5
		prim_cipher_pkg_prince_nibble_red16 = ((vect[0+:4] ^ vect[4+:4]) ^ vect[8+:4]) ^ vect[12+:4];
	endfunction
	function automatic [31:0] prim_cipher_pkg_prince_mult_prime_32bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:94:59
		input reg [31:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:95:5
		reg [31:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:97:5
			state_out[0+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:98:5
			state_out[4+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:99:5
			state_out[8+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:100:5
			state_out[12+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:102:5
			state_out[16+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:103:5
			state_out[20+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:104:5
			state_out[24+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:105:5
			state_out[28+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:106:5
			prim_cipher_pkg_prince_mult_prime_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_prince_mult_prime_64bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:110:59
		input reg [63:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:111:5
		reg [63:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:113:5
			state_out[0+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:114:5
			state_out[4+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:115:5
			state_out[8+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:116:5
			state_out[12+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:118:5
			state_out[16+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:119:5
			state_out[20+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:120:5
			state_out[24+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:121:5
			state_out[28+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:123:5
			state_out[32+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[32+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:124:5
			state_out[36+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[32+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:125:5
			state_out[40+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[32+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:126:5
			state_out[44+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[32+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:128:5
			state_out[48+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[48+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:129:5
			state_out[52+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[48+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:130:5
			state_out[56+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[48+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:131:5
			state_out[60+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[48+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:132:5
			prim_cipher_pkg_prince_mult_prime_64bit = state_out;
		end
	endfunction
	function automatic [31:0] prim_cipher_pkg_prince_shiftrows_32bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:67:58
		input reg [31:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:68:58
		input reg [63:0] shifts;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:69:5
		reg [31:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:71:5
			begin : sv2v_autoblock_1
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:71:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:71:10
				for (k = 0; k < 16; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:73:7
						state_out[k * 2+:2] = state_in[shifts[k * 4+:4] * 2+:2];
					end
			end
			prim_cipher_pkg_prince_shiftrows_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_prince_shiftrows_64bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:78:58
		input reg [63:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:79:58
		input reg [63:0] shifts;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:80:5
		reg [63:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:82:5
			begin : sv2v_autoblock_2
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:82:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:82:10
				for (k = 0; k < 16; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:83:7
						state_out[k * 4+:4] = state_in[shifts[k * 4+:4] * 4+:4];
					end
			end
			prim_cipher_pkg_prince_shiftrows_64bit = state_out;
		end
	endfunction
	function automatic [7:0] prim_cipher_pkg_sbox4_8bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:325:45
		input reg [7:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:325:67
		input reg [63:0] sbox4;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:326:5
		reg [7:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:5
			begin : sv2v_autoblock_3
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:10
				for (k = 0; k < 2; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:329:7
						state_out[k * 4+:4] = sbox4[state_in[k * 4+:4] * 4+:4];
					end
			end
			prim_cipher_pkg_sbox4_8bit = state_out;
		end
	endfunction
	function automatic [31:0] prim_cipher_pkg_sbox4_32bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:343:47
		input reg [31:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:343:70
		input reg [63:0] sbox4;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:344:5
		reg [31:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:5
			begin : sv2v_autoblock_4
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:10
				for (k = 0; k < 4; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:347:7
						state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
					end
			end
			prim_cipher_pkg_sbox4_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_sbox4_64bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:352:47
		input reg [63:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:352:70
		input reg [63:0] sbox4;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:353:5
		reg [63:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:355:5
			begin : sv2v_autoblock_5
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:355:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:355:10
				for (k = 0; k < 8; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:356:7
						state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
					end
			end
			prim_cipher_pkg_sbox4_64bit = state_out;
		end
	endfunction
	generate
		for (_gv_k_11 = 1; _gv_k_11 <= NumRoundsHalf; _gv_k_11 = _gv_k_11 + 1) begin : gen_fwd_pass
			localparam k = _gv_k_11;
			// Trace: design.sv:33378:5
			reg [DataWidth - 1:0] data_state_round;
			if (DataWidth == 64) begin : gen_fwd_d64
				// Trace: design.sv:33380:7
				always @(*) begin : p_fwd_d64
					if (_sv2v_0)
						;
					// Trace: design.sv:33381:9
					data_state_round = prim_cipher_pkg_sbox4_64bit(data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? k - 1 : ((NumRoundsHalf * 2) + 1) - (k - 1)) * DataWidth+:DataWidth], prim_cipher_pkg_PRINCE_SBOX4);
					// Trace: design.sv:33383:9
					data_state_round = prim_cipher_pkg_prince_mult_prime_64bit(data_state_round);
					// Trace: design.sv:33384:9
					data_state_round = prim_cipher_pkg_prince_shiftrows_64bit(data_state_round, prim_cipher_pkg_PRINCE_SHIFT_ROWS64);
				end
			end
			else begin : gen_fwd_d32
				// Trace: design.sv:33388:7
				always @(*) begin : p_fwd_d32
					if (_sv2v_0)
						;
					// Trace: design.sv:33389:9
					data_state_round = prim_cipher_pkg_sbox4_32bit(data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? k - 1 : ((NumRoundsHalf * 2) + 1) - (k - 1)) * DataWidth+:DataWidth], prim_cipher_pkg_PRINCE_SBOX4);
					// Trace: design.sv:33391:9
					data_state_round = prim_cipher_pkg_prince_mult_prime_32bit(data_state_round);
					// Trace: design.sv:33392:9
					data_state_round = prim_cipher_pkg_prince_shiftrows_32bit(data_state_round, prim_cipher_pkg_PRINCE_SHIFT_ROWS64);
				end
			end
			// Trace: design.sv:33396:5
			wire [DataWidth - 1:0] data_state_xor;
			// Trace: design.sv:33397:5
			assign data_state_xor = data_state_round ^ prim_cipher_pkg_PRINCE_ROUND_CONST[(k * 64) + (DataWidth - 1)-:DataWidth];
			if ((k % 2) == 1) begin : gen_fwd_key_odd
				// Trace: design.sv:33401:7
				wire [DataWidth * 1:1] sv2v_tmp_10B0B;
				assign sv2v_tmp_10B0B = data_state_xor ^ k0_new_d;
				always @(*) data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? k : ((NumRoundsHalf * 2) + 1) - k) * DataWidth+:DataWidth] = sv2v_tmp_10B0B;
			end
			else begin : gen_fwd_key_even
				// Trace: design.sv:33403:7
				wire [DataWidth * 1:1] sv2v_tmp_AB0D5;
				assign sv2v_tmp_AB0D5 = data_state_xor ^ k1_d;
				always @(*) data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? k : ((NumRoundsHalf * 2) + 1) - k) * DataWidth+:DataWidth] = sv2v_tmp_AB0D5;
			end
		end
	endgenerate
	// Trace: design.sv:33408:3
	reg [DataWidth - 1:0] data_state_middle_d;
	reg [DataWidth - 1:0] data_state_middle_q;
	reg [DataWidth - 1:0] data_state_middle;
	// Trace: design.sv:33409:3
	localparam [63:0] prim_cipher_pkg_PRINCE_SBOX4_INV = 64'h1ce5046a98df237b;
	generate
		if (DataWidth == 64) begin : gen_middle_d64
			// Trace: design.sv:33410:5
			always @(*) begin : p_middle_d64
				if (_sv2v_0)
					;
				// Trace: design.sv:33411:7
				data_state_middle_d = prim_cipher_pkg_sbox4_64bit(data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? NumRoundsHalf : ((NumRoundsHalf * 2) + 1) - NumRoundsHalf) * DataWidth+:DataWidth], prim_cipher_pkg_PRINCE_SBOX4);
				// Trace: design.sv:33413:7
				data_state_middle = prim_cipher_pkg_prince_mult_prime_64bit(data_state_middle_q);
				// Trace: design.sv:33414:7
				data_state_middle = prim_cipher_pkg_sbox4_64bit(data_state_middle, prim_cipher_pkg_PRINCE_SBOX4_INV);
			end
		end
		else begin : gen_middle_d32
			// Trace: design.sv:33418:5
			always @(*) begin : p_middle_d32
				if (_sv2v_0)
					;
				// Trace: design.sv:33419:7
				data_state_middle_d = prim_cipher_pkg_sbox4_32bit(data_state_middle[NumRoundsHalf], prim_cipher_pkg_PRINCE_SBOX4);
				// Trace: design.sv:33421:7
				data_state_middle = prim_cipher_pkg_prince_mult_prime_32bit(data_state_middle_q);
				// Trace: design.sv:33422:7
				data_state_middle = prim_cipher_pkg_sbox4_32bit(data_state_middle, prim_cipher_pkg_PRINCE_SBOX4_INV);
			end
		end
	endgenerate
	// Trace: design.sv:33427:3
	generate
		if (HalfwayDataReg) begin : gen_data_reg
			// Trace: design.sv:33428:5
			reg valid_q;
			// Trace: design.sv:33429:5
			always @(posedge clk_i or negedge rst_ni) begin : p_data_reg
				// Trace: design.sv:33430:7
				if (!rst_ni) begin
					// Trace: design.sv:33431:9
					valid_q <= 1'b0;
					// Trace: design.sv:33432:9
					data_state_middle_q <= 1'sb0;
				end
				else begin
					// Trace: design.sv:33434:9
					valid_q <= valid_i;
					// Trace: design.sv:33435:9
					if (valid_i)
						// Trace: design.sv:33436:11
						data_state_middle_q <= data_state_middle_d;
				end
			end
			// Trace: design.sv:33440:5
			assign valid_o = valid_q;
		end
		else begin : gen_no_data_reg
			// Trace: design.sv:33443:5
			wire [DataWidth:1] sv2v_tmp_F3D64;
			assign sv2v_tmp_F3D64 = data_state_middle_d;
			always @(*) data_state_middle_q = sv2v_tmp_F3D64;
			// Trace: design.sv:33444:5
			assign valid_o = valid_i;
		end
	endgenerate
	// Trace: design.sv:33447:3
	wire [DataWidth * 1:1] sv2v_tmp_93EC1;
	assign sv2v_tmp_93EC1 = data_state_middle;
	always @(*) data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? NumRoundsHalf + 1 : ((NumRoundsHalf * 2) + 1) - (NumRoundsHalf + 1)) * DataWidth+:DataWidth] = sv2v_tmp_93EC1;
	// Trace: design.sv:33450:3
	genvar _gv_k_12;
	localparam [63:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS64_INV = 64'hf258be147ad0369c;
	generate
		for (_gv_k_12 = 1; _gv_k_12 <= NumRoundsHalf; _gv_k_12 = _gv_k_12 + 1) begin : gen_bwd_pass
			localparam k = _gv_k_12;
			// Trace: design.sv:33451:5
			wire [DataWidth - 1:0] data_state_xor0;
			wire [DataWidth - 1:0] data_state_xor1;
			if ((((NumRoundsHalf + k) + 1) % 2) == 1) begin : gen_bkwd_key_odd
				// Trace: design.sv:33454:7
				assign data_state_xor0 = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? NumRoundsHalf + k : ((NumRoundsHalf * 2) + 1) - (NumRoundsHalf + k)) * DataWidth+:DataWidth] ^ k0_new_q;
			end
			else begin : gen_bkwd_key_even
				// Trace: design.sv:33456:7
				assign data_state_xor0 = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? NumRoundsHalf + k : ((NumRoundsHalf * 2) + 1) - (NumRoundsHalf + k)) * DataWidth+:DataWidth] ^ k1_q;
			end
			// Trace: design.sv:33459:5
			assign data_state_xor1 = data_state_xor0 ^ prim_cipher_pkg_PRINCE_ROUND_CONST[(((10 - NumRoundsHalf) + k) * 64) + (DataWidth - 1)-:DataWidth];
			// Trace: design.sv:33462:5
			reg [DataWidth - 1:0] data_state_bwd;
			if (DataWidth == 64) begin : gen_bwd_d64
				// Trace: design.sv:33464:7
				always @(*) begin : p_bwd_d64
					if (_sv2v_0)
						;
					// Trace: design.sv:33465:9
					data_state_bwd = prim_cipher_pkg_prince_shiftrows_64bit(data_state_xor1, prim_cipher_pkg_PRINCE_SHIFT_ROWS64_INV);
					// Trace: design.sv:33467:9
					data_state_bwd = prim_cipher_pkg_prince_mult_prime_64bit(data_state_bwd);
					// Trace: design.sv:33468:9
					data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? (NumRoundsHalf + k) + 1 : ((NumRoundsHalf * 2) + 1) - ((NumRoundsHalf + k) + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_64bit(data_state_bwd, prim_cipher_pkg_PRINCE_SBOX4_INV);
				end
			end
			else begin : gen_bwd_d32
				// Trace: design.sv:33472:7
				always @(*) begin : p_bwd_d32
					if (_sv2v_0)
						;
					// Trace: design.sv:33473:9
					data_state_bwd = prim_cipher_pkg_prince_shiftrows_32bit(data_state_xor1, prim_cipher_pkg_PRINCE_SHIFT_ROWS64_INV);
					// Trace: design.sv:33475:9
					data_state_bwd = prim_cipher_pkg_prince_mult_prime_32bit(data_state_bwd);
					// Trace: design.sv:33476:9
					data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? (NumRoundsHalf + k) + 1 : ((NumRoundsHalf * 2) + 1) - ((NumRoundsHalf + k) + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_32bit(data_state_bwd, prim_cipher_pkg_PRINCE_SBOX4_INV);
				end
			end
		end
	endgenerate
	// Trace: design.sv:33483:3
	always @(*) begin : p_post_round_xor
		if (_sv2v_0)
			;
		// Trace: design.sv:33484:5
		data_o = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? (2 * NumRoundsHalf) + 1 : ((NumRoundsHalf * 2) + 1) - ((2 * NumRoundsHalf) + 1)) * DataWidth+:DataWidth] ^ prim_cipher_pkg_PRINCE_ROUND_CONST[DataWidth + 703-:DataWidth];
		// Trace: design.sv:33486:5
		data_o = data_o ^ k1_q;
		// Trace: design.sv:33487:5
		data_o = data_o ^ k0_prime_q;
	end
	initial _sv2v_0 = 0;
endmodule
module prim_diff_decode (
	clk_i,
	rst_ni,
	diff_pi,
	diff_ni,
	level_o,
	rise_o,
	fall_o,
	event_o,
	sigint_o
);
	reg _sv2v_0;
	// Trace: design.sv:33521:13
	parameter [0:0] AsyncOn = 1'b0;
	// Trace: design.sv:33523:3
	input clk_i;
	// Trace: design.sv:33524:3
	input rst_ni;
	// Trace: design.sv:33526:3
	input diff_pi;
	// Trace: design.sv:33527:3
	input diff_ni;
	// Trace: design.sv:33530:3
	output wire level_o;
	// Trace: design.sv:33531:3
	output reg rise_o;
	// Trace: design.sv:33532:3
	output reg fall_o;
	// Trace: design.sv:33534:3
	output wire event_o;
	// Trace: design.sv:33536:3
	output reg sigint_o;
	// Trace: design.sv:33539:3
	reg level_d;
	reg level_q;
	// Trace: design.sv:33544:3
	generate
		if (AsyncOn) begin : gen_async
			// Trace: design.sv:33546:5
			// removed localparam type state_e
			// Trace: design.sv:33547:5
			reg [1:0] state_d;
			reg [1:0] state_q;
			// Trace: design.sv:33548:5
			wire diff_p_edge;
			wire diff_n_edge;
			wire diff_check_ok;
			wire level;
			// Trace: design.sv:33551:5
			reg diff_pq;
			reg diff_nq;
			wire diff_pd;
			wire diff_nd;
			// Trace: design.sv:33553:5
			prim_flop_2sync #(
				.Width(1),
				.ResetValue(1'sb0)
			) i_sync_p(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(diff_pi),
				.q_o(diff_pd)
			);
			// Trace: design.sv:33563:5
			prim_flop_2sync #(
				.Width(1),
				.ResetValue(1'b1)
			) i_sync_n(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(diff_ni),
				.q_o(diff_nd)
			);
			// Trace: design.sv:33574:5
			assign diff_p_edge = diff_pq ^ diff_pd;
			// Trace: design.sv:33575:5
			assign diff_n_edge = diff_nq ^ diff_nd;
			// Trace: design.sv:33578:5
			assign diff_check_ok = diff_pd ^ diff_nd;
			// Trace: design.sv:33581:5
			assign level = diff_pd;
			// Trace: design.sv:33584:5
			assign level_o = level_d;
			// Trace: design.sv:33585:5
			assign event_o = rise_o | fall_o;
			// Trace: design.sv:33606:5
			always @(*) begin : p_diff_fsm
				if (_sv2v_0)
					;
				// Trace: design.sv:33608:7
				state_d = state_q;
				// Trace: design.sv:33609:7
				level_d = level_q;
				// Trace: design.sv:33610:7
				rise_o = 1'b0;
				// Trace: design.sv:33611:7
				fall_o = 1'b0;
				// Trace: design.sv:33612:7
				sigint_o = 1'b0;
				// Trace: design.sv:33614:7
				(* full_case, parallel_case *)
				case (state_q)
					2'd0:
						// Trace: design.sv:33618:11
						if (diff_check_ok) begin
							// Trace: design.sv:33619:13
							level_d = level;
							// Trace: design.sv:33620:13
							if (diff_p_edge && diff_n_edge) begin
								begin
									// Trace: design.sv:33621:15
									if (level)
										// Trace: design.sv:33622:17
										rise_o = 1'b1;
									else
										// Trace: design.sv:33624:17
										fall_o = 1'b1;
								end
							end
						end
						else
							// Trace: design.sv:33628:13
							if (diff_p_edge || diff_n_edge)
								// Trace: design.sv:33629:15
								state_d = 2'd1;
							else begin
								// Trace: design.sv:33631:15
								state_d = 2'd2;
								// Trace: design.sv:33632:15
								sigint_o = 1'b1;
							end
					2'd1:
						// Trace: design.sv:33638:11
						if (diff_check_ok) begin
							// Trace: design.sv:33639:13
							state_d = 2'd0;
							// Trace: design.sv:33640:13
							level_d = level;
							// Trace: design.sv:33641:13
							if (level)
								// Trace: design.sv:33641:24
								rise_o = 1'b1;
							else
								// Trace: design.sv:33642:24
								fall_o = 1'b1;
						end
						else begin
							// Trace: design.sv:33644:13
							state_d = 2'd2;
							// Trace: design.sv:33645:13
							sigint_o = 1'b1;
						end
					2'd2: begin
						// Trace: design.sv:33651:11
						sigint_o = 1'b1;
						// Trace: design.sv:33652:11
						if (diff_check_ok) begin
							// Trace: design.sv:33653:13
							state_d = 2'd0;
							// Trace: design.sv:33654:13
							sigint_o = 1'b0;
						end
					end
					default:
						;
				endcase
			end
			// Trace: design.sv:33661:5
			always @(posedge clk_i or negedge rst_ni) begin : p_sync_reg
				// Trace: design.sv:33662:7
				if (!rst_ni) begin
					// Trace: design.sv:33663:9
					state_q <= 2'd0;
					// Trace: design.sv:33664:9
					diff_pq <= 1'b0;
					// Trace: design.sv:33665:9
					diff_nq <= 1'b1;
					// Trace: design.sv:33666:9
					level_q <= 1'b0;
				end
				else begin
					// Trace: design.sv:33668:9
					state_q <= state_d;
					// Trace: design.sv:33669:9
					diff_pq <= diff_pd;
					// Trace: design.sv:33670:9
					diff_nq <= diff_nd;
					// Trace: design.sv:33671:9
					level_q <= level_d;
				end
			end
		end
		else begin : gen_no_async
			// Trace: design.sv:33679:5
			reg diff_pq;
			wire diff_pd;
			// Trace: design.sv:33682:5
			assign diff_pd = diff_pi;
			// Trace: design.sv:33685:5
			wire [1:1] sv2v_tmp_5CA36;
			assign sv2v_tmp_5CA36 = ~(diff_pi ^ diff_ni);
			always @(*) sigint_o = sv2v_tmp_5CA36;
			// Trace: design.sv:33687:5
			assign level_o = (sigint_o ? level_q : diff_pi);
			// Trace: design.sv:33688:5
			wire [1:1] sv2v_tmp_AB662;
			assign sv2v_tmp_AB662 = level_o;
			always @(*) level_d = sv2v_tmp_AB662;
			// Trace: design.sv:33691:5
			wire [1:1] sv2v_tmp_8926B;
			assign sv2v_tmp_8926B = (~diff_pq & diff_pi) & ~sigint_o;
			always @(*) rise_o = sv2v_tmp_8926B;
			// Trace: design.sv:33692:5
			wire [1:1] sv2v_tmp_A5341;
			assign sv2v_tmp_A5341 = (diff_pq & ~diff_pi) & ~sigint_o;
			always @(*) fall_o = sv2v_tmp_A5341;
			// Trace: design.sv:33693:5
			assign event_o = rise_o | fall_o;
			// Trace: design.sv:33695:5
			always @(posedge clk_i or negedge rst_ni) begin : p_edge_reg
				// Trace: design.sv:33696:7
				if (!rst_ni) begin
					// Trace: design.sv:33697:9
					diff_pq <= 1'b0;
					// Trace: design.sv:33698:9
					level_q <= 1'b0;
				end
				else begin
					// Trace: design.sv:33700:9
					diff_pq <= diff_pd;
					// Trace: design.sv:33701:9
					level_q <= level_d;
				end
			end
		end
	endgenerate
	// Trace: design.sv:33719:3
	initial _sv2v_0 = 0;
endmodule
module prim_generic_clock_mux2 (
	clk0_i,
	clk1_i,
	sel_i,
	clk_o
);
	// Trace: design.sv:33767:13
	parameter [0:0] NoFpgaBufG = 1'b0;
	// Trace: design.sv:33769:3
	input clk0_i;
	// Trace: design.sv:33770:3
	input clk1_i;
	// Trace: design.sv:33771:3
	input sel_i;
	// Trace: design.sv:33772:3
	output wire clk_o;
	// Trace: design.sv:33775:3
	assign clk_o = (sel_i ? clk1_i : clk0_i);
endmodule
// removed package "tlul_pkg"
module ibex_alu (
	operator_i,
	operand_a_i,
	operand_b_i,
	instr_first_cycle_i,
	multdiv_operand_a_i,
	multdiv_operand_b_i,
	multdiv_sel_i,
	imd_val_q_i,
	imd_val_d_o,
	imd_val_we_o,
	adder_result_o,
	adder_result_ext_o,
	result_o,
	comparison_result_o,
	is_equal_result_o
);
	reg _sv2v_0;
	// Trace: design.sv:33979:13
	// removed localparam type ibex_pkg_rv32b_e
	parameter integer RV32B = 32'sd0;
	// Trace: design.sv:33981:3
	// removed localparam type ibex_pkg_alu_op_e
	input wire [6:0] operator_i;
	// Trace: design.sv:33982:3
	input wire [31:0] operand_a_i;
	// Trace: design.sv:33983:3
	input wire [31:0] operand_b_i;
	// Trace: design.sv:33985:3
	input wire instr_first_cycle_i;
	// Trace: design.sv:33987:3
	input wire [32:0] multdiv_operand_a_i;
	// Trace: design.sv:33988:3
	input wire [32:0] multdiv_operand_b_i;
	// Trace: design.sv:33990:3
	input wire multdiv_sel_i;
	// Trace: design.sv:33992:3
	input wire [63:0] imd_val_q_i;
	// Trace: design.sv:33993:3
	output reg [63:0] imd_val_d_o;
	// Trace: design.sv:33994:3
	output reg [1:0] imd_val_we_o;
	// Trace: design.sv:33996:3
	output wire [31:0] adder_result_o;
	// Trace: design.sv:33997:3
	output wire [33:0] adder_result_ext_o;
	// Trace: design.sv:33999:3
	output reg [31:0] result_o;
	// Trace: design.sv:34000:3
	output wire comparison_result_o;
	// Trace: design.sv:34001:3
	output wire is_equal_result_o;
	// Trace: design.sv:34003:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:34005:3
	wire [31:0] operand_a_rev;
	// Trace: design.sv:34006:3
	wire [32:0] operand_b_neg;
	// Trace: design.sv:34009:3
	genvar _gv_k_13;
	generate
		for (_gv_k_13 = 0; _gv_k_13 < 32; _gv_k_13 = _gv_k_13 + 1) begin : gen_rev_operand_a
			localparam k = _gv_k_13;
			// Trace: design.sv:34010:5
			assign operand_a_rev[k] = operand_a_i[31 - k];
		end
	endgenerate
	// Trace: design.sv:34017:3
	reg adder_op_a_shift1;
	// Trace: design.sv:34018:3
	reg adder_op_a_shift2;
	// Trace: design.sv:34019:3
	reg adder_op_a_shift3;
	// Trace: design.sv:34020:3
	reg adder_op_b_negate;
	// Trace: design.sv:34021:3
	reg [32:0] adder_in_a;
	reg [32:0] adder_in_b;
	// Trace: design.sv:34022:3
	wire [31:0] adder_result;
	// Trace: design.sv:34024:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34025:5
		adder_op_a_shift1 = 1'b0;
		// Trace: design.sv:34026:5
		adder_op_a_shift2 = 1'b0;
		// Trace: design.sv:34027:5
		adder_op_a_shift3 = 1'b0;
		// Trace: design.sv:34028:5
		adder_op_b_negate = 1'b0;
		// Trace: design.sv:34029:5
		(* full_case, parallel_case *)
		case (operator_i)
			7'd1, 7'd29, 7'd30, 7'd27, 7'd28, 7'd25, 7'd26, 7'd43, 7'd44, 7'd31, 7'd32, 7'd33, 7'd34:
				// Trace: design.sv:34041:27
				adder_op_b_negate = 1'b1;
			7'd22:
				if (RV32B != 32'sd0)
					// Trace: design.sv:34044:43
					adder_op_a_shift1 = 1'b1;
			7'd23:
				if (RV32B != 32'sd0)
					// Trace: design.sv:34045:43
					adder_op_a_shift2 = 1'b1;
			7'd24:
				if (RV32B != 32'sd0)
					// Trace: design.sv:34046:43
					adder_op_a_shift3 = 1'b1;
			default:
				;
		endcase
	end
	// Trace: design.sv:34053:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34054:5
		(* full_case, parallel_case *)
		case (1'b1)
			multdiv_sel_i:
				// Trace: design.sv:34055:26
				adder_in_a = multdiv_operand_a_i;
			adder_op_a_shift1:
				// Trace: design.sv:34056:26
				adder_in_a = {operand_a_i[30:0], 2'b01};
			adder_op_a_shift2:
				// Trace: design.sv:34057:26
				adder_in_a = {operand_a_i[29:0], 3'b001};
			adder_op_a_shift3:
				// Trace: design.sv:34058:26
				adder_in_a = {operand_a_i[28:0], 4'b0001};
			default:
				// Trace: design.sv:34059:26
				adder_in_a = {operand_a_i, 1'b1};
		endcase
	end
	// Trace: design.sv:34064:3
	assign operand_b_neg = {operand_b_i, 1'b0} ^ {33 {1'b1}};
	// Trace: design.sv:34065:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34066:5
		(* full_case, parallel_case *)
		case (1'b1)
			multdiv_sel_i:
				// Trace: design.sv:34067:26
				adder_in_b = multdiv_operand_b_i;
			adder_op_b_negate:
				// Trace: design.sv:34068:26
				adder_in_b = operand_b_neg;
			default:
				// Trace: design.sv:34069:26
				adder_in_b = {operand_b_i, 1'b0};
		endcase
	end
	// Trace: design.sv:34074:3
	assign adder_result_ext_o = $unsigned(adder_in_a) + $unsigned(adder_in_b);
	// Trace: design.sv:34076:3
	assign adder_result = adder_result_ext_o[32:1];
	// Trace: design.sv:34078:3
	assign adder_result_o = adder_result;
	// Trace: design.sv:34084:3
	wire is_equal;
	// Trace: design.sv:34085:3
	reg is_greater_equal;
	// Trace: design.sv:34086:3
	reg cmp_signed;
	// Trace: design.sv:34088:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34089:5
		(* full_case, parallel_case *)
		case (operator_i)
			7'd27, 7'd25, 7'd43, 7'd31, 7'd33:
				// Trace: design.sv:34095:16
				cmp_signed = 1'b1;
			default:
				// Trace: design.sv:34097:16
				cmp_signed = 1'b0;
		endcase
	end
	// Trace: design.sv:34101:3
	assign is_equal = adder_result == 32'b00000000000000000000000000000000;
	// Trace: design.sv:34102:3
	assign is_equal_result_o = is_equal;
	// Trace: design.sv:34105:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34106:5
		if ((operand_a_i[31] ^ operand_b_i[31]) == 1'b0)
			// Trace: design.sv:34107:7
			is_greater_equal = adder_result[31] == 1'b0;
		else
			// Trace: design.sv:34109:7
			is_greater_equal = operand_a_i[31] ^ cmp_signed;
	end
	// Trace: design.sv:34126:3
	reg cmp_result;
	// Trace: design.sv:34128:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34129:5
		(* full_case, parallel_case *)
		case (operator_i)
			7'd29:
				// Trace: design.sv:34130:27
				cmp_result = is_equal;
			7'd30:
				// Trace: design.sv:34131:27
				cmp_result = ~is_equal;
			7'd27, 7'd28, 7'd33, 7'd34:
				// Trace: design.sv:34133:27
				cmp_result = is_greater_equal;
			7'd25, 7'd26, 7'd31, 7'd32, 7'd43, 7'd44:
				// Trace: design.sv:34136:27
				cmp_result = ~is_greater_equal;
			default:
				// Trace: design.sv:34138:16
				cmp_result = is_equal;
		endcase
	end
	// Trace: design.sv:34142:3
	assign comparison_result_o = cmp_result;
	// Trace: design.sv:34211:3
	reg shift_left;
	// Trace: design.sv:34212:3
	wire shift_ones;
	// Trace: design.sv:34213:3
	wire shift_arith;
	// Trace: design.sv:34214:3
	wire shift_funnel;
	// Trace: design.sv:34215:3
	wire shift_sbmode;
	// Trace: design.sv:34216:3
	reg [5:0] shift_amt;
	// Trace: design.sv:34217:3
	wire [5:0] shift_amt_compl;
	// Trace: design.sv:34219:3
	reg [31:0] shift_operand;
	// Trace: design.sv:34220:3
	reg signed [32:0] shift_result_ext_signed;
	// Trace: design.sv:34221:3
	reg [32:0] shift_result_ext;
	// Trace: design.sv:34222:3
	reg unused_shift_result_ext;
	// Trace: design.sv:34223:3
	reg [31:0] shift_result;
	// Trace: design.sv:34224:3
	reg [31:0] shift_result_rev;
	// Trace: design.sv:34227:3
	wire bfp_op;
	// Trace: design.sv:34228:3
	wire [4:0] bfp_len;
	// Trace: design.sv:34229:3
	wire [4:0] bfp_off;
	// Trace: design.sv:34230:3
	wire [31:0] bfp_mask;
	// Trace: design.sv:34231:3
	wire [31:0] bfp_mask_rev;
	// Trace: design.sv:34232:3
	wire [31:0] bfp_result;
	// Trace: design.sv:34235:3
	assign bfp_op = (RV32B != 32'sd0 ? operator_i == 7'd55 : 1'b0);
	// Trace: design.sv:34236:3
	assign bfp_len = {~(|operand_b_i[27:24]), operand_b_i[27:24]};
	// Trace: design.sv:34237:3
	assign bfp_off = operand_b_i[20:16];
	// Trace: design.sv:34238:3
	assign bfp_mask = (RV32B != 32'sd0 ? ~(32'hffffffff << bfp_len) : {32 {1'sb0}});
	// Trace: design.sv:34239:3
	genvar _gv_i_38;
	generate
		for (_gv_i_38 = 0; _gv_i_38 < 32; _gv_i_38 = _gv_i_38 + 1) begin : gen_rev_bfp_mask
			localparam i = _gv_i_38;
			// Trace: design.sv:34240:5
			assign bfp_mask_rev[i] = bfp_mask[31 - i];
		end
	endgenerate
	// Trace: design.sv:34243:3
	assign bfp_result = (RV32B != 32'sd0 ? (~shift_result & operand_a_i) | ((operand_b_i & bfp_mask) << bfp_off) : {32 {1'sb0}});
	// Trace: design.sv:34248:3
	wire [1:1] sv2v_tmp_BA5F8;
	assign sv2v_tmp_BA5F8 = operand_b_i[5] & shift_funnel;
	always @(*) shift_amt[5] = sv2v_tmp_BA5F8;
	// Trace: design.sv:34249:3
	assign shift_amt_compl = 32 - operand_b_i[4:0];
	// Trace: design.sv:34251:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34252:5
		if (bfp_op)
			// Trace: design.sv:34253:7
			shift_amt[4:0] = bfp_off;
		else
			// Trace: design.sv:34255:7
			shift_amt[4:0] = (instr_first_cycle_i ? (operand_b_i[5] && shift_funnel ? shift_amt_compl[4:0] : operand_b_i[4:0]) : (operand_b_i[5] && shift_funnel ? operand_b_i[4:0] : shift_amt_compl[4:0]));
	end
	// Trace: design.sv:34262:3
	assign shift_sbmode = (RV32B != 32'sd0 ? ((operator_i == 7'd49) | (operator_i == 7'd50)) | (operator_i == 7'd51) : 1'b0);
	// Trace: design.sv:34273:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34274:5
		(* full_case, parallel_case *)
		case (operator_i)
			7'd10:
				// Trace: design.sv:34275:16
				shift_left = 1'b1;
			7'd12:
				// Trace: design.sv:34276:16
				shift_left = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b1 : 1'b0);
			7'd55:
				// Trace: design.sv:34277:16
				shift_left = (RV32B != 32'sd0 ? 1'b1 : 1'b0);
			7'd14:
				// Trace: design.sv:34278:16
				shift_left = (RV32B != 32'sd0 ? instr_first_cycle_i : 0);
			7'd13:
				// Trace: design.sv:34279:16
				shift_left = (RV32B != 32'sd0 ? ~instr_first_cycle_i : 0);
			7'd47:
				// Trace: design.sv:34280:16
				shift_left = (RV32B != 32'sd0 ? (shift_amt[5] ? ~instr_first_cycle_i : instr_first_cycle_i) : 1'b0);
			7'd48:
				// Trace: design.sv:34282:16
				shift_left = (RV32B != 32'sd0 ? (shift_amt[5] ? instr_first_cycle_i : ~instr_first_cycle_i) : 1'b0);
			default:
				// Trace: design.sv:34284:16
				shift_left = 1'b0;
		endcase
		if (shift_sbmode)
			// Trace: design.sv:34287:7
			shift_left = 1'b1;
	end
	// Trace: design.sv:34291:3
	assign shift_arith = operator_i == 7'd8;
	// Trace: design.sv:34292:3
	assign shift_ones = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? (operator_i == 7'd12) | (operator_i == 7'd11) : 1'b0);
	// Trace: design.sv:34294:3
	assign shift_funnel = (RV32B != 32'sd0 ? (operator_i == 7'd47) | (operator_i == 7'd48) : 1'b0);
	// Trace: design.sv:34298:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34301:5
		if (RV32B == 32'sd0)
			// Trace: design.sv:34302:7
			shift_operand = (shift_left ? operand_a_rev : operand_a_i);
		else
			// Trace: design.sv:34304:7
			(* full_case, parallel_case *)
			case (1'b1)
				bfp_op:
					// Trace: design.sv:34305:23
					shift_operand = bfp_mask_rev;
				shift_sbmode:
					// Trace: design.sv:34306:23
					shift_operand = 32'h80000000;
				default:
					// Trace: design.sv:34307:23
					shift_operand = (shift_left ? operand_a_rev : operand_a_i);
			endcase
		// Trace: design.sv:34311:5
		shift_result_ext_signed = $signed({shift_ones | (shift_arith & shift_operand[31]), shift_operand}) >>> shift_amt[4:0];
		// Trace: design.sv:34313:5
		shift_result_ext = $unsigned(shift_result_ext_signed);
		// Trace: design.sv:34315:5
		shift_result = shift_result_ext[31:0];
		// Trace: design.sv:34316:5
		unused_shift_result_ext = shift_result_ext[32];
		begin : sv2v_autoblock_1
			// Trace: design.sv:34318:10
			reg [31:0] i;
			// Trace: design.sv:34318:10
			for (i = 0; i < 32; i = i + 1)
				begin
					// Trace: design.sv:34319:7
					shift_result_rev[i] = shift_result[31 - i];
				end
		end
		// Trace: design.sv:34322:5
		shift_result = (shift_left ? shift_result_rev : shift_result);
	end
	// Trace: design.sv:34330:3
	wire bwlogic_or;
	// Trace: design.sv:34331:3
	wire bwlogic_and;
	// Trace: design.sv:34332:3
	wire [31:0] bwlogic_operand_b;
	// Trace: design.sv:34333:3
	wire [31:0] bwlogic_or_result;
	// Trace: design.sv:34334:3
	wire [31:0] bwlogic_and_result;
	// Trace: design.sv:34335:3
	wire [31:0] bwlogic_xor_result;
	// Trace: design.sv:34336:3
	reg [31:0] bwlogic_result;
	// Trace: design.sv:34338:3
	reg bwlogic_op_b_negate;
	// Trace: design.sv:34340:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34341:5
		(* full_case, parallel_case *)
		case (operator_i)
			7'd5, 7'd6, 7'd7:
				// Trace: design.sv:34345:17
				bwlogic_op_b_negate = (RV32B != 32'sd0 ? 1'b1 : 1'b0);
			7'd46:
				// Trace: design.sv:34346:17
				bwlogic_op_b_negate = (RV32B != 32'sd0 ? ~instr_first_cycle_i : 1'b0);
			default:
				// Trace: design.sv:34347:17
				bwlogic_op_b_negate = 1'b0;
		endcase
	end
	// Trace: design.sv:34351:3
	assign bwlogic_operand_b = (bwlogic_op_b_negate ? operand_b_neg[32:1] : operand_b_i);
	// Trace: design.sv:34353:3
	assign bwlogic_or_result = operand_a_i | bwlogic_operand_b;
	// Trace: design.sv:34354:3
	assign bwlogic_and_result = operand_a_i & bwlogic_operand_b;
	// Trace: design.sv:34355:3
	assign bwlogic_xor_result = operand_a_i ^ bwlogic_operand_b;
	// Trace: design.sv:34357:3
	assign bwlogic_or = (operator_i == 7'd3) | (operator_i == 7'd6);
	// Trace: design.sv:34358:3
	assign bwlogic_and = (operator_i == 7'd4) | (operator_i == 7'd7);
	// Trace: design.sv:34360:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:34361:5
		(* full_case, parallel_case *)
		case (1'b1)
			bwlogic_or:
				// Trace: design.sv:34362:20
				bwlogic_result = bwlogic_or_result;
			bwlogic_and:
				// Trace: design.sv:34363:20
				bwlogic_result = bwlogic_and_result;
			default:
				// Trace: design.sv:34364:20
				bwlogic_result = bwlogic_xor_result;
		endcase
	end
	// Trace: design.sv:34368:3
	wire [5:0] bitcnt_result;
	// Trace: design.sv:34369:3
	wire [31:0] minmax_result;
	// Trace: design.sv:34370:3
	reg [31:0] pack_result;
	// Trace: design.sv:34371:3
	wire [31:0] sext_result;
	// Trace: design.sv:34372:3
	reg [31:0] singlebit_result;
	// Trace: design.sv:34373:3
	reg [31:0] rev_result;
	// Trace: design.sv:34374:3
	reg [31:0] shuffle_result;
	// Trace: design.sv:34375:3
	wire [31:0] xperm_result;
	// Trace: design.sv:34376:3
	reg [31:0] butterfly_result;
	// Trace: design.sv:34377:3
	reg [31:0] invbutterfly_result;
	// Trace: design.sv:34378:3
	reg [31:0] clmul_result;
	// Trace: design.sv:34379:3
	reg [31:0] multicycle_result;
	// Trace: design.sv:34381:3
	generate
		if (RV32B != 32'sd0) begin : g_alu_rvb
			// Trace: design.sv:34392:5
			wire zbe_op;
			// Trace: design.sv:34393:5
			wire bitcnt_ctz;
			// Trace: design.sv:34394:5
			wire bitcnt_clz;
			// Trace: design.sv:34395:5
			wire bitcnt_cz;
			// Trace: design.sv:34396:5
			reg [31:0] bitcnt_bits;
			// Trace: design.sv:34397:5
			wire [31:0] bitcnt_mask_op;
			// Trace: design.sv:34398:5
			reg [31:0] bitcnt_bit_mask;
			// Trace: design.sv:34399:5
			reg [191:0] bitcnt_partial;
			// Trace: design.sv:34400:5
			wire [31:0] bitcnt_partial_lsb_d;
			// Trace: design.sv:34401:5
			wire [31:0] bitcnt_partial_msb_d;
			// Trace: design.sv:34404:5
			assign bitcnt_ctz = operator_i == 7'd41;
			// Trace: design.sv:34405:5
			assign bitcnt_clz = operator_i == 7'd40;
			// Trace: design.sv:34406:5
			assign bitcnt_cz = bitcnt_ctz | bitcnt_clz;
			// Trace: design.sv:34407:5
			assign bitcnt_result = bitcnt_partial[0+:6];
			// Trace: design.sv:34413:5
			assign bitcnt_mask_op = (bitcnt_clz ? operand_a_rev : operand_a_i);
			// Trace: design.sv:34415:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:34416:7
				bitcnt_bit_mask = bitcnt_mask_op;
				// Trace: design.sv:34417:7
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 1);
				// Trace: design.sv:34418:7
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 2);
				// Trace: design.sv:34419:7
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 4);
				// Trace: design.sv:34420:7
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 8);
				// Trace: design.sv:34421:7
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 16);
				// Trace: design.sv:34422:7
				bitcnt_bit_mask = ~bitcnt_bit_mask;
			end
			// Trace: design.sv:34425:5
			assign zbe_op = (operator_i == 7'd53) | (operator_i == 7'd54);
			// Trace: design.sv:34427:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:34428:7
				case (1'b1)
					zbe_op:
						// Trace: design.sv:34429:22
						bitcnt_bits = operand_b_i;
					bitcnt_cz:
						// Trace: design.sv:34430:22
						bitcnt_bits = bitcnt_bit_mask & ~bitcnt_mask_op;
					default:
						// Trace: design.sv:34431:22
						bitcnt_bits = operand_a_i;
				endcase
			end
			// Trace: design.sv:34476:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:34477:7
				bitcnt_partial = {32 {6'b000000}};
				// Trace: design.sv:34479:7
				begin : sv2v_autoblock_2
					// Trace: design.sv:34479:12
					reg [31:0] i;
					// Trace: design.sv:34479:12
					for (i = 1; i < 32; i = i + 2)
						begin
							// Trace: design.sv:34480:9
							bitcnt_partial[(31 - i) * 6+:6] = {5'h00, bitcnt_bits[i]} + {5'h00, bitcnt_bits[i - 1]};
						end
				end
				begin : sv2v_autoblock_3
					// Trace: design.sv:34483:12
					reg [31:0] i;
					// Trace: design.sv:34483:12
					for (i = 3; i < 32; i = i + 4)
						begin
							// Trace: design.sv:34484:9
							bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(33 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
						end
				end
				begin : sv2v_autoblock_4
					// Trace: design.sv:34487:12
					reg [31:0] i;
					// Trace: design.sv:34487:12
					for (i = 7; i < 32; i = i + 8)
						begin
							// Trace: design.sv:34488:9
							bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(35 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
						end
				end
				begin : sv2v_autoblock_5
					// Trace: design.sv:34491:12
					reg [31:0] i;
					// Trace: design.sv:34491:12
					for (i = 15; i < 32; i = i + 16)
						begin
							// Trace: design.sv:34492:9
							bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(39 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
						end
				end
				// Trace: design.sv:34495:7
				bitcnt_partial[0+:6] = bitcnt_partial[96+:6] + bitcnt_partial[0+:6];
				// Trace: design.sv:34499:7
				bitcnt_partial[48+:6] = bitcnt_partial[96+:6] + bitcnt_partial[48+:6];
				begin : sv2v_autoblock_6
					// Trace: design.sv:34502:12
					reg [31:0] i;
					// Trace: design.sv:34502:12
					for (i = 11; i < 32; i = i + 8)
						begin
							// Trace: design.sv:34503:9
							bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(35 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
						end
				end
				begin : sv2v_autoblock_7
					// Trace: design.sv:34507:12
					reg [31:0] i;
					// Trace: design.sv:34507:12
					for (i = 5; i < 32; i = i + 4)
						begin
							// Trace: design.sv:34508:9
							bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(33 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
						end
				end
				// Trace: design.sv:34511:7
				bitcnt_partial[186+:6] = {5'h00, bitcnt_bits[0]};
				begin : sv2v_autoblock_8
					// Trace: design.sv:34512:12
					reg [31:0] i;
					// Trace: design.sv:34512:12
					for (i = 2; i < 32; i = i + 2)
						begin
							// Trace: design.sv:34513:9
							bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(32 - i) * 6+:6] + {5'h00, bitcnt_bits[i]};
						end
				end
			end
			// Trace: design.sv:34521:5
			assign minmax_result = (cmp_result ? operand_a_i : operand_b_i);
			// Trace: design.sv:34527:5
			wire packu;
			// Trace: design.sv:34528:5
			wire packh;
			// Trace: design.sv:34529:5
			assign packu = operator_i == 7'd36;
			// Trace: design.sv:34530:5
			assign packh = operator_i == 7'd37;
			// Trace: design.sv:34532:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:34533:7
				(* full_case, parallel_case *)
				case (1'b1)
					packu:
						// Trace: design.sv:34534:18
						pack_result = {operand_b_i[31:16], operand_a_i[31:16]};
					packh:
						// Trace: design.sv:34535:18
						pack_result = {16'h0000, operand_b_i[7:0], operand_a_i[7:0]};
					default:
						// Trace: design.sv:34536:18
						pack_result = {operand_b_i[15:0], operand_a_i[15:0]};
				endcase
			end
			// Trace: design.sv:34544:5
			assign sext_result = (operator_i == 7'd38 ? {{24 {operand_a_i[7]}}, operand_a_i[7:0]} : {{16 {operand_a_i[15]}}, operand_a_i[15:0]});
			// Trace: design.sv:34551:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:34552:7
				(* full_case, parallel_case *)
				case (operator_i)
					7'd49:
						// Trace: design.sv:34553:19
						singlebit_result = operand_a_i | shift_result;
					7'd50:
						// Trace: design.sv:34554:19
						singlebit_result = operand_a_i & ~shift_result;
					7'd51:
						// Trace: design.sv:34555:19
						singlebit_result = operand_a_i ^ shift_result;
					default:
						// Trace: design.sv:34556:19
						singlebit_result = {31'h00000000, shift_result[0]};
				endcase
			end
			// Trace: design.sv:34568:5
			wire [4:0] zbp_shift_amt;
			// Trace: design.sv:34569:5
			wire gorc_op;
			// Trace: design.sv:34571:5
			assign gorc_op = operator_i == 7'd16;
			// Trace: design.sv:34572:5
			assign zbp_shift_amt[2:0] = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? shift_amt[2:0] : {3 {shift_amt[0]}});
			// Trace: design.sv:34574:5
			assign zbp_shift_amt[4:3] = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? shift_amt[4:3] : {2 {shift_amt[3]}});
			// Trace: design.sv:34577:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:34578:7
				rev_result = operand_a_i;
				// Trace: design.sv:34580:7
				if (zbp_shift_amt[0])
					// Trace: design.sv:34581:9
					rev_result = ((gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h55555555) << 1)) | ((rev_result & 32'haaaaaaaa) >> 1);
				if (zbp_shift_amt[1])
					// Trace: design.sv:34587:9
					rev_result = ((gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h33333333) << 2)) | ((rev_result & 32'hcccccccc) >> 2);
				if (zbp_shift_amt[2])
					// Trace: design.sv:34593:9
					rev_result = ((gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h0f0f0f0f) << 4)) | ((rev_result & 32'hf0f0f0f0) >> 4);
				if (zbp_shift_amt[3])
					// Trace: design.sv:34599:9
					rev_result = ((((RV32B == 32'sd2) || (RV32B == 32'sd3)) && gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h00ff00ff) << 8)) | ((rev_result & 32'hff00ff00) >> 8);
				if (zbp_shift_amt[4])
					// Trace: design.sv:34606:9
					rev_result = ((((RV32B == 32'sd2) || (RV32B == 32'sd3)) && gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h0000ffff) << 16)) | ((rev_result & 32'hffff0000) >> 16);
			end
			// Trace: design.sv:34613:5
			wire crc_hmode;
			// Trace: design.sv:34614:5
			wire crc_bmode;
			// Trace: design.sv:34615:5
			wire [31:0] clmul_result_rev;
			if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin : gen_alu_rvb_otearlgrey_full
				// Trace: design.sv:34623:7
				localparam [127:0] SHUFFLE_MASK_L = 128'h00ff00000f000f003030303044444444;
				// Trace: design.sv:34625:7
				localparam [127:0] SHUFFLE_MASK_R = 128'h0000ff0000f000f00c0c0c0c22222222;
				// Trace: design.sv:34628:7
				localparam [127:0] FLIP_MASK_L = 128'h22001100004400004411000011000000;
				// Trace: design.sv:34630:7
				localparam [127:0] FLIP_MASK_R = 128'h00880044000022000000882200000088;
				// Trace: design.sv:34633:7
				wire [31:0] SHUFFLE_MASK_NOT [0:3];
				genvar _gv_i_39;
				for (_gv_i_39 = 0; _gv_i_39 < 4; _gv_i_39 = _gv_i_39 + 1) begin : gen_shuffle_mask_not
					localparam i = _gv_i_39;
					// Trace: design.sv:34635:9
					assign SHUFFLE_MASK_NOT[i] = ~(SHUFFLE_MASK_L[(3 - i) * 32+:32] | SHUFFLE_MASK_R[(3 - i) * 32+:32]);
				end
				// Trace: design.sv:34638:7
				wire shuffle_flip;
				// Trace: design.sv:34639:7
				assign shuffle_flip = operator_i == 7'd18;
				// Trace: design.sv:34641:7
				reg [3:0] shuffle_mode;
				// Trace: design.sv:34643:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:34644:9
					shuffle_result = operand_a_i;
					// Trace: design.sv:34646:9
					if (shuffle_flip) begin
						// Trace: design.sv:34647:11
						shuffle_mode[3] = shift_amt[0];
						// Trace: design.sv:34648:11
						shuffle_mode[2] = shift_amt[1];
						// Trace: design.sv:34649:11
						shuffle_mode[1] = shift_amt[2];
						// Trace: design.sv:34650:11
						shuffle_mode[0] = shift_amt[3];
					end
					else
						// Trace: design.sv:34652:11
						shuffle_mode = shift_amt[3:0];
					if (shuffle_flip)
						// Trace: design.sv:34656:11
						shuffle_result = ((((((((shuffle_result & 32'h88224411) | ((shuffle_result << 6) & FLIP_MASK_L[96+:32])) | ((shuffle_result >> 6) & FLIP_MASK_R[96+:32])) | ((shuffle_result << 9) & FLIP_MASK_L[64+:32])) | ((shuffle_result >> 9) & FLIP_MASK_R[64+:32])) | ((shuffle_result << 15) & FLIP_MASK_L[32+:32])) | ((shuffle_result >> 15) & FLIP_MASK_R[32+:32])) | ((shuffle_result << 21) & FLIP_MASK_L[0+:32])) | ((shuffle_result >> 21) & FLIP_MASK_R[0+:32]);
					if (shuffle_mode[3])
						// Trace: design.sv:34668:11
						shuffle_result = (shuffle_result & SHUFFLE_MASK_NOT[0]) | (((shuffle_result << 8) & SHUFFLE_MASK_L[96+:32]) | ((shuffle_result >> 8) & SHUFFLE_MASK_R[96+:32]));
					if (shuffle_mode[2])
						// Trace: design.sv:34673:11
						shuffle_result = (shuffle_result & SHUFFLE_MASK_NOT[1]) | (((shuffle_result << 4) & SHUFFLE_MASK_L[64+:32]) | ((shuffle_result >> 4) & SHUFFLE_MASK_R[64+:32]));
					if (shuffle_mode[1])
						// Trace: design.sv:34678:11
						shuffle_result = (shuffle_result & SHUFFLE_MASK_NOT[2]) | (((shuffle_result << 2) & SHUFFLE_MASK_L[32+:32]) | ((shuffle_result >> 2) & SHUFFLE_MASK_R[32+:32]));
					if (shuffle_mode[0])
						// Trace: design.sv:34683:11
						shuffle_result = (shuffle_result & SHUFFLE_MASK_NOT[3]) | (((shuffle_result << 1) & SHUFFLE_MASK_L[0+:32]) | ((shuffle_result >> 1) & SHUFFLE_MASK_R[0+:32]));
					if (shuffle_flip)
						// Trace: design.sv:34689:11
						shuffle_result = ((((((((shuffle_result & 32'h88224411) | ((shuffle_result << 6) & FLIP_MASK_L[96+:32])) | ((shuffle_result >> 6) & FLIP_MASK_R[96+:32])) | ((shuffle_result << 9) & FLIP_MASK_L[64+:32])) | ((shuffle_result >> 9) & FLIP_MASK_R[64+:32])) | ((shuffle_result << 15) & FLIP_MASK_L[32+:32])) | ((shuffle_result >> 15) & FLIP_MASK_R[32+:32])) | ((shuffle_result << 21) & FLIP_MASK_L[0+:32])) | ((shuffle_result >> 21) & FLIP_MASK_R[0+:32]);
				end
				// Trace: design.sv:34711:7
				wire [23:0] sel_n;
				// Trace: design.sv:34712:7
				wire [7:0] vld_n;
				// Trace: design.sv:34713:7
				wire [7:0] sel_b;
				// Trace: design.sv:34714:7
				wire [3:0] vld_b;
				// Trace: design.sv:34715:7
				wire [1:0] sel_h;
				// Trace: design.sv:34716:7
				wire [1:0] vld_h;
				genvar _gv_i_40;
				for (_gv_i_40 = 0; _gv_i_40 < 8; _gv_i_40 = _gv_i_40 + 1) begin : gen_sel_vld_n
					localparam i = _gv_i_40;
					// Trace: design.sv:34722:9
					assign sel_n[i * 3+:3] = operand_b_i[i * 4+:3];
					// Trace: design.sv:34723:9
					assign vld_n[i] = ~|operand_b_i[(i * 4) + 3+:1];
				end
				genvar _gv_i_41;
				for (_gv_i_41 = 0; _gv_i_41 < 4; _gv_i_41 = _gv_i_41 + 1) begin : gen_sel_vld_b
					localparam i = _gv_i_41;
					// Trace: design.sv:34730:9
					assign sel_b[i * 2+:2] = operand_b_i[i * 8+:2];
					// Trace: design.sv:34731:9
					assign vld_b[i] = ~|operand_b_i[(i * 8) + 2+:6];
				end
				genvar _gv_i_42;
				for (_gv_i_42 = 0; _gv_i_42 < 2; _gv_i_42 = _gv_i_42 + 1) begin : gen_sel_vld_h
					localparam i = _gv_i_42;
					// Trace: design.sv:34738:9
					assign sel_h[i+:1] = operand_b_i[i * 16+:1];
					// Trace: design.sv:34739:9
					assign vld_h[i] = ~|operand_b_i[(i * 16) + 1+:15];
				end
				// Trace: design.sv:34744:7
				reg [23:0] sel;
				// Trace: design.sv:34745:7
				reg [7:0] vld;
				// Trace: design.sv:34746:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:34747:9
					(* full_case, parallel_case *)
					case (operator_i)
						7'd19: begin
							// Trace: design.sv:34750:13
							sel = sel_n;
							// Trace: design.sv:34751:13
							vld = vld_n;
						end
						7'd20:
							// Trace: design.sv:34756:13
							begin : sv2v_autoblock_9
								// Trace: design.sv:34756:18
								reg signed [31:0] b;
								// Trace: design.sv:34756:18
								for (b = 0; b < 4; b = b + 1)
									begin
										// Trace: design.sv:34757:15
										sel[((b * 2) + 0) * 3+:3] = {sel_b[b * 2+:2], 1'b0};
										// Trace: design.sv:34758:15
										sel[((b * 2) + 1) * 3+:3] = {sel_b[b * 2+:2], 1'b1};
										// Trace: design.sv:34759:15
										vld[b * 2+:2] = {2 {vld_b[b]}};
									end
							end
						7'd21:
							// Trace: design.sv:34765:13
							begin : sv2v_autoblock_10
								// Trace: design.sv:34765:18
								reg signed [31:0] h;
								// Trace: design.sv:34765:18
								for (h = 0; h < 2; h = h + 1)
									begin
										// Trace: design.sv:34766:15
										sel[((h * 4) + 0) * 3+:3] = {sel_h[h+:1], 2'b00};
										// Trace: design.sv:34767:15
										sel[((h * 4) + 1) * 3+:3] = {sel_h[h+:1], 2'b01};
										// Trace: design.sv:34768:15
										sel[((h * 4) + 2) * 3+:3] = {sel_h[h+:1], 2'b10};
										// Trace: design.sv:34769:15
										sel[((h * 4) + 3) * 3+:3] = {sel_h[h+:1], 2'b11};
										// Trace: design.sv:34770:15
										vld[h * 4+:4] = {4 {vld_h[h]}};
									end
							end
						default: begin
							// Trace: design.sv:34776:13
							sel = sel_n;
							// Trace: design.sv:34777:13
							vld = 1'sb0;
						end
					endcase
				end
				// Trace: design.sv:34783:7
				wire [31:0] val_n;
				// Trace: design.sv:34784:7
				wire [31:0] xperm_n;
				// Trace: design.sv:34785:7
				assign val_n = operand_a_i;
				genvar _gv_i_43;
				for (_gv_i_43 = 0; _gv_i_43 < 8; _gv_i_43 = _gv_i_43 + 1) begin : gen_xperm_n
					localparam i = _gv_i_43;
					// Trace: design.sv:34787:9
					assign xperm_n[i * 4+:4] = (vld[i] ? val_n[sel[i * 3+:3] * 4+:4] : {4 {1'sb0}});
				end
				// Trace: design.sv:34789:7
				assign xperm_result = xperm_n;
				// Trace: design.sv:34852:7
				wire clmul_rmode;
				// Trace: design.sv:34853:7
				wire clmul_hmode;
				// Trace: design.sv:34854:7
				reg [31:0] clmul_op_a;
				// Trace: design.sv:34855:7
				reg [31:0] clmul_op_b;
				// Trace: design.sv:34856:7
				wire [31:0] operand_b_rev;
				// Trace: design.sv:34857:7
				wire [31:0] clmul_and_stage [0:31];
				// Trace: design.sv:34858:7
				wire [31:0] clmul_xor_stage1 [0:15];
				// Trace: design.sv:34859:7
				wire [31:0] clmul_xor_stage2 [0:7];
				// Trace: design.sv:34860:7
				wire [31:0] clmul_xor_stage3 [0:3];
				// Trace: design.sv:34861:7
				wire [31:0] clmul_xor_stage4 [0:1];
				// Trace: design.sv:34863:7
				wire [31:0] clmul_result_raw;
				genvar _gv_i_44;
				for (_gv_i_44 = 0; _gv_i_44 < 32; _gv_i_44 = _gv_i_44 + 1) begin : gen_rev_operand_b
					localparam i = _gv_i_44;
					// Trace: design.sv:34866:9
					assign operand_b_rev[i] = operand_b_i[31 - i];
				end
				// Trace: design.sv:34869:7
				assign clmul_rmode = operator_i == 7'd57;
				// Trace: design.sv:34870:7
				assign clmul_hmode = operator_i == 7'd58;
				// Trace: design.sv:34873:7
				localparam [31:0] CRC32_POLYNOMIAL = 32'h04c11db7;
				// Trace: design.sv:34874:7
				localparam [31:0] CRC32_MU_REV = 32'hf7011641;
				// Trace: design.sv:34876:7
				localparam [31:0] CRC32C_POLYNOMIAL = 32'h1edc6f41;
				// Trace: design.sv:34877:7
				localparam [31:0] CRC32C_MU_REV = 32'hdea713f1;
				// Trace: design.sv:34879:7
				wire crc_op;
				// Trace: design.sv:34881:7
				wire crc_cpoly;
				// Trace: design.sv:34883:7
				reg [31:0] crc_operand;
				// Trace: design.sv:34884:7
				wire [31:0] crc_poly;
				// Trace: design.sv:34885:7
				wire [31:0] crc_mu_rev;
				// Trace: design.sv:34887:7
				assign crc_op = (((((operator_i == 7'd64) | (operator_i == 7'd63)) | (operator_i == 7'd62)) | (operator_i == 7'd61)) | (operator_i == 7'd60)) | (operator_i == 7'd59);
				// Trace: design.sv:34891:7
				assign crc_cpoly = ((operator_i == 7'd64) | (operator_i == 7'd62)) | (operator_i == 7'd60);
				// Trace: design.sv:34895:7
				assign crc_hmode = (operator_i == 7'd61) | (operator_i == 7'd62);
				// Trace: design.sv:34896:7
				assign crc_bmode = (operator_i == 7'd59) | (operator_i == 7'd60);
				// Trace: design.sv:34898:7
				assign crc_poly = (crc_cpoly ? CRC32C_POLYNOMIAL : CRC32_POLYNOMIAL);
				// Trace: design.sv:34899:7
				assign crc_mu_rev = (crc_cpoly ? CRC32C_MU_REV : CRC32_MU_REV);
				// Trace: design.sv:34901:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:34902:9
					(* full_case, parallel_case *)
					case (1'b1)
						crc_bmode:
							// Trace: design.sv:34903:22
							crc_operand = {operand_a_i[7:0], 24'h000000};
						crc_hmode:
							// Trace: design.sv:34904:22
							crc_operand = {operand_a_i[15:0], 16'h0000};
						default:
							// Trace: design.sv:34905:22
							crc_operand = operand_a_i;
					endcase
				end
				// Trace: design.sv:34910:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:34911:9
					if (crc_op) begin
						// Trace: design.sv:34912:11
						clmul_op_a = (instr_first_cycle_i ? crc_operand : imd_val_q_i[32+:32]);
						// Trace: design.sv:34913:11
						clmul_op_b = (instr_first_cycle_i ? crc_mu_rev : crc_poly);
					end
					else begin
						// Trace: design.sv:34915:11
						clmul_op_a = (clmul_rmode | clmul_hmode ? operand_a_rev : operand_a_i);
						// Trace: design.sv:34916:11
						clmul_op_b = (clmul_rmode | clmul_hmode ? operand_b_rev : operand_b_i);
					end
				end
				genvar _gv_i_45;
				for (_gv_i_45 = 0; _gv_i_45 < 32; _gv_i_45 = _gv_i_45 + 1) begin : gen_clmul_and_op
					localparam i = _gv_i_45;
					// Trace: design.sv:34921:9
					assign clmul_and_stage[i] = (clmul_op_b[i] ? clmul_op_a << i : {32 {1'sb0}});
				end
				genvar _gv_i_46;
				for (_gv_i_46 = 0; _gv_i_46 < 16; _gv_i_46 = _gv_i_46 + 1) begin : gen_clmul_xor_op_l1
					localparam i = _gv_i_46;
					// Trace: design.sv:34925:9
					assign clmul_xor_stage1[i] = clmul_and_stage[2 * i] ^ clmul_and_stage[(2 * i) + 1];
				end
				genvar _gv_i_47;
				for (_gv_i_47 = 0; _gv_i_47 < 8; _gv_i_47 = _gv_i_47 + 1) begin : gen_clmul_xor_op_l2
					localparam i = _gv_i_47;
					// Trace: design.sv:34929:9
					assign clmul_xor_stage2[i] = clmul_xor_stage1[2 * i] ^ clmul_xor_stage1[(2 * i) + 1];
				end
				genvar _gv_i_48;
				for (_gv_i_48 = 0; _gv_i_48 < 4; _gv_i_48 = _gv_i_48 + 1) begin : gen_clmul_xor_op_l3
					localparam i = _gv_i_48;
					// Trace: design.sv:34933:9
					assign clmul_xor_stage3[i] = clmul_xor_stage2[2 * i] ^ clmul_xor_stage2[(2 * i) + 1];
				end
				genvar _gv_i_49;
				for (_gv_i_49 = 0; _gv_i_49 < 2; _gv_i_49 = _gv_i_49 + 1) begin : gen_clmul_xor_op_l4
					localparam i = _gv_i_49;
					// Trace: design.sv:34937:9
					assign clmul_xor_stage4[i] = clmul_xor_stage3[2 * i] ^ clmul_xor_stage3[(2 * i) + 1];
				end
				// Trace: design.sv:34940:7
				assign clmul_result_raw = clmul_xor_stage4[0] ^ clmul_xor_stage4[1];
				genvar _gv_i_50;
				for (_gv_i_50 = 0; _gv_i_50 < 32; _gv_i_50 = _gv_i_50 + 1) begin : gen_rev_clmul_result
					localparam i = _gv_i_50;
					// Trace: design.sv:34943:9
					assign clmul_result_rev[i] = clmul_result_raw[31 - i];
				end
				// Trace: design.sv:34948:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:34949:9
					case (1'b1)
						clmul_rmode:
							// Trace: design.sv:34950:24
							clmul_result = clmul_result_rev;
						clmul_hmode:
							// Trace: design.sv:34951:24
							clmul_result = {1'b0, clmul_result_rev[31:1]};
						default:
							// Trace: design.sv:34952:24
							clmul_result = clmul_result_raw;
					endcase
				end
			end
			else begin : gen_alu_rvb_not_otearlgrey_full
				// Trace: design.sv:34956:7
				wire [32:1] sv2v_tmp_4A308;
				assign sv2v_tmp_4A308 = 1'sb0;
				always @(*) shuffle_result = sv2v_tmp_4A308;
				// Trace: design.sv:34957:7
				assign xperm_result = 1'sb0;
				// Trace: design.sv:34958:7
				wire [32:1] sv2v_tmp_31DA6;
				assign sv2v_tmp_31DA6 = 1'sb0;
				always @(*) clmul_result = sv2v_tmp_31DA6;
				// Trace: design.sv:34960:7
				assign clmul_result_rev = 1'sb0;
				// Trace: design.sv:34961:7
				assign crc_bmode = 1'sb0;
				// Trace: design.sv:34962:7
				assign crc_hmode = 1'sb0;
			end
			if (RV32B == 32'sd3) begin : gen_alu_rvb_full
				// Trace: design.sv:35019:7
				reg [191:0] bitcnt_partial_q;
				genvar _gv_i_51;
				for (_gv_i_51 = 0; _gv_i_51 < 32; _gv_i_51 = _gv_i_51 + 1) begin : gen_bitcnt_reg_in_lsb
					localparam i = _gv_i_51;
					// Trace: design.sv:35024:9
					assign bitcnt_partial_lsb_d[i] = bitcnt_partial[(31 - i) * 6];
				end
				genvar _gv_i_52;
				for (_gv_i_52 = 0; _gv_i_52 < 16; _gv_i_52 = _gv_i_52 + 1) begin : gen_bitcnt_reg_in_b1
					localparam i = _gv_i_52;
					// Trace: design.sv:35028:9
					assign bitcnt_partial_msb_d[i] = bitcnt_partial[((31 - ((2 * i) + 1)) * 6) + 1];
				end
				genvar _gv_i_53;
				for (_gv_i_53 = 0; _gv_i_53 < 8; _gv_i_53 = _gv_i_53 + 1) begin : gen_bitcnt_reg_in_b2
					localparam i = _gv_i_53;
					// Trace: design.sv:35032:9
					assign bitcnt_partial_msb_d[16 + i] = bitcnt_partial[((31 - ((4 * i) + 3)) * 6) + 2];
				end
				genvar _gv_i_54;
				for (_gv_i_54 = 0; _gv_i_54 < 4; _gv_i_54 = _gv_i_54 + 1) begin : gen_bitcnt_reg_in_b3
					localparam i = _gv_i_54;
					// Trace: design.sv:35036:9
					assign bitcnt_partial_msb_d[24 + i] = bitcnt_partial[((31 - ((8 * i) + 7)) * 6) + 3];
				end
				genvar _gv_i_55;
				for (_gv_i_55 = 0; _gv_i_55 < 2; _gv_i_55 = _gv_i_55 + 1) begin : gen_bitcnt_reg_in_b4
					localparam i = _gv_i_55;
					// Trace: design.sv:35040:9
					assign bitcnt_partial_msb_d[28 + i] = bitcnt_partial[((31 - ((16 * i) + 15)) * 6) + 4];
				end
				// Trace: design.sv:35043:7
				assign bitcnt_partial_msb_d[30] = bitcnt_partial[5];
				// Trace: design.sv:35044:7
				assign bitcnt_partial_msb_d[31] = 1'b0;
				// Trace: design.sv:35048:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:35049:9
					bitcnt_partial_q = {32 {6'b000000}};
					// Trace: design.sv:35051:9
					begin : sv2v_autoblock_11
						// Trace: design.sv:35051:14
						reg [31:0] i;
						// Trace: design.sv:35051:14
						for (i = 0; i < 32; i = i + 1)
							begin : gen_bitcnt_reg_out_lsb
								// Trace: design.sv:35052:11
								bitcnt_partial_q[(31 - i) * 6] = imd_val_q_i[32 + i];
							end
					end
					begin : sv2v_autoblock_12
						// Trace: design.sv:35055:14
						reg [31:0] i;
						// Trace: design.sv:35055:14
						for (i = 0; i < 16; i = i + 1)
							begin : gen_bitcnt_reg_out_b1
								// Trace: design.sv:35056:11
								bitcnt_partial_q[((31 - ((2 * i) + 1)) * 6) + 1] = imd_val_q_i[0 + i];
							end
					end
					begin : sv2v_autoblock_13
						// Trace: design.sv:35059:14
						reg [31:0] i;
						// Trace: design.sv:35059:14
						for (i = 0; i < 8; i = i + 1)
							begin : gen_bitcnt_reg_out_b2
								// Trace: design.sv:35060:11
								bitcnt_partial_q[((31 - ((4 * i) + 3)) * 6) + 2] = imd_val_q_i[16 + i];
							end
					end
					begin : sv2v_autoblock_14
						// Trace: design.sv:35063:14
						reg [31:0] i;
						// Trace: design.sv:35063:14
						for (i = 0; i < 4; i = i + 1)
							begin : gen_bitcnt_reg_out_b3
								// Trace: design.sv:35064:11
								bitcnt_partial_q[((31 - ((8 * i) + 7)) * 6) + 3] = imd_val_q_i[24 + i];
							end
					end
					begin : sv2v_autoblock_15
						// Trace: design.sv:35067:14
						reg [31:0] i;
						// Trace: design.sv:35067:14
						for (i = 0; i < 2; i = i + 1)
							begin : gen_bitcnt_reg_out_b4
								// Trace: design.sv:35068:11
								bitcnt_partial_q[((31 - ((16 * i) + 15)) * 6) + 4] = imd_val_q_i[28 + i];
							end
					end
					// Trace: design.sv:35071:9
					bitcnt_partial_q[5] = imd_val_q_i[30];
				end
				// Trace: design.sv:35074:7
				wire [31:0] butterfly_mask_l [0:4];
				// Trace: design.sv:35075:7
				wire [31:0] butterfly_mask_r [0:4];
				// Trace: design.sv:35076:7
				wire [31:0] butterfly_mask_not [0:4];
				// Trace: design.sv:35077:7
				wire [31:0] lrotc_stage [0:4];
				genvar _gv_stg_1;
				for (_gv_stg_1 = 0; _gv_stg_1 < 5; _gv_stg_1 = _gv_stg_1 + 1) begin : gen_butterfly_ctrl_stage
					localparam stg = _gv_stg_1;
					genvar _gv_seg_1;
					for (_gv_seg_1 = 0; _gv_seg_1 < (2 ** stg); _gv_seg_1 = _gv_seg_1 + 1) begin : gen_butterfly_ctrl
						localparam seg = _gv_seg_1;
						// Trace: design.sv:35087:11
						assign lrotc_stage[stg][((2 * (16 >> stg)) * (seg + 1)) - 1:(2 * (16 >> stg)) * seg] = {{16 >> stg {1'b0}}, {16 >> stg {1'b1}}} << bitcnt_partial_q[((32 - ((16 >> stg) * ((2 * seg) + 1))) * 6) + ($clog2(16 >> stg) >= 0 ? $clog2(16 >> stg) : ($clog2(16 >> stg) + ($clog2(16 >> stg) >= 0 ? $clog2(16 >> stg) + 1 : 1 - $clog2(16 >> stg))) - 1)-:($clog2(16 >> stg) >= 0 ? $clog2(16 >> stg) + 1 : 1 - $clog2(16 >> stg))];
						// Trace: design.sv:35091:11
						assign butterfly_mask_l[stg][((16 >> stg) * ((2 * seg) + 2)) - 1:(16 >> stg) * ((2 * seg) + 1)] = ~lrotc_stage[stg][((16 >> stg) * ((2 * seg) + 2)) - 1:(16 >> stg) * ((2 * seg) + 1)];
						// Trace: design.sv:35094:11
						assign butterfly_mask_r[stg][((16 >> stg) * ((2 * seg) + 1)) - 1:(16 >> stg) * (2 * seg)] = ~lrotc_stage[stg][((16 >> stg) * ((2 * seg) + 2)) - 1:(16 >> stg) * ((2 * seg) + 1)];
						// Trace: design.sv:35097:11
						assign butterfly_mask_l[stg][((16 >> stg) * ((2 * seg) + 1)) - 1:(16 >> stg) * (2 * seg)] = 1'sb0;
						// Trace: design.sv:35098:11
						assign butterfly_mask_r[stg][((16 >> stg) * ((2 * seg) + 2)) - 1:(16 >> stg) * ((2 * seg) + 1)] = 1'sb0;
					end
				end
				genvar _gv_stg_2;
				for (_gv_stg_2 = 0; _gv_stg_2 < 5; _gv_stg_2 = _gv_stg_2 + 1) begin : gen_butterfly_not
					localparam stg = _gv_stg_2;
					// Trace: design.sv:35104:9
					assign butterfly_mask_not[stg] = ~(butterfly_mask_l[stg] | butterfly_mask_r[stg]);
				end
				// Trace: design.sv:35108:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:35109:9
					butterfly_result = operand_a_i;
					// Trace: design.sv:35111:9
					butterfly_result = ((butterfly_result & butterfly_mask_not[0]) | ((butterfly_result & butterfly_mask_l[0]) >> 16)) | ((butterfly_result & butterfly_mask_r[0]) << 16);
					// Trace: design.sv:35115:9
					butterfly_result = ((butterfly_result & butterfly_mask_not[1]) | ((butterfly_result & butterfly_mask_l[1]) >> 8)) | ((butterfly_result & butterfly_mask_r[1]) << 8);
					// Trace: design.sv:35119:9
					butterfly_result = ((butterfly_result & butterfly_mask_not[2]) | ((butterfly_result & butterfly_mask_l[2]) >> 4)) | ((butterfly_result & butterfly_mask_r[2]) << 4);
					// Trace: design.sv:35123:9
					butterfly_result = ((butterfly_result & butterfly_mask_not[3]) | ((butterfly_result & butterfly_mask_l[3]) >> 2)) | ((butterfly_result & butterfly_mask_r[3]) << 2);
					// Trace: design.sv:35127:9
					butterfly_result = ((butterfly_result & butterfly_mask_not[4]) | ((butterfly_result & butterfly_mask_l[4]) >> 1)) | ((butterfly_result & butterfly_mask_r[4]) << 1);
					// Trace: design.sv:35131:9
					butterfly_result = butterfly_result & operand_b_i;
				end
				// Trace: design.sv:35134:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:35135:9
					invbutterfly_result = operand_a_i & operand_b_i;
					// Trace: design.sv:35137:9
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[4]) | ((invbutterfly_result & butterfly_mask_l[4]) >> 1)) | ((invbutterfly_result & butterfly_mask_r[4]) << 1);
					// Trace: design.sv:35141:9
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[3]) | ((invbutterfly_result & butterfly_mask_l[3]) >> 2)) | ((invbutterfly_result & butterfly_mask_r[3]) << 2);
					// Trace: design.sv:35145:9
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[2]) | ((invbutterfly_result & butterfly_mask_l[2]) >> 4)) | ((invbutterfly_result & butterfly_mask_r[2]) << 4);
					// Trace: design.sv:35149:9
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[1]) | ((invbutterfly_result & butterfly_mask_l[1]) >> 8)) | ((invbutterfly_result & butterfly_mask_r[1]) << 8);
					// Trace: design.sv:35153:9
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[0]) | ((invbutterfly_result & butterfly_mask_l[0]) >> 16)) | ((invbutterfly_result & butterfly_mask_r[0]) << 16);
				end
			end
			else begin : gen_alu_rvb_not_full
				// Trace: design.sv:35158:7
				wire [31:0] unused_imd_val_q_1;
				// Trace: design.sv:35159:7
				assign unused_imd_val_q_1 = imd_val_q_i[0+:32];
				// Trace: design.sv:35160:7
				wire [32:1] sv2v_tmp_98122;
				assign sv2v_tmp_98122 = 1'sb0;
				always @(*) butterfly_result = sv2v_tmp_98122;
				// Trace: design.sv:35161:7
				wire [32:1] sv2v_tmp_B39E0;
				assign sv2v_tmp_B39E0 = 1'sb0;
				always @(*) invbutterfly_result = sv2v_tmp_B39E0;
				// Trace: design.sv:35163:7
				assign bitcnt_partial_lsb_d = 1'sb0;
				// Trace: design.sv:35164:7
				assign bitcnt_partial_msb_d = 1'sb0;
			end
			// Trace: design.sv:35174:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:35175:7
				(* full_case, parallel_case *)
				case (operator_i)
					7'd45: begin
						// Trace: design.sv:35177:11
						multicycle_result = (operand_b_i == 32'h00000000 ? operand_a_i : imd_val_q_i[32+:32]);
						// Trace: design.sv:35178:11
						imd_val_d_o = {operand_a_i, 32'h00000000};
						// Trace: design.sv:35179:11
						if (instr_first_cycle_i)
							// Trace: design.sv:35180:13
							imd_val_we_o = 2'b01;
						else
							// Trace: design.sv:35182:13
							imd_val_we_o = 2'b00;
					end
					7'd46: begin
						// Trace: design.sv:35187:11
						multicycle_result = imd_val_q_i[32+:32] | bwlogic_and_result;
						// Trace: design.sv:35188:11
						imd_val_d_o = {bwlogic_and_result, 32'h00000000};
						// Trace: design.sv:35189:11
						if (instr_first_cycle_i)
							// Trace: design.sv:35190:13
							imd_val_we_o = 2'b01;
						else
							// Trace: design.sv:35192:13
							imd_val_we_o = 2'b00;
					end
					7'd48, 7'd47, 7'd14, 7'd13: begin
						// Trace: design.sv:35198:11
						if (shift_amt[4:0] == 5'h00)
							// Trace: design.sv:35199:13
							multicycle_result = (shift_amt[5] ? operand_a_i : imd_val_q_i[32+:32]);
						else
							// Trace: design.sv:35201:13
							multicycle_result = imd_val_q_i[32+:32] | shift_result;
						// Trace: design.sv:35203:11
						imd_val_d_o = {shift_result, 32'h00000000};
						if (instr_first_cycle_i)
							// Trace: design.sv:35205:13
							imd_val_we_o = 2'b01;
						else
							// Trace: design.sv:35207:13
							imd_val_we_o = 2'b00;
					end
					7'd63, 7'd64, 7'd61, 7'd62, 7'd59, 7'd60:
						// Trace: design.sv:35214:11
						if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
							// Trace: design.sv:35215:13
							(* full_case, parallel_case *)
							case (1'b1)
								crc_bmode:
									// Trace: design.sv:35216:26
									multicycle_result = clmul_result_rev ^ (operand_a_i >> 8);
								crc_hmode:
									// Trace: design.sv:35217:26
									multicycle_result = clmul_result_rev ^ (operand_a_i >> 16);
								default:
									// Trace: design.sv:35218:26
									multicycle_result = clmul_result_rev;
							endcase
							// Trace: design.sv:35220:13
							imd_val_d_o = {clmul_result_rev, 32'h00000000};
							if (instr_first_cycle_i)
								// Trace: design.sv:35222:15
								imd_val_we_o = 2'b01;
							else
								// Trace: design.sv:35224:15
								imd_val_we_o = 2'b00;
						end
						else begin
							// Trace: design.sv:35227:13
							imd_val_d_o = {operand_a_i, 32'h00000000};
							// Trace: design.sv:35228:13
							imd_val_we_o = 2'b00;
							// Trace: design.sv:35229:13
							multicycle_result = 1'sb0;
						end
					7'd53, 7'd54:
						// Trace: design.sv:35234:11
						if (RV32B == 32'sd3) begin
							// Trace: design.sv:35235:13
							multicycle_result = (operator_i == 7'd54 ? butterfly_result : invbutterfly_result);
							// Trace: design.sv:35237:13
							imd_val_d_o = {bitcnt_partial_lsb_d, bitcnt_partial_msb_d};
							// Trace: design.sv:35238:13
							if (instr_first_cycle_i)
								// Trace: design.sv:35239:15
								imd_val_we_o = 2'b11;
							else
								// Trace: design.sv:35241:15
								imd_val_we_o = 2'b00;
						end
						else begin
							// Trace: design.sv:35244:13
							imd_val_d_o = {operand_a_i, 32'h00000000};
							// Trace: design.sv:35245:13
							imd_val_we_o = 2'b00;
							// Trace: design.sv:35246:13
							multicycle_result = 1'sb0;
						end
					default: begin
						// Trace: design.sv:35251:11
						imd_val_d_o = {operand_a_i, 32'h00000000};
						// Trace: design.sv:35252:11
						imd_val_we_o = 2'b00;
						// Trace: design.sv:35253:11
						multicycle_result = 1'sb0;
					end
				endcase
			end
		end
		else begin : g_no_alu_rvb
			// Trace: design.sv:35260:5
			wire [63:0] unused_imd_val_q;
			// Trace: design.sv:35261:5
			assign unused_imd_val_q = imd_val_q_i;
			// Trace: design.sv:35262:5
			wire [31:0] unused_butterfly_result;
			// Trace: design.sv:35263:5
			assign unused_butterfly_result = butterfly_result;
			// Trace: design.sv:35264:5
			wire [31:0] unused_invbutterfly_result;
			// Trace: design.sv:35265:5
			assign unused_invbutterfly_result = invbutterfly_result;
			// Trace: design.sv:35267:5
			assign bitcnt_result = 1'sb0;
			// Trace: design.sv:35268:5
			assign minmax_result = 1'sb0;
			// Trace: design.sv:35269:5
			wire [32:1] sv2v_tmp_A0513;
			assign sv2v_tmp_A0513 = 1'sb0;
			always @(*) pack_result = sv2v_tmp_A0513;
			// Trace: design.sv:35270:5
			assign sext_result = 1'sb0;
			// Trace: design.sv:35271:5
			wire [32:1] sv2v_tmp_75CE4;
			assign sv2v_tmp_75CE4 = 1'sb0;
			always @(*) singlebit_result = sv2v_tmp_75CE4;
			// Trace: design.sv:35272:5
			wire [32:1] sv2v_tmp_FA09A;
			assign sv2v_tmp_FA09A = 1'sb0;
			always @(*) rev_result = sv2v_tmp_FA09A;
			// Trace: design.sv:35273:5
			wire [32:1] sv2v_tmp_4A308;
			assign sv2v_tmp_4A308 = 1'sb0;
			always @(*) shuffle_result = sv2v_tmp_4A308;
			// Trace: design.sv:35274:5
			assign xperm_result = 1'sb0;
			// Trace: design.sv:35275:5
			wire [32:1] sv2v_tmp_98122;
			assign sv2v_tmp_98122 = 1'sb0;
			always @(*) butterfly_result = sv2v_tmp_98122;
			// Trace: design.sv:35276:5
			wire [32:1] sv2v_tmp_B39E0;
			assign sv2v_tmp_B39E0 = 1'sb0;
			always @(*) invbutterfly_result = sv2v_tmp_B39E0;
			// Trace: design.sv:35277:5
			wire [32:1] sv2v_tmp_31DA6;
			assign sv2v_tmp_31DA6 = 1'sb0;
			always @(*) clmul_result = sv2v_tmp_31DA6;
			// Trace: design.sv:35278:5
			wire [32:1] sv2v_tmp_BC1B9;
			assign sv2v_tmp_BC1B9 = 1'sb0;
			always @(*) multicycle_result = sv2v_tmp_BC1B9;
			// Trace: design.sv:35280:5
			wire [64:1] sv2v_tmp_42A49;
			assign sv2v_tmp_42A49 = {2 {32'b00000000000000000000000000000000}};
			always @(*) imd_val_d_o = sv2v_tmp_42A49;
			// Trace: design.sv:35281:5
			wire [2:1] sv2v_tmp_0E15E;
			assign sv2v_tmp_0E15E = {2 {1'b0}};
			always @(*) imd_val_we_o = sv2v_tmp_0E15E;
		end
	endgenerate
	// Trace: design.sv:35288:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:35289:5
		result_o = 1'sb0;
		// Trace: design.sv:35291:5
		(* full_case, parallel_case *)
		case (operator_i)
			7'd2, 7'd5, 7'd3, 7'd6, 7'd4, 7'd7:
				// Trace: design.sv:35295:27
				result_o = bwlogic_result;
			7'd0, 7'd1, 7'd22, 7'd23, 7'd24:
				// Trace: design.sv:35301:19
				result_o = adder_result;
			7'd10, 7'd9, 7'd8, 7'd12, 7'd11:
				// Trace: design.sv:35307:26
				result_o = shift_result;
			7'd17, 7'd18:
				// Trace: design.sv:35310:29
				result_o = shuffle_result;
			7'd19, 7'd20, 7'd21:
				// Trace: design.sv:35313:46
				result_o = xperm_result;
			7'd29, 7'd30, 7'd27, 7'd28, 7'd25, 7'd26, 7'd43, 7'd44:
				// Trace: design.sv:35319:27
				result_o = {31'h00000000, cmp_result};
			7'd31, 7'd33, 7'd32, 7'd34:
				// Trace: design.sv:35323:27
				result_o = minmax_result;
			7'd40, 7'd41, 7'd42:
				// Trace: design.sv:35327:17
				result_o = {26'h0000000, bitcnt_result};
			7'd35, 7'd37, 7'd36:
				// Trace: design.sv:35331:18
				result_o = pack_result;
			7'd38, 7'd39:
				// Trace: design.sv:35334:29
				result_o = sext_result;
			7'd46, 7'd45, 7'd47, 7'd48, 7'd14, 7'd13, 7'd63, 7'd64, 7'd61, 7'd62, 7'd59, 7'd60, 7'd53, 7'd54:
				// Trace: design.sv:35346:39
				result_o = multicycle_result;
			7'd49, 7'd50, 7'd51, 7'd52:
				// Trace: design.sv:35350:27
				result_o = singlebit_result;
			7'd15, 7'd16:
				// Trace: design.sv:35353:27
				result_o = rev_result;
			7'd55:
				// Trace: design.sv:35356:16
				result_o = bfp_result;
			7'd56, 7'd57, 7'd58:
				// Trace: design.sv:35360:19
				result_o = clmul_result;
			default:
				;
		endcase
	end
	// Trace: design.sv:35366:3
	wire unused_shift_amt_compl;
	// Trace: design.sv:35367:3
	assign unused_shift_amt_compl = shift_amt_compl[5];
	initial _sv2v_0 = 0;
endmodule
module ibex_branch_predict (
	clk_i,
	rst_ni,
	fetch_rdata_i,
	fetch_pc_i,
	fetch_valid_i,
	predict_branch_taken_o,
	predict_branch_pc_o
);
	reg _sv2v_0;
	// Trace: design.sv:35390:3
	input wire clk_i;
	// Trace: design.sv:35391:3
	input wire rst_ni;
	// Trace: design.sv:35394:3
	input wire [31:0] fetch_rdata_i;
	// Trace: design.sv:35395:3
	input wire [31:0] fetch_pc_i;
	// Trace: design.sv:35396:3
	input wire fetch_valid_i;
	// Trace: design.sv:35399:3
	output wire predict_branch_taken_o;
	// Trace: design.sv:35400:3
	output wire [31:0] predict_branch_pc_o;
	// Trace: design.sv:35402:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:35404:3
	wire [31:0] imm_j_type;
	// Trace: design.sv:35405:3
	wire [31:0] imm_b_type;
	// Trace: design.sv:35406:3
	wire [31:0] imm_cj_type;
	// Trace: design.sv:35407:3
	wire [31:0] imm_cb_type;
	// Trace: design.sv:35409:3
	reg [31:0] branch_imm;
	// Trace: design.sv:35411:3
	wire [31:0] instr;
	// Trace: design.sv:35413:3
	wire instr_j;
	// Trace: design.sv:35414:3
	wire instr_b;
	// Trace: design.sv:35415:3
	wire instr_cj;
	// Trace: design.sv:35416:3
	wire instr_cb;
	// Trace: design.sv:35418:3
	wire instr_b_taken;
	// Trace: design.sv:35421:3
	assign instr = fetch_rdata_i;
	// Trace: design.sv:35427:3
	assign imm_j_type = {{12 {instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};
	// Trace: design.sv:35428:3
	assign imm_b_type = {{19 {instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
	// Trace: design.sv:35431:3
	assign imm_cj_type = {{20 {instr[12]}}, instr[12], instr[8], instr[10:9], instr[6], instr[7], instr[2], instr[11], instr[5:3], 1'b0};
	// Trace: design.sv:35434:3
	assign imm_cb_type = {{23 {instr[12]}}, instr[12], instr[6:5], instr[2], instr[11:10], instr[4:3], 1'b0};
	// Trace: design.sv:35440:3
	// removed localparam type ibex_pkg_opcode_e
	assign instr_b = instr[6:0] == 7'h63;
	// Trace: design.sv:35441:3
	assign instr_j = instr[6:0] == 7'h6f;
	// Trace: design.sv:35444:3
	assign instr_cb = (instr[1:0] == 2'b01) & ((instr[15:13] == 3'b110) | (instr[15:13] == 3'b111));
	// Trace: design.sv:35445:3
	assign instr_cj = (instr[1:0] == 2'b01) & ((instr[15:13] == 3'b101) | (instr[15:13] == 3'b001));
	// Trace: design.sv:35448:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:35449:5
		branch_imm = imm_b_type;
		// Trace: design.sv:35451:5
		(* full_case, parallel_case *)
		case (1'b1)
			instr_j:
				// Trace: design.sv:35452:18
				branch_imm = imm_j_type;
			instr_b:
				// Trace: design.sv:35453:18
				branch_imm = imm_b_type;
			instr_cj:
				// Trace: design.sv:35454:18
				branch_imm = imm_cj_type;
			instr_cb:
				// Trace: design.sv:35455:18
				branch_imm = imm_cb_type;
			default:
				;
		endcase
	end
	// Trace: design.sv:35463:3
	assign instr_b_taken = (instr_b & imm_b_type[31]) | (instr_cb & imm_cb_type[31]);
	// Trace: design.sv:35466:3
	assign predict_branch_taken_o = fetch_valid_i & ((instr_j | instr_cj) | instr_b_taken);
	// Trace: design.sv:35468:3
	assign predict_branch_pc_o = fetch_pc_i + branch_imm;
	initial _sv2v_0 = 0;
endmodule
module ibex_compressed_decoder (
	clk_i,
	rst_ni,
	valid_i,
	instr_i,
	instr_o,
	is_compressed_o,
	illegal_instr_o
);
	reg _sv2v_0;
	// Trace: design.sv:35486:3
	input wire clk_i;
	// Trace: design.sv:35487:3
	input wire rst_ni;
	// Trace: design.sv:35488:3
	input wire valid_i;
	// Trace: design.sv:35489:3
	input wire [31:0] instr_i;
	// Trace: design.sv:35490:3
	output reg [31:0] instr_o;
	// Trace: design.sv:35491:3
	output wire is_compressed_o;
	// Trace: design.sv:35492:3
	output reg illegal_instr_o;
	// Trace: design.sv:35494:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:35498:3
	wire unused_valid;
	// Trace: design.sv:35499:3
	assign unused_valid = valid_i;
	// Trace: design.sv:35505:3
	// removed localparam type ibex_pkg_opcode_e
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:35507:5
		instr_o = instr_i;
		// Trace: design.sv:35508:5
		illegal_instr_o = 1'b0;
		// Trace: design.sv:35511:5
		(* full_case, parallel_case *)
		case (instr_i[1:0])
			2'b00:
				// Trace: design.sv:35514:9
				(* full_case, parallel_case *)
				case (instr_i[15:13])
					3'b000: begin
						// Trace: design.sv:35517:13
						instr_o = {2'b00, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], 7'h13};
						// Trace: design.sv:35519:13
						if (instr_i[12:5] == 8'b00000000)
							// Trace: design.sv:35519:41
							illegal_instr_o = 1'b1;
					end
					3'b010:
						// Trace: design.sv:35524:13
						instr_o = {5'b00000, instr_i[5], instr_i[12:10], instr_i[6], 4'b0001, instr_i[9:7], 5'b01001, instr_i[4:2], 7'h03};
					3'b110:
						// Trace: design.sv:35530:13
						instr_o = {5'b00000, instr_i[5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b010, instr_i[11:10], instr_i[6], 9'h023};
					3'b001, 3'b011, 3'b100, 3'b101, 3'b111:
						// Trace: design.sv:35540:13
						illegal_instr_o = 1'b1;
					default:
						// Trace: design.sv:35544:13
						illegal_instr_o = 1'b1;
				endcase
			2'b01:
				// Trace: design.sv:35555:9
				(* full_case, parallel_case *)
				case (instr_i[15:13])
					3'b000:
						// Trace: design.sv:35559:13
						instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], 7'h13};
					3'b001, 3'b101:
						// Trace: design.sv:35566:13
						instr_o = {instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], {9 {instr_i[12]}}, 4'b0000, ~instr_i[15], 7'h6f};
					3'b010:
						// Trace: design.sv:35574:13
						instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 8'b00000000, instr_i[11:7], 7'h13};
					3'b011: begin
						// Trace: design.sv:35581:13
						instr_o = {{15 {instr_i[12]}}, instr_i[6:2], instr_i[11:7], 7'h37};
						// Trace: design.sv:35583:13
						if (instr_i[11:7] == 5'h02)
							// Trace: design.sv:35585:15
							instr_o = {{3 {instr_i[12]}}, instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 24'h010113};
						if ({instr_i[12], instr_i[6:2]} == 6'b000000)
							// Trace: design.sv:35589:54
							illegal_instr_o = 1'b1;
					end
					3'b100:
						// Trace: design.sv:35593:13
						(* full_case, parallel_case *)
						case (instr_i[11:10])
							2'b00, 2'b01: begin
								// Trace: design.sv:35599:17
								instr_o = {1'b0, instr_i[10], 5'b00000, instr_i[6:2], 2'b01, instr_i[9:7], 5'b10101, instr_i[9:7], 7'h13};
								// Trace: design.sv:35601:17
								if (instr_i[12] == 1'b1)
									// Trace: design.sv:35601:43
									illegal_instr_o = 1'b1;
							end
							2'b10:
								// Trace: design.sv:35606:17
								instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 2'b01, instr_i[9:7], 5'b11101, instr_i[9:7], 7'h13};
							2'b11:
								// Trace: design.sv:35611:17
								(* full_case, parallel_case *)
								case ({instr_i[12], instr_i[6:5]})
									3'b000:
										// Trace: design.sv:35614:21
										instr_o = {9'b010000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b00001, instr_i[9:7], 7'h33};
									3'b001:
										// Trace: design.sv:35620:21
										instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b10001, instr_i[9:7], 7'h33};
									3'b010:
										// Trace: design.sv:35626:21
										instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b11001, instr_i[9:7], 7'h33};
									3'b011:
										// Trace: design.sv:35632:21
										instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b11101, instr_i[9:7], 7'h33};
									3'b100, 3'b101, 3'b110, 3'b111:
										// Trace: design.sv:35642:21
										illegal_instr_o = 1'b1;
									default:
										// Trace: design.sv:35646:21
										illegal_instr_o = 1'b1;
								endcase
							default:
								// Trace: design.sv:35652:17
								illegal_instr_o = 1'b1;
						endcase
					3'b110, 3'b111:
						// Trace: design.sv:35660:13
						instr_o = {{4 {instr_i[12]}}, instr_i[6:5], instr_i[2], 7'b0000001, instr_i[9:7], 2'b00, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], 7'h63};
					default:
						// Trace: design.sv:35666:13
						illegal_instr_o = 1'b1;
				endcase
			2'b10:
				// Trace: design.sv:35677:9
				(* full_case, parallel_case *)
				case (instr_i[15:13])
					3'b000: begin
						// Trace: design.sv:35681:13
						instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b001, instr_i[11:7], 7'h13};
						// Trace: design.sv:35682:13
						if (instr_i[12] == 1'b1)
							// Trace: design.sv:35682:39
							illegal_instr_o = 1'b1;
					end
					3'b010: begin
						// Trace: design.sv:35687:13
						instr_o = {4'b0000, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], 7'h03};
						// Trace: design.sv:35689:13
						if (instr_i[11:7] == 5'b00000)
							// Trace: design.sv:35689:41
							illegal_instr_o = 1'b1;
					end
					3'b100:
						// Trace: design.sv:35693:13
						if (instr_i[12] == 1'b0) begin
							begin
								// Trace: design.sv:35694:15
								if (instr_i[6:2] != 5'b00000)
									// Trace: design.sv:35697:17
									instr_o = {7'b0000000, instr_i[6:2], 8'b00000000, instr_i[11:7], 7'h33};
								else begin
									// Trace: design.sv:35700:17
									instr_o = {12'b000000000000, instr_i[11:7], 15'h0067};
									// Trace: design.sv:35701:17
									if (instr_i[11:7] == 5'b00000)
										// Trace: design.sv:35701:44
										illegal_instr_o = 1'b1;
								end
							end
						end
						else
							// Trace: design.sv:35704:15
							if (instr_i[6:2] != 5'b00000)
								// Trace: design.sv:35707:17
								instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], 7'h33};
							else
								// Trace: design.sv:35709:17
								if (instr_i[11:7] == 5'b00000)
									// Trace: design.sv:35711:19
									instr_o = 32'h00100073;
								else
									// Trace: design.sv:35714:19
									instr_o = {12'b000000000000, instr_i[11:7], 15'h00e7};
					3'b110:
						// Trace: design.sv:35722:13
						instr_o = {4'b0000, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 9'h023};
					3'b001, 3'b011, 3'b101, 3'b111:
						// Trace: design.sv:35730:13
						illegal_instr_o = 1'b1;
					default:
						// Trace: design.sv:35734:13
						illegal_instr_o = 1'b1;
				endcase
			2'b11:
				;
			default:
				// Trace: design.sv:35743:9
				illegal_instr_o = 1'b1;
		endcase
	end
	// Trace: design.sv:35748:3
	assign is_compressed_o = instr_i[1:0] != 2'b11;
	initial _sv2v_0 = 0;
endmodule
module ibex_controller (
	clk_i,
	rst_ni,
	ctrl_busy_o,
	illegal_insn_i,
	ecall_insn_i,
	mret_insn_i,
	dret_insn_i,
	wfi_insn_i,
	ebrk_insn_i,
	csr_pipe_flush_i,
	instr_valid_i,
	instr_i,
	instr_compressed_i,
	instr_is_compressed_i,
	instr_bp_taken_i,
	instr_fetch_err_i,
	instr_fetch_err_plus2_i,
	pc_id_i,
	instr_valid_clear_o,
	id_in_ready_o,
	controller_run_o,
	instr_req_o,
	pc_set_o,
	pc_mux_o,
	nt_branch_mispredict_o,
	exc_pc_mux_o,
	exc_cause_o,
	lsu_addr_last_i,
	load_err_i,
	store_err_i,
	wb_exception_o,
	id_exception_o,
	branch_set_i,
	branch_not_set_i,
	jump_set_i,
	csr_mstatus_mie_i,
	irq_pending_i,
	irqs_i,
	irq_nm_i,
	nmi_mode_o,
	debug_req_i,
	debug_cause_o,
	debug_csr_save_o,
	debug_mode_o,
	debug_single_step_i,
	debug_ebreakm_i,
	debug_ebreaku_i,
	trigger_match_i,
	wake_from_sleep_o,
	csr_save_if_o,
	csr_save_id_o,
	csr_save_wb_o,
	csr_restore_mret_id_o,
	csr_restore_dret_id_o,
	csr_save_cause_o,
	csr_mtval_o,
	priv_mode_i,
	csr_mstatus_tw_i,
	stall_id_i,
	stall_wb_i,
	flush_id_o,
	ready_wb_i,
	perf_jump_o,
	perf_tbranch_o
);
	reg _sv2v_0;
	// Trace: design.sv:35786:13
	parameter [0:0] WritebackStage = 0;
	// Trace: design.sv:35787:13
	parameter [0:0] BranchPredictor = 0;
	// Trace: design.sv:35789:3
	input wire clk_i;
	// Trace: design.sv:35790:3
	input wire rst_ni;
	// Trace: design.sv:35792:3
	output reg ctrl_busy_o;
	// Trace: design.sv:35795:3
	input wire illegal_insn_i;
	// Trace: design.sv:35796:3
	input wire ecall_insn_i;
	// Trace: design.sv:35797:3
	input wire mret_insn_i;
	// Trace: design.sv:35798:3
	input wire dret_insn_i;
	// Trace: design.sv:35799:3
	input wire wfi_insn_i;
	// Trace: design.sv:35800:3
	input wire ebrk_insn_i;
	// Trace: design.sv:35801:3
	input wire csr_pipe_flush_i;
	// Trace: design.sv:35804:3
	input wire instr_valid_i;
	// Trace: design.sv:35805:3
	input wire [31:0] instr_i;
	// Trace: design.sv:35806:3
	input wire [15:0] instr_compressed_i;
	// Trace: design.sv:35807:3
	input wire instr_is_compressed_i;
	// Trace: design.sv:35808:3
	input wire instr_bp_taken_i;
	// Trace: design.sv:35809:3
	input wire instr_fetch_err_i;
	// Trace: design.sv:35810:3
	input wire instr_fetch_err_plus2_i;
	// Trace: design.sv:35811:3
	input wire [31:0] pc_id_i;
	// Trace: design.sv:35814:3
	output wire instr_valid_clear_o;
	// Trace: design.sv:35815:3
	output wire id_in_ready_o;
	// Trace: design.sv:35816:3
	output reg controller_run_o;
	// Trace: design.sv:35820:3
	output reg instr_req_o;
	// Trace: design.sv:35821:3
	output reg pc_set_o;
	// Trace: design.sv:35822:3
	// removed localparam type ibex_pkg_pc_sel_e
	output reg [2:0] pc_mux_o;
	// Trace: design.sv:35824:3
	output reg nt_branch_mispredict_o;
	// Trace: design.sv:35826:3
	// removed localparam type ibex_pkg_exc_pc_sel_e
	output reg [1:0] exc_pc_mux_o;
	// Trace: design.sv:35827:3
	// removed localparam type ibex_pkg_exc_cause_e
	output reg [5:0] exc_cause_o;
	// Trace: design.sv:35830:3
	input wire [31:0] lsu_addr_last_i;
	// Trace: design.sv:35831:3
	input wire load_err_i;
	// Trace: design.sv:35832:3
	input wire store_err_i;
	// Trace: design.sv:35833:3
	output wire wb_exception_o;
	// Trace: design.sv:35834:3
	output wire id_exception_o;
	// Trace: design.sv:35837:3
	input wire branch_set_i;
	// Trace: design.sv:35839:3
	input wire branch_not_set_i;
	// Trace: design.sv:35840:3
	input wire jump_set_i;
	// Trace: design.sv:35843:3
	input wire csr_mstatus_mie_i;
	// Trace: design.sv:35844:3
	input wire irq_pending_i;
	// Trace: design.sv:35845:3
	// removed localparam type ibex_pkg_irqs_t
	input wire [17:0] irqs_i;
	// Trace: design.sv:35847:3
	input wire irq_nm_i;
	// Trace: design.sv:35848:3
	output wire nmi_mode_o;
	// Trace: design.sv:35851:3
	input wire debug_req_i;
	// Trace: design.sv:35852:3
	// removed localparam type ibex_pkg_dbg_cause_e
	output reg [2:0] debug_cause_o;
	// Trace: design.sv:35853:3
	output reg debug_csr_save_o;
	// Trace: design.sv:35854:3
	output wire debug_mode_o;
	// Trace: design.sv:35855:3
	input wire debug_single_step_i;
	// Trace: design.sv:35856:3
	input wire debug_ebreakm_i;
	// Trace: design.sv:35857:3
	input wire debug_ebreaku_i;
	// Trace: design.sv:35858:3
	input wire trigger_match_i;
	// Trace: design.sv:35861:3
	output wire wake_from_sleep_o;
	// Trace: design.sv:35863:3
	output reg csr_save_if_o;
	// Trace: design.sv:35864:3
	output reg csr_save_id_o;
	// Trace: design.sv:35865:3
	output reg csr_save_wb_o;
	// Trace: design.sv:35866:3
	output reg csr_restore_mret_id_o;
	// Trace: design.sv:35867:3
	output reg csr_restore_dret_id_o;
	// Trace: design.sv:35868:3
	output reg csr_save_cause_o;
	// Trace: design.sv:35869:3
	output reg [31:0] csr_mtval_o;
	// Trace: design.sv:35870:3
	// removed localparam type ibex_pkg_priv_lvl_e
	input wire [1:0] priv_mode_i;
	// Trace: design.sv:35871:3
	input wire csr_mstatus_tw_i;
	// Trace: design.sv:35874:3
	input wire stall_id_i;
	// Trace: design.sv:35875:3
	input wire stall_wb_i;
	// Trace: design.sv:35876:3
	output wire flush_id_o;
	// Trace: design.sv:35877:3
	input wire ready_wb_i;
	// Trace: design.sv:35880:3
	output reg perf_jump_o;
	// Trace: design.sv:35882:3
	output reg perf_tbranch_o;
	// Trace: design.sv:35885:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:35888:3
	// removed localparam type ctrl_fsm_e
	// Trace: design.sv:35893:3
	reg [3:0] ctrl_fsm_cs;
	reg [3:0] ctrl_fsm_ns;
	// Trace: design.sv:35895:3
	reg nmi_mode_q;
	reg nmi_mode_d;
	// Trace: design.sv:35896:3
	reg debug_mode_q;
	reg debug_mode_d;
	// Trace: design.sv:35897:3
	reg load_err_q;
	wire load_err_d;
	// Trace: design.sv:35898:3
	reg store_err_q;
	wire store_err_d;
	// Trace: design.sv:35899:3
	reg exc_req_q;
	wire exc_req_d;
	// Trace: design.sv:35900:3
	reg illegal_insn_q;
	wire illegal_insn_d;
	// Trace: design.sv:35904:3
	reg instr_fetch_err_prio;
	// Trace: design.sv:35905:3
	reg illegal_insn_prio;
	// Trace: design.sv:35906:3
	reg ecall_insn_prio;
	// Trace: design.sv:35907:3
	reg ebrk_insn_prio;
	// Trace: design.sv:35908:3
	reg store_err_prio;
	// Trace: design.sv:35909:3
	reg load_err_prio;
	// Trace: design.sv:35911:3
	wire stall;
	// Trace: design.sv:35912:3
	reg halt_if;
	// Trace: design.sv:35913:3
	reg retain_id;
	// Trace: design.sv:35914:3
	reg flush_id;
	// Trace: design.sv:35915:3
	wire illegal_dret;
	// Trace: design.sv:35916:3
	wire illegal_umode;
	// Trace: design.sv:35917:3
	wire exc_req_lsu;
	// Trace: design.sv:35918:3
	wire special_req;
	// Trace: design.sv:35919:3
	wire special_req_pc_change;
	// Trace: design.sv:35920:3
	wire special_req_flush_only;
	// Trace: design.sv:35921:3
	wire do_single_step_d;
	// Trace: design.sv:35922:3
	reg do_single_step_q;
	// Trace: design.sv:35923:3
	wire enter_debug_mode_prio_d;
	// Trace: design.sv:35924:3
	reg enter_debug_mode_prio_q;
	// Trace: design.sv:35925:3
	wire enter_debug_mode;
	// Trace: design.sv:35926:3
	wire ebreak_into_debug;
	// Trace: design.sv:35927:3
	wire handle_irq;
	// Trace: design.sv:35928:3
	wire id_wb_pending;
	// Trace: design.sv:35930:3
	reg [3:0] mfip_id;
	// Trace: design.sv:35931:3
	wire unused_irq_timer;
	// Trace: design.sv:35933:3
	wire ecall_insn;
	// Trace: design.sv:35934:3
	wire mret_insn;
	// Trace: design.sv:35935:3
	wire dret_insn;
	// Trace: design.sv:35936:3
	wire wfi_insn;
	// Trace: design.sv:35937:3
	wire ebrk_insn;
	// Trace: design.sv:35938:3
	wire csr_pipe_flush;
	// Trace: design.sv:35939:3
	wire instr_fetch_err;
	// Trace: design.sv:35959:3
	assign load_err_d = load_err_i;
	// Trace: design.sv:35960:3
	assign store_err_d = store_err_i;
	// Trace: design.sv:35963:3
	assign ecall_insn = ecall_insn_i & instr_valid_i;
	// Trace: design.sv:35964:3
	assign mret_insn = mret_insn_i & instr_valid_i;
	// Trace: design.sv:35965:3
	assign dret_insn = dret_insn_i & instr_valid_i;
	// Trace: design.sv:35966:3
	assign wfi_insn = wfi_insn_i & instr_valid_i;
	// Trace: design.sv:35967:3
	assign ebrk_insn = ebrk_insn_i & instr_valid_i;
	// Trace: design.sv:35968:3
	assign csr_pipe_flush = csr_pipe_flush_i & instr_valid_i;
	// Trace: design.sv:35969:3
	assign instr_fetch_err = instr_fetch_err_i & instr_valid_i;
	// Trace: design.sv:35973:3
	assign illegal_dret = dret_insn & ~debug_mode_q;
	// Trace: design.sv:35976:3
	assign illegal_umode = (priv_mode_i != 2'b11) & (mret_insn | (csr_mstatus_tw_i & wfi_insn));
	// Trace: design.sv:35985:3
	assign illegal_insn_d = ((illegal_insn_i | illegal_dret) | illegal_umode) & (ctrl_fsm_cs != 4'd6);
	// Trace: design.sv:35992:3
	assign exc_req_d = (((ecall_insn | ebrk_insn) | illegal_insn_d) | instr_fetch_err) & (ctrl_fsm_cs != 4'd6);
	// Trace: design.sv:35996:3
	assign exc_req_lsu = store_err_i | load_err_i;
	// Trace: design.sv:35998:3
	assign id_exception_o = exc_req_d;
	// Trace: design.sv:36006:3
	assign special_req_flush_only = wfi_insn | csr_pipe_flush;
	// Trace: design.sv:36009:3
	assign special_req_pc_change = ((mret_insn | dret_insn) | exc_req_d) | exc_req_lsu;
	// Trace: design.sv:36012:3
	assign special_req = special_req_pc_change | special_req_flush_only;
	// Trace: design.sv:36015:3
	assign id_wb_pending = instr_valid_i | ~ready_wb_i;
	// Trace: design.sv:36018:3
	generate
		if (WritebackStage) begin : g_wb_exceptions
			// Trace: design.sv:36019:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:36020:7
				instr_fetch_err_prio = 0;
				// Trace: design.sv:36021:7
				illegal_insn_prio = 0;
				// Trace: design.sv:36022:7
				ecall_insn_prio = 0;
				// Trace: design.sv:36023:7
				ebrk_insn_prio = 0;
				// Trace: design.sv:36024:7
				store_err_prio = 0;
				// Trace: design.sv:36025:7
				load_err_prio = 0;
				// Trace: design.sv:36030:7
				if (store_err_q)
					// Trace: design.sv:36031:9
					store_err_prio = 1'b1;
				else if (load_err_q)
					// Trace: design.sv:36033:9
					load_err_prio = 1'b1;
				else if (instr_fetch_err)
					// Trace: design.sv:36035:9
					instr_fetch_err_prio = 1'b1;
				else if (illegal_insn_q)
					// Trace: design.sv:36037:9
					illegal_insn_prio = 1'b1;
				else if (ecall_insn)
					// Trace: design.sv:36039:9
					ecall_insn_prio = 1'b1;
				else if (ebrk_insn)
					// Trace: design.sv:36041:9
					ebrk_insn_prio = 1'b1;
			end
			// Trace: design.sv:36046:5
			assign wb_exception_o = ((load_err_q | store_err_q) | load_err_i) | store_err_i;
		end
		else begin : g_no_wb_exceptions
			// Trace: design.sv:36048:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:36049:7
				instr_fetch_err_prio = 0;
				// Trace: design.sv:36050:7
				illegal_insn_prio = 0;
				// Trace: design.sv:36051:7
				ecall_insn_prio = 0;
				// Trace: design.sv:36052:7
				ebrk_insn_prio = 0;
				// Trace: design.sv:36053:7
				store_err_prio = 0;
				// Trace: design.sv:36054:7
				load_err_prio = 0;
				// Trace: design.sv:36056:7
				if (instr_fetch_err)
					// Trace: design.sv:36057:9
					instr_fetch_err_prio = 1'b1;
				else if (illegal_insn_q)
					// Trace: design.sv:36059:9
					illegal_insn_prio = 1'b1;
				else if (ecall_insn)
					// Trace: design.sv:36061:9
					ecall_insn_prio = 1'b1;
				else if (ebrk_insn)
					// Trace: design.sv:36063:9
					ebrk_insn_prio = 1'b1;
				else if (store_err_q)
					// Trace: design.sv:36065:9
					store_err_prio = 1'b1;
				else if (load_err_q)
					// Trace: design.sv:36067:9
					load_err_prio = 1'b1;
			end
			// Trace: design.sv:36070:5
			assign wb_exception_o = 1'b0;
		end
	endgenerate
	// Trace: design.sv:36097:3
	assign do_single_step_d = (instr_valid_i ? ~debug_mode_q & debug_single_step_i : do_single_step_q);
	// Trace: design.sv:36108:3
	assign enter_debug_mode_prio_d = (debug_req_i | do_single_step_d) & ~debug_mode_q;
	// Trace: design.sv:36109:3
	assign enter_debug_mode = enter_debug_mode_prio_d | (trigger_match_i & ~debug_mode_q);
	// Trace: design.sv:36113:3
	assign ebreak_into_debug = (priv_mode_i == 2'b11 ? debug_ebreakm_i : (priv_mode_i == 2'b00 ? debug_ebreaku_i : 1'b0));
	// Trace: design.sv:36121:3
	assign handle_irq = (~debug_mode_q & ~nmi_mode_q) & (irq_nm_i | (irq_pending_i & csr_mstatus_mie_i));
	// Trace: design.sv:36125:3
	always @(*) begin : gen_mfip_id
		if (_sv2v_0)
			;
		// Trace: design.sv:36126:5
		mfip_id = 4'd0;
		// Trace: design.sv:36128:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:36128:10
			reg signed [31:0] i;
			// Trace: design.sv:36128:10
			for (i = 14; i >= 0; i = i - 1)
				begin
					// Trace: design.sv:36129:7
					if (irqs_i[0 + i])
						// Trace: design.sv:36130:9
						mfip_id = i[3:0];
				end
		end
	end
	// Trace: design.sv:36135:3
	assign unused_irq_timer = irqs_i[16];
	// Trace: design.sv:36141:3
	function automatic [5:0] sv2v_cast_6;
		input reg [5:0] inp;
		sv2v_cast_6 = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:36143:5
		instr_req_o = 1'b1;
		// Trace: design.sv:36145:5
		csr_save_if_o = 1'b0;
		// Trace: design.sv:36146:5
		csr_save_id_o = 1'b0;
		// Trace: design.sv:36147:5
		csr_save_wb_o = 1'b0;
		// Trace: design.sv:36148:5
		csr_restore_mret_id_o = 1'b0;
		// Trace: design.sv:36149:5
		csr_restore_dret_id_o = 1'b0;
		// Trace: design.sv:36150:5
		csr_save_cause_o = 1'b0;
		// Trace: design.sv:36151:5
		csr_mtval_o = 1'sb0;
		// Trace: design.sv:36157:5
		pc_mux_o = 3'd0;
		// Trace: design.sv:36158:5
		pc_set_o = 1'b0;
		// Trace: design.sv:36159:5
		nt_branch_mispredict_o = 1'b0;
		// Trace: design.sv:36161:5
		exc_pc_mux_o = 2'd1;
		// Trace: design.sv:36162:5
		exc_cause_o = 6'h00;
		// Trace: design.sv:36164:5
		ctrl_fsm_ns = ctrl_fsm_cs;
		// Trace: design.sv:36166:5
		ctrl_busy_o = 1'b1;
		// Trace: design.sv:36168:5
		halt_if = 1'b0;
		// Trace: design.sv:36169:5
		retain_id = 1'b0;
		// Trace: design.sv:36170:5
		flush_id = 1'b0;
		// Trace: design.sv:36172:5
		debug_csr_save_o = 1'b0;
		// Trace: design.sv:36173:5
		debug_cause_o = 3'h1;
		// Trace: design.sv:36174:5
		debug_mode_d = debug_mode_q;
		// Trace: design.sv:36175:5
		nmi_mode_d = nmi_mode_q;
		// Trace: design.sv:36177:5
		perf_tbranch_o = 1'b0;
		// Trace: design.sv:36178:5
		perf_jump_o = 1'b0;
		// Trace: design.sv:36180:5
		controller_run_o = 1'b0;
		// Trace: design.sv:36182:5
		(* full_case, parallel_case *)
		case (ctrl_fsm_cs)
			4'd0: begin
				// Trace: design.sv:36184:9
				instr_req_o = 1'b0;
				// Trace: design.sv:36185:9
				pc_mux_o = 3'd0;
				// Trace: design.sv:36186:9
				pc_set_o = 1'b1;
				// Trace: design.sv:36187:9
				ctrl_fsm_ns = 4'd1;
			end
			4'd1: begin
				// Trace: design.sv:36192:9
				instr_req_o = 1'b1;
				// Trace: design.sv:36193:9
				pc_mux_o = 3'd0;
				// Trace: design.sv:36194:9
				pc_set_o = 1'b1;
				// Trace: design.sv:36196:9
				ctrl_fsm_ns = 4'd4;
			end
			4'd2: begin
				// Trace: design.sv:36200:9
				ctrl_busy_o = 1'b0;
				// Trace: design.sv:36201:9
				instr_req_o = 1'b0;
				// Trace: design.sv:36202:9
				halt_if = 1'b1;
				// Trace: design.sv:36203:9
				flush_id = 1'b1;
				// Trace: design.sv:36204:9
				ctrl_fsm_ns = 4'd3;
			end
			4'd3: begin
				// Trace: design.sv:36210:9
				instr_req_o = 1'b0;
				// Trace: design.sv:36211:9
				halt_if = 1'b1;
				// Trace: design.sv:36212:9
				flush_id = 1'b1;
				// Trace: design.sv:36216:9
				if (wake_from_sleep_o)
					// Trace: design.sv:36217:11
					ctrl_fsm_ns = 4'd4;
				else
					// Trace: design.sv:36220:11
					ctrl_busy_o = 1'b0;
			end
			4'd4: begin
				// Trace: design.sv:36227:9
				if (id_in_ready_o)
					// Trace: design.sv:36228:11
					ctrl_fsm_ns = 4'd5;
				if (handle_irq) begin
					// Trace: design.sv:36237:11
					ctrl_fsm_ns = 4'd7;
					// Trace: design.sv:36238:11
					halt_if = 1'b1;
				end
				if (enter_debug_mode) begin
					// Trace: design.sv:36243:11
					ctrl_fsm_ns = 4'd8;
					// Trace: design.sv:36246:11
					halt_if = 1'b1;
				end
			end
			4'd5: begin
				// Trace: design.sv:36257:9
				controller_run_o = 1'b1;
				// Trace: design.sv:36262:9
				pc_mux_o = 3'd1;
				// Trace: design.sv:36266:9
				if (special_req) begin
					// Trace: design.sv:36270:11
					retain_id = 1'b1;
					// Trace: design.sv:36278:11
					if (ready_wb_i | wb_exception_o)
						// Trace: design.sv:36279:13
						ctrl_fsm_ns = 4'd6;
				end
				if (branch_set_i || jump_set_i) begin
					// Trace: design.sv:36285:11
					pc_set_o = (BranchPredictor ? ~instr_bp_taken_i : 1'b1);
					// Trace: design.sv:36287:11
					perf_tbranch_o = branch_set_i;
					// Trace: design.sv:36288:11
					perf_jump_o = jump_set_i;
				end
				if (BranchPredictor) begin
					begin
						// Trace: design.sv:36292:11
						if (instr_bp_taken_i & branch_not_set_i)
							// Trace: design.sv:36295:13
							nt_branch_mispredict_o = 1'b1;
					end
				end
				if ((enter_debug_mode || handle_irq) && (stall || id_wb_pending))
					// Trace: design.sv:36302:11
					halt_if = 1'b1;
				if ((!stall && !special_req) && !id_wb_pending) begin
					begin
						// Trace: design.sv:36306:11
						if (enter_debug_mode) begin
							// Trace: design.sv:36308:13
							ctrl_fsm_ns = 4'd8;
							// Trace: design.sv:36311:13
							halt_if = 1'b1;
						end
						else if (handle_irq) begin
							// Trace: design.sv:36314:13
							ctrl_fsm_ns = 4'd7;
							// Trace: design.sv:36320:13
							halt_if = 1'b1;
						end
					end
				end
			end
			4'd7: begin
				// Trace: design.sv:36327:9
				pc_mux_o = 3'd2;
				// Trace: design.sv:36328:9
				exc_pc_mux_o = 2'd1;
				// Trace: design.sv:36330:9
				if (handle_irq) begin
					// Trace: design.sv:36331:11
					pc_set_o = 1'b1;
					// Trace: design.sv:36333:11
					csr_save_if_o = 1'b1;
					// Trace: design.sv:36334:11
					csr_save_cause_o = 1'b1;
					// Trace: design.sv:36337:11
					if (irq_nm_i && !nmi_mode_q) begin
						// Trace: design.sv:36338:13
						exc_cause_o = 6'h3f;
						// Trace: design.sv:36339:13
						nmi_mode_d = 1'b1;
					end
					else if (irqs_i[14-:15] != 15'b000000000000000)
						// Trace: design.sv:36345:13
						exc_cause_o = sv2v_cast_6({2'b11, mfip_id});
					else if (irqs_i[15])
						// Trace: design.sv:36347:13
						exc_cause_o = 6'h2b;
					else if (irqs_i[17])
						// Trace: design.sv:36349:13
						exc_cause_o = 6'h23;
					else
						// Trace: design.sv:36351:13
						exc_cause_o = 6'h27;
				end
				// Trace: design.sv:36355:9
				ctrl_fsm_ns = 4'd5;
			end
			4'd8: begin
				// Trace: design.sv:36359:9
				pc_mux_o = 3'd2;
				// Trace: design.sv:36360:9
				exc_pc_mux_o = 2'd2;
				// Trace: design.sv:36364:9
				flush_id = 1'b1;
				// Trace: design.sv:36365:9
				pc_set_o = 1'b1;
				// Trace: design.sv:36367:9
				csr_save_if_o = 1'b1;
				// Trace: design.sv:36368:9
				debug_csr_save_o = 1'b1;
				// Trace: design.sv:36370:9
				csr_save_cause_o = 1'b1;
				// Trace: design.sv:36371:9
				if (trigger_match_i)
					// Trace: design.sv:36372:11
					debug_cause_o = 3'h2;
				else if (debug_single_step_i)
					// Trace: design.sv:36374:11
					debug_cause_o = 3'h4;
				else
					// Trace: design.sv:36376:11
					debug_cause_o = 3'h3;
				// Trace: design.sv:36380:9
				debug_mode_d = 1'b1;
				// Trace: design.sv:36382:9
				ctrl_fsm_ns = 4'd5;
			end
			4'd9: begin
				// Trace: design.sv:36393:9
				flush_id = 1'b1;
				// Trace: design.sv:36394:9
				pc_mux_o = 3'd2;
				// Trace: design.sv:36395:9
				pc_set_o = 1'b1;
				// Trace: design.sv:36396:9
				exc_pc_mux_o = 2'd2;
				// Trace: design.sv:36399:9
				if (ebreak_into_debug && !debug_mode_q) begin
					// Trace: design.sv:36402:11
					csr_save_cause_o = 1'b1;
					// Trace: design.sv:36403:11
					csr_save_id_o = 1'b1;
					// Trace: design.sv:36406:11
					debug_csr_save_o = 1'b1;
					// Trace: design.sv:36407:11
					debug_cause_o = 3'h1;
				end
				// Trace: design.sv:36411:9
				debug_mode_d = 1'b1;
				// Trace: design.sv:36413:9
				ctrl_fsm_ns = 4'd5;
			end
			4'd6: begin
				// Trace: design.sv:36418:9
				halt_if = 1'b1;
				// Trace: design.sv:36419:9
				flush_id = 1'b1;
				// Trace: design.sv:36420:9
				ctrl_fsm_ns = 4'd5;
				// Trace: design.sv:36427:9
				if ((exc_req_q || store_err_q) || load_err_q) begin
					// Trace: design.sv:36428:11
					pc_set_o = 1'b1;
					// Trace: design.sv:36429:11
					pc_mux_o = 3'd2;
					// Trace: design.sv:36430:11
					exc_pc_mux_o = (debug_mode_q ? 2'd3 : 2'd0);
					// Trace: design.sv:36432:11
					if (WritebackStage) begin : g_writeback_mepc_save
						// Trace: design.sv:36436:13
						csr_save_id_o = ~(store_err_q | load_err_q);
						// Trace: design.sv:36437:13
						csr_save_wb_o = store_err_q | load_err_q;
					end
					else begin : g_no_writeback_mepc_save
						// Trace: design.sv:36439:13
						csr_save_id_o = 1'b0;
					end
					// Trace: design.sv:36442:11
					csr_save_cause_o = 1'b1;
					(* full_case, parallel_case *)
					case (1'b1)
						instr_fetch_err_prio: begin
							// Trace: design.sv:36447:15
							exc_cause_o = 6'h01;
							// Trace: design.sv:36448:15
							csr_mtval_o = (instr_fetch_err_plus2_i ? pc_id_i + 32'd2 : pc_id_i);
						end
						illegal_insn_prio: begin
							// Trace: design.sv:36451:15
							exc_cause_o = 6'h02;
							// Trace: design.sv:36452:15
							csr_mtval_o = (instr_is_compressed_i ? {16'b0000000000000000, instr_compressed_i} : instr_i);
						end
						ecall_insn_prio:
							// Trace: design.sv:36455:15
							exc_cause_o = (priv_mode_i == 2'b11 ? 6'h0b : 6'h08);
						ebrk_insn_prio:
							// Trace: design.sv:36459:15
							if (debug_mode_q | ebreak_into_debug) begin
								// Trace: design.sv:36473:17
								pc_set_o = 1'b0;
								// Trace: design.sv:36474:17
								csr_save_id_o = 1'b0;
								// Trace: design.sv:36475:17
								csr_save_cause_o = 1'b0;
								// Trace: design.sv:36476:17
								ctrl_fsm_ns = 4'd9;
								// Trace: design.sv:36477:17
								flush_id = 1'b0;
							end
							else
								// Trace: design.sv:36488:17
								exc_cause_o = 6'h03;
						store_err_prio: begin
							// Trace: design.sv:36492:15
							exc_cause_o = 6'h07;
							// Trace: design.sv:36493:15
							csr_mtval_o = lsu_addr_last_i;
						end
						load_err_prio: begin
							// Trace: design.sv:36496:15
							exc_cause_o = 6'h05;
							// Trace: design.sv:36497:15
							csr_mtval_o = lsu_addr_last_i;
						end
						default:
							;
					endcase
				end
				else
					// Trace: design.sv:36503:11
					if (mret_insn) begin
						// Trace: design.sv:36504:13
						pc_mux_o = 3'd3;
						// Trace: design.sv:36505:13
						pc_set_o = 1'b1;
						// Trace: design.sv:36506:13
						csr_restore_mret_id_o = 1'b1;
						// Trace: design.sv:36507:13
						if (nmi_mode_q)
							// Trace: design.sv:36508:15
							nmi_mode_d = 1'b0;
					end
					else if (dret_insn) begin
						// Trace: design.sv:36511:13
						pc_mux_o = 3'd4;
						// Trace: design.sv:36512:13
						pc_set_o = 1'b1;
						// Trace: design.sv:36513:13
						debug_mode_d = 1'b0;
						// Trace: design.sv:36514:13
						csr_restore_dret_id_o = 1'b1;
					end
					else if (wfi_insn)
						// Trace: design.sv:36516:13
						ctrl_fsm_ns = 4'd2;
					else if (csr_pipe_flush && handle_irq)
						// Trace: design.sv:36519:13
						ctrl_fsm_ns = 4'd7;
				if (enter_debug_mode_prio_q && !(ebrk_insn_prio && ebreak_into_debug))
					// Trace: design.sv:36533:11
					ctrl_fsm_ns = 4'd8;
			end
			default: begin
				// Trace: design.sv:36538:9
				instr_req_o = 1'b0;
				// Trace: design.sv:36539:9
				ctrl_fsm_ns = 4'd0;
			end
		endcase
	end
	// Trace: design.sv:36544:3
	assign flush_id_o = flush_id;
	// Trace: design.sv:36547:3
	assign debug_mode_o = debug_mode_q;
	// Trace: design.sv:36550:3
	assign nmi_mode_o = nmi_mode_q;
	// Trace: design.sv:36559:3
	assign stall = stall_id_i | stall_wb_i;
	// Trace: design.sv:36562:3
	assign id_in_ready_o = (~stall & ~halt_if) & ~retain_id;
	// Trace: design.sv:36569:3
	assign instr_valid_clear_o = ~(stall | retain_id) | flush_id;
	// Trace: design.sv:36572:3
	always @(posedge clk_i or negedge rst_ni) begin : update_regs
		// Trace: design.sv:36573:5
		if (!rst_ni) begin
			// Trace: design.sv:36574:7
			ctrl_fsm_cs <= 4'd0;
			// Trace: design.sv:36575:7
			nmi_mode_q <= 1'b0;
			// Trace: design.sv:36576:7
			do_single_step_q <= 1'b0;
			// Trace: design.sv:36577:7
			debug_mode_q <= 1'b0;
			// Trace: design.sv:36578:7
			enter_debug_mode_prio_q <= 1'b0;
			// Trace: design.sv:36579:7
			load_err_q <= 1'b0;
			// Trace: design.sv:36580:7
			store_err_q <= 1'b0;
			// Trace: design.sv:36581:7
			exc_req_q <= 1'b0;
			// Trace: design.sv:36582:7
			illegal_insn_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:36584:7
			ctrl_fsm_cs <= ctrl_fsm_ns;
			// Trace: design.sv:36585:7
			nmi_mode_q <= nmi_mode_d;
			// Trace: design.sv:36586:7
			do_single_step_q <= do_single_step_d;
			// Trace: design.sv:36587:7
			debug_mode_q <= debug_mode_d;
			// Trace: design.sv:36588:7
			enter_debug_mode_prio_q <= enter_debug_mode_prio_d;
			// Trace: design.sv:36589:7
			load_err_q <= load_err_d;
			// Trace: design.sv:36590:7
			store_err_q <= store_err_d;
			// Trace: design.sv:36591:7
			exc_req_q <= exc_req_d;
			// Trace: design.sv:36592:7
			illegal_insn_q <= illegal_insn_d;
		end
	end
	// Trace: design.sv:36596:3
	assign wake_from_sleep_o = (((irq_nm_i || irq_pending_i) || debug_req_i) || debug_mode_q) || debug_single_step_i;
	initial _sv2v_0 = 0;
endmodule
module ibex_cs_registers (
	clk_i,
	rst_ni,
	hart_id_i,
	priv_mode_id_o,
	priv_mode_lsu_o,
	csr_mstatus_tw_o,
	csr_mtvec_o,
	csr_mtvec_init_i,
	boot_addr_i,
	csr_access_i,
	csr_addr_i,
	csr_wdata_i,
	csr_op_i,
	csr_op_en_i,
	csr_rdata_o,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	irq_fast_i,
	nmi_mode_i,
	irq_pending_o,
	irqs_o,
	csr_mstatus_mie_o,
	csr_mepc_o,
	csr_pmp_cfg_o,
	csr_pmp_addr_o,
	csr_pmp_mseccfg_o,
	debug_mode_i,
	debug_cause_i,
	debug_csr_save_i,
	csr_depc_o,
	debug_single_step_o,
	debug_ebreakm_o,
	debug_ebreaku_o,
	trigger_match_o,
	pc_if_i,
	pc_id_i,
	pc_wb_i,
	data_ind_timing_o,
	dummy_instr_en_o,
	dummy_instr_mask_o,
	dummy_instr_seed_en_o,
	dummy_instr_seed_o,
	icache_enable_o,
	csr_shadow_err_o,
	csr_save_if_i,
	csr_save_id_i,
	csr_save_wb_i,
	csr_restore_mret_i,
	csr_restore_dret_i,
	csr_save_cause_i,
	csr_mcause_i,
	csr_mtval_i,
	illegal_csr_insn_o,
	double_fault_seen_o,
	instr_ret_i,
	instr_ret_compressed_i,
	instr_ret_spec_i,
	instr_ret_compressed_spec_i,
	iside_wait_i,
	jump_i,
	branch_i,
	branch_taken_i,
	mem_load_i,
	mem_store_i,
	dside_wait_i,
	mul_wait_i,
	div_wait_i
);
	reg _sv2v_0;
	// Trace: design.sv:36719:13
	parameter [0:0] DbgTriggerEn = 0;
	// Trace: design.sv:36720:13
	parameter [31:0] DbgHwBreakNum = 1;
	// Trace: design.sv:36721:13
	parameter [0:0] DataIndTiming = 1'b0;
	// Trace: design.sv:36722:13
	parameter [0:0] DummyInstructions = 1'b0;
	// Trace: design.sv:36723:13
	parameter [0:0] ShadowCSR = 1'b0;
	// Trace: design.sv:36724:13
	parameter [0:0] ICache = 1'b0;
	// Trace: design.sv:36725:13
	parameter [31:0] MHPMCounterNum = 10;
	// Trace: design.sv:36726:13
	parameter [31:0] MHPMCounterWidth = 40;
	// Trace: design.sv:36727:13
	parameter [0:0] PMPEnable = 0;
	// Trace: design.sv:36728:13
	parameter [31:0] PMPGranularity = 0;
	// Trace: design.sv:36729:13
	parameter [31:0] PMPNumRegions = 4;
	// Trace: design.sv:36730:13
	parameter [0:0] RV32E = 0;
	// Trace: design.sv:36731:13
	// removed localparam type ibex_pkg_rv32m_e
	parameter integer RV32M = 32'sd2;
	// Trace: design.sv:36732:13
	// removed localparam type ibex_pkg_rv32b_e
	parameter integer RV32B = 32'sd0;
	// Trace: design.sv:36735:3
	input wire clk_i;
	// Trace: design.sv:36736:3
	input wire rst_ni;
	// Trace: design.sv:36739:3
	input wire [31:0] hart_id_i;
	// Trace: design.sv:36742:3
	// removed localparam type ibex_pkg_priv_lvl_e
	output wire [1:0] priv_mode_id_o;
	// Trace: design.sv:36743:3
	output wire [1:0] priv_mode_lsu_o;
	// Trace: design.sv:36744:3
	output wire csr_mstatus_tw_o;
	// Trace: design.sv:36747:3
	output wire [31:0] csr_mtvec_o;
	// Trace: design.sv:36748:3
	input wire csr_mtvec_init_i;
	// Trace: design.sv:36749:3
	input wire [31:0] boot_addr_i;
	// Trace: design.sv:36752:3
	input wire csr_access_i;
	// Trace: design.sv:36753:3
	// removed localparam type ibex_pkg_csr_num_e
	input wire [11:0] csr_addr_i;
	// Trace: design.sv:36754:3
	input wire [31:0] csr_wdata_i;
	// Trace: design.sv:36755:3
	// removed localparam type ibex_pkg_csr_op_e
	input wire [1:0] csr_op_i;
	// Trace: design.sv:36756:3
	input csr_op_en_i;
	// Trace: design.sv:36757:3
	output wire [31:0] csr_rdata_o;
	// Trace: design.sv:36760:3
	input wire irq_software_i;
	// Trace: design.sv:36761:3
	input wire irq_timer_i;
	// Trace: design.sv:36762:3
	input wire irq_external_i;
	// Trace: design.sv:36763:3
	input wire [14:0] irq_fast_i;
	// Trace: design.sv:36764:3
	input wire nmi_mode_i;
	// Trace: design.sv:36765:3
	output wire irq_pending_o;
	// Trace: design.sv:36766:3
	// removed localparam type ibex_pkg_irqs_t
	output wire [17:0] irqs_o;
	// Trace: design.sv:36767:3
	output wire csr_mstatus_mie_o;
	// Trace: design.sv:36768:3
	output wire [31:0] csr_mepc_o;
	// Trace: design.sv:36771:3
	// removed localparam type ibex_pkg_pmp_cfg_mode_e
	// removed localparam type ibex_pkg_pmp_cfg_t
	output wire [(PMPNumRegions * 6) - 1:0] csr_pmp_cfg_o;
	// Trace: design.sv:36772:3
	output wire [(PMPNumRegions * 34) - 1:0] csr_pmp_addr_o;
	// Trace: design.sv:36773:3
	// removed localparam type ibex_pkg_pmp_mseccfg_t
	output wire [2:0] csr_pmp_mseccfg_o;
	// Trace: design.sv:36776:3
	input wire debug_mode_i;
	// Trace: design.sv:36777:3
	// removed localparam type ibex_pkg_dbg_cause_e
	input wire [2:0] debug_cause_i;
	// Trace: design.sv:36778:3
	input wire debug_csr_save_i;
	// Trace: design.sv:36779:3
	output wire [31:0] csr_depc_o;
	// Trace: design.sv:36780:3
	output wire debug_single_step_o;
	// Trace: design.sv:36781:3
	output wire debug_ebreakm_o;
	// Trace: design.sv:36782:3
	output wire debug_ebreaku_o;
	// Trace: design.sv:36783:3
	output wire trigger_match_o;
	// Trace: design.sv:36785:3
	input wire [31:0] pc_if_i;
	// Trace: design.sv:36786:3
	input wire [31:0] pc_id_i;
	// Trace: design.sv:36787:3
	input wire [31:0] pc_wb_i;
	// Trace: design.sv:36790:3
	output wire data_ind_timing_o;
	// Trace: design.sv:36791:3
	output wire dummy_instr_en_o;
	// Trace: design.sv:36792:3
	output wire [2:0] dummy_instr_mask_o;
	// Trace: design.sv:36793:3
	output wire dummy_instr_seed_en_o;
	// Trace: design.sv:36794:3
	output wire [31:0] dummy_instr_seed_o;
	// Trace: design.sv:36795:3
	output wire icache_enable_o;
	// Trace: design.sv:36796:3
	output wire csr_shadow_err_o;
	// Trace: design.sv:36799:3
	input wire csr_save_if_i;
	// Trace: design.sv:36800:3
	input wire csr_save_id_i;
	// Trace: design.sv:36801:3
	input wire csr_save_wb_i;
	// Trace: design.sv:36802:3
	input wire csr_restore_mret_i;
	// Trace: design.sv:36803:3
	input wire csr_restore_dret_i;
	// Trace: design.sv:36804:3
	input wire csr_save_cause_i;
	// Trace: design.sv:36805:3
	// removed localparam type ibex_pkg_exc_cause_e
	input wire [5:0] csr_mcause_i;
	// Trace: design.sv:36806:3
	input wire [31:0] csr_mtval_i;
	// Trace: design.sv:36807:3
	output wire illegal_csr_insn_o;
	// Trace: design.sv:36810:3
	output reg double_fault_seen_o;
	// Trace: design.sv:36812:3
	input wire instr_ret_i;
	// Trace: design.sv:36813:3
	input wire instr_ret_compressed_i;
	// Trace: design.sv:36814:3
	input wire instr_ret_spec_i;
	// Trace: design.sv:36815:3
	input wire instr_ret_compressed_spec_i;
	// Trace: design.sv:36816:3
	input wire iside_wait_i;
	// Trace: design.sv:36817:3
	input wire jump_i;
	// Trace: design.sv:36818:3
	input wire branch_i;
	// Trace: design.sv:36819:3
	input wire branch_taken_i;
	// Trace: design.sv:36820:3
	input wire mem_load_i;
	// Trace: design.sv:36821:3
	input wire mem_store_i;
	// Trace: design.sv:36822:3
	input wire dside_wait_i;
	// Trace: design.sv:36823:3
	input wire mul_wait_i;
	// Trace: design.sv:36824:3
	input wire div_wait_i;
	// Trace: design.sv:36827:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:36829:3
	localparam [31:0] RV32BEnabled = (RV32B == 32'sd0 ? 0 : 1);
	// Trace: design.sv:36830:3
	localparam [31:0] RV32MEnabled = (RV32M == 32'sd0 ? 0 : 1);
	// Trace: design.sv:36831:3
	localparam [31:0] PMPAddrWidth = (PMPGranularity > 0 ? 33 - PMPGranularity : 32);
	// Trace: design.sv:36834:3
	localparam [1:0] ibex_pkg_CSR_MISA_MXL = 2'd1;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	localparam [31:0] MISA_VALUE = (((((((((((0 | (RV32BEnabled << 1)) | 4) | 0) | (sv2v_cast_32(RV32E) << 4)) | 0) | (sv2v_cast_32(!RV32E) << 8)) | (RV32MEnabled << 12)) | 0) | 0) | 1048576) | 0) | (sv2v_cast_32(ibex_pkg_CSR_MISA_MXL) << 30);
	// Trace: design.sv:36849:3
	// removed localparam type status_t
	// Trace: design.sv:36857:3
	// removed localparam type status_stk_t
	// Trace: design.sv:36862:3
	// removed localparam type ibex_pkg_x_debug_ver_e
	// removed localparam type dcsr_t
	// Trace: design.sv:36881:3
	// removed localparam type cpu_ctrl_t
	// Trace: design.sv:36891:3
	reg [31:0] exception_pc;
	// Trace: design.sv:36894:3
	reg [1:0] priv_lvl_q;
	reg [1:0] priv_lvl_d;
	// Trace: design.sv:36895:3
	wire [5:0] mstatus_q;
	reg [5:0] mstatus_d;
	// Trace: design.sv:36896:3
	wire mstatus_err;
	// Trace: design.sv:36897:3
	reg mstatus_en;
	// Trace: design.sv:36898:3
	wire [17:0] mie_q;
	wire [17:0] mie_d;
	// Trace: design.sv:36899:3
	reg mie_en;
	// Trace: design.sv:36900:3
	wire [31:0] mscratch_q;
	// Trace: design.sv:36901:3
	reg mscratch_en;
	// Trace: design.sv:36902:3
	wire [31:0] mepc_q;
	reg [31:0] mepc_d;
	// Trace: design.sv:36903:3
	reg mepc_en;
	// Trace: design.sv:36904:3
	wire [5:0] mcause_q;
	reg [5:0] mcause_d;
	// Trace: design.sv:36905:3
	reg mcause_en;
	// Trace: design.sv:36906:3
	wire [31:0] mtval_q;
	reg [31:0] mtval_d;
	// Trace: design.sv:36907:3
	reg mtval_en;
	// Trace: design.sv:36908:3
	wire [31:0] mtvec_q;
	reg [31:0] mtvec_d;
	// Trace: design.sv:36909:3
	wire mtvec_err;
	// Trace: design.sv:36910:3
	reg mtvec_en;
	// Trace: design.sv:36911:3
	wire [17:0] mip;
	// Trace: design.sv:36912:3
	wire [31:0] dcsr_q;
	reg [31:0] dcsr_d;
	// Trace: design.sv:36913:3
	reg dcsr_en;
	// Trace: design.sv:36914:3
	wire [31:0] depc_q;
	reg [31:0] depc_d;
	// Trace: design.sv:36915:3
	reg depc_en;
	// Trace: design.sv:36916:3
	wire [31:0] dscratch0_q;
	// Trace: design.sv:36917:3
	wire [31:0] dscratch1_q;
	// Trace: design.sv:36918:3
	reg dscratch0_en;
	reg dscratch1_en;
	// Trace: design.sv:36922:3
	wire [2:0] mstack_q;
	reg [2:0] mstack_d;
	// Trace: design.sv:36923:3
	reg mstack_en;
	// Trace: design.sv:36924:3
	wire [31:0] mstack_epc_q;
	reg [31:0] mstack_epc_d;
	// Trace: design.sv:36925:3
	wire [5:0] mstack_cause_q;
	reg [5:0] mstack_cause_d;
	// Trace: design.sv:36928:3
	localparam [31:0] ibex_pkg_PMP_MAX_REGIONS = 16;
	reg [31:0] pmp_addr_rdata [0:15];
	// Trace: design.sv:36929:3
	localparam [31:0] ibex_pkg_PMP_CFG_W = 8;
	wire [7:0] pmp_cfg_rdata [0:15];
	// Trace: design.sv:36930:3
	wire pmp_csr_err;
	// Trace: design.sv:36931:3
	wire [2:0] pmp_mseccfg;
	// Trace: design.sv:36934:3
	wire [31:0] mcountinhibit;
	// Trace: design.sv:36936:3
	reg [MHPMCounterNum + 2:0] mcountinhibit_d;
	reg [MHPMCounterNum + 2:0] mcountinhibit_q;
	// Trace: design.sv:36937:3
	reg mcountinhibit_we;
	// Trace: design.sv:36942:3
	wire [63:0] mhpmcounter [0:31];
	// Trace: design.sv:36943:3
	reg [31:0] mhpmcounter_we;
	// Trace: design.sv:36944:3
	reg [31:0] mhpmcounterh_we;
	// Trace: design.sv:36945:3
	reg [31:0] mhpmcounter_incr;
	// Trace: design.sv:36946:3
	reg [31:0] mhpmevent [0:31];
	// Trace: design.sv:36947:3
	wire [4:0] mhpmcounter_idx;
	// Trace: design.sv:36948:3
	wire unused_mhpmcounter_we_1;
	// Trace: design.sv:36949:3
	wire unused_mhpmcounterh_we_1;
	// Trace: design.sv:36950:3
	wire unused_mhpmcounter_incr_1;
	// Trace: design.sv:36952:3
	wire [63:0] minstret_next;
	wire [63:0] minstret_raw;
	// Trace: design.sv:36955:3
	wire [31:0] tselect_rdata;
	// Trace: design.sv:36956:3
	wire [31:0] tmatch_control_rdata;
	// Trace: design.sv:36957:3
	wire [31:0] tmatch_value_rdata;
	// Trace: design.sv:36960:3
	wire [7:0] cpuctrl_q;
	reg [7:0] cpuctrl_d;
	wire [7:0] cpuctrl_wdata_raw;
	wire [7:0] cpuctrl_wdata;
	// Trace: design.sv:36961:3
	reg cpuctrl_we;
	// Trace: design.sv:36962:3
	wire cpuctrl_err;
	// Trace: design.sv:36965:3
	reg [31:0] csr_wdata_int;
	// Trace: design.sv:36966:3
	reg [31:0] csr_rdata_int;
	// Trace: design.sv:36967:3
	wire csr_we_int;
	// Trace: design.sv:36968:3
	wire csr_wr;
	// Trace: design.sv:36971:3
	reg illegal_csr;
	// Trace: design.sv:36972:3
	wire illegal_csr_priv;
	// Trace: design.sv:36973:3
	wire illegal_csr_write;
	// Trace: design.sv:36975:3
	wire [7:0] unused_boot_addr;
	// Trace: design.sv:36976:3
	wire [2:0] unused_csr_addr;
	// Trace: design.sv:36978:3
	assign unused_boot_addr = boot_addr_i[7:0];
	// Trace: design.sv:36984:3
	wire [11:0] csr_addr;
	// Trace: design.sv:36985:3
	assign csr_addr = {csr_addr_i};
	// Trace: design.sv:36986:3
	assign unused_csr_addr = csr_addr[7:5];
	// Trace: design.sv:36987:3
	assign mhpmcounter_idx = csr_addr[4:0];
	// Trace: design.sv:36990:3
	assign illegal_csr_priv = csr_addr[9:8] > {priv_lvl_q};
	// Trace: design.sv:36991:3
	assign illegal_csr_write = (csr_addr[11:10] == 2'b11) && csr_wr;
	// Trace: design.sv:36992:3
	assign illegal_csr_insn_o = csr_access_i & ((illegal_csr | illegal_csr_write) | illegal_csr_priv);
	// Trace: design.sv:36995:3
	assign mip[17] = irq_software_i;
	// Trace: design.sv:36996:3
	assign mip[16] = irq_timer_i;
	// Trace: design.sv:36997:3
	assign mip[15] = irq_external_i;
	// Trace: design.sv:36998:3
	assign mip[14-:15] = irq_fast_i;
	// Trace: design.sv:37001:3
	localparam [31:0] ibex_pkg_CSR_MARCHID_VALUE = 32'h00000016;
	localparam [31:0] ibex_pkg_CSR_MEIX_BIT = 11;
	localparam [31:0] ibex_pkg_CSR_MFIX_BIT_HIGH = 30;
	localparam [31:0] ibex_pkg_CSR_MFIX_BIT_LOW = 16;
	localparam [31:0] ibex_pkg_CSR_MIMPID_VALUE = 32'b00000000000000000000000000000000;
	localparam [31:0] ibex_pkg_CSR_MSECCFG_MML_BIT = 0;
	localparam [31:0] ibex_pkg_CSR_MSECCFG_MMWP_BIT = 1;
	localparam [31:0] ibex_pkg_CSR_MSECCFG_RLB_BIT = 2;
	localparam [31:0] ibex_pkg_CSR_MSIX_BIT = 3;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MIE_BIT = 3;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MPIE_BIT = 7;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MPP_BIT_HIGH = 12;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MPP_BIT_LOW = 11;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MPRV_BIT = 17;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_TW_BIT = 21;
	localparam [31:0] ibex_pkg_CSR_MTIX_BIT = 7;
	localparam [31:0] ibex_pkg_CSR_MVENDORID_VALUE = 32'b00000000000000000000000000000000;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:37002:5
		csr_rdata_int = 1'sb0;
		// Trace: design.sv:37003:5
		illegal_csr = 1'b0;
		// Trace: design.sv:37005:5
		(* full_case, parallel_case *)
		case (csr_addr_i)
			12'hf11:
				// Trace: design.sv:37007:22
				csr_rdata_int = ibex_pkg_CSR_MVENDORID_VALUE;
			12'hf12:
				// Trace: design.sv:37009:20
				csr_rdata_int = ibex_pkg_CSR_MARCHID_VALUE;
			12'hf13:
				// Trace: design.sv:37011:19
				csr_rdata_int = ibex_pkg_CSR_MIMPID_VALUE;
			12'hf14:
				// Trace: design.sv:37013:20
				csr_rdata_int = hart_id_i;
			12'h300: begin
				// Trace: design.sv:37017:9
				csr_rdata_int = 1'sb0;
				// Trace: design.sv:37018:9
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_MIE_BIT] = mstatus_q[5];
				// Trace: design.sv:37019:9
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_MPIE_BIT] = mstatus_q[4];
				// Trace: design.sv:37020:9
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_MPP_BIT_HIGH:ibex_pkg_CSR_MSTATUS_MPP_BIT_LOW] = mstatus_q[3-:2];
				// Trace: design.sv:37021:9
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_MPRV_BIT] = mstatus_q[1];
				// Trace: design.sv:37022:9
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_TW_BIT] = mstatus_q[0];
			end
			12'h301:
				// Trace: design.sv:37026:17
				csr_rdata_int = MISA_VALUE;
			12'h304: begin
				// Trace: design.sv:37030:9
				csr_rdata_int = 1'sb0;
				// Trace: design.sv:37031:9
				csr_rdata_int[ibex_pkg_CSR_MSIX_BIT] = mie_q[17];
				// Trace: design.sv:37032:9
				csr_rdata_int[ibex_pkg_CSR_MTIX_BIT] = mie_q[16];
				// Trace: design.sv:37033:9
				csr_rdata_int[ibex_pkg_CSR_MEIX_BIT] = mie_q[15];
				// Trace: design.sv:37034:9
				csr_rdata_int[ibex_pkg_CSR_MFIX_BIT_HIGH:ibex_pkg_CSR_MFIX_BIT_LOW] = mie_q[14-:15];
			end
			12'h306:
				// Trace: design.sv:37039:9
				csr_rdata_int = 1'sb0;
			12'h340:
				// Trace: design.sv:37042:21
				csr_rdata_int = mscratch_q;
			12'h305:
				// Trace: design.sv:37045:18
				csr_rdata_int = mtvec_q;
			12'h341:
				// Trace: design.sv:37048:17
				csr_rdata_int = mepc_q;
			12'h342:
				// Trace: design.sv:37051:19
				csr_rdata_int = {mcause_q[5], 26'b00000000000000000000000000, mcause_q[4:0]};
			12'h343:
				// Trace: design.sv:37054:18
				csr_rdata_int = mtval_q;
			12'h344: begin
				// Trace: design.sv:37058:9
				csr_rdata_int = 1'sb0;
				// Trace: design.sv:37059:9
				csr_rdata_int[ibex_pkg_CSR_MSIX_BIT] = mip[17];
				// Trace: design.sv:37060:9
				csr_rdata_int[ibex_pkg_CSR_MTIX_BIT] = mip[16];
				// Trace: design.sv:37061:9
				csr_rdata_int[ibex_pkg_CSR_MEIX_BIT] = mip[15];
				// Trace: design.sv:37062:9
				csr_rdata_int[ibex_pkg_CSR_MFIX_BIT_HIGH:ibex_pkg_CSR_MFIX_BIT_LOW] = mip[14-:15];
			end
			12'h747:
				// Trace: design.sv:37066:9
				if (PMPEnable) begin
					// Trace: design.sv:37067:11
					csr_rdata_int = 1'sb0;
					// Trace: design.sv:37068:11
					csr_rdata_int[ibex_pkg_CSR_MSECCFG_MML_BIT] = pmp_mseccfg[0];
					// Trace: design.sv:37069:11
					csr_rdata_int[ibex_pkg_CSR_MSECCFG_MMWP_BIT] = pmp_mseccfg[1];
					// Trace: design.sv:37070:11
					csr_rdata_int[ibex_pkg_CSR_MSECCFG_RLB_BIT] = pmp_mseccfg[2];
				end
				else
					// Trace: design.sv:37072:11
					illegal_csr = 1'b1;
			12'h757:
				// Trace: design.sv:37077:9
				if (PMPEnable)
					// Trace: design.sv:37078:11
					csr_rdata_int = 1'sb0;
				else
					// Trace: design.sv:37080:11
					illegal_csr = 1'b1;
			12'h3a0:
				// Trace: design.sv:37085:22
				csr_rdata_int = {pmp_cfg_rdata[3], pmp_cfg_rdata[2], pmp_cfg_rdata[1], pmp_cfg_rdata[0]};
			12'h3a1:
				// Trace: design.sv:37087:22
				csr_rdata_int = {pmp_cfg_rdata[7], pmp_cfg_rdata[6], pmp_cfg_rdata[5], pmp_cfg_rdata[4]};
			12'h3a2:
				// Trace: design.sv:37089:22
				csr_rdata_int = {pmp_cfg_rdata[11], pmp_cfg_rdata[10], pmp_cfg_rdata[9], pmp_cfg_rdata[8]};
			12'h3a3:
				// Trace: design.sv:37091:22
				csr_rdata_int = {pmp_cfg_rdata[15], pmp_cfg_rdata[14], pmp_cfg_rdata[13], pmp_cfg_rdata[12]};
			12'h3b0:
				// Trace: design.sv:37093:22
				csr_rdata_int = pmp_addr_rdata[0];
			12'h3b1:
				// Trace: design.sv:37094:22
				csr_rdata_int = pmp_addr_rdata[1];
			12'h3b2:
				// Trace: design.sv:37095:22
				csr_rdata_int = pmp_addr_rdata[2];
			12'h3b3:
				// Trace: design.sv:37096:22
				csr_rdata_int = pmp_addr_rdata[3];
			12'h3b4:
				// Trace: design.sv:37097:22
				csr_rdata_int = pmp_addr_rdata[4];
			12'h3b5:
				// Trace: design.sv:37098:22
				csr_rdata_int = pmp_addr_rdata[5];
			12'h3b6:
				// Trace: design.sv:37099:22
				csr_rdata_int = pmp_addr_rdata[6];
			12'h3b7:
				// Trace: design.sv:37100:22
				csr_rdata_int = pmp_addr_rdata[7];
			12'h3b8:
				// Trace: design.sv:37101:22
				csr_rdata_int = pmp_addr_rdata[8];
			12'h3b9:
				// Trace: design.sv:37102:22
				csr_rdata_int = pmp_addr_rdata[9];
			12'h3ba:
				// Trace: design.sv:37103:22
				csr_rdata_int = pmp_addr_rdata[10];
			12'h3bb:
				// Trace: design.sv:37104:22
				csr_rdata_int = pmp_addr_rdata[11];
			12'h3bc:
				// Trace: design.sv:37105:22
				csr_rdata_int = pmp_addr_rdata[12];
			12'h3bd:
				// Trace: design.sv:37106:22
				csr_rdata_int = pmp_addr_rdata[13];
			12'h3be:
				// Trace: design.sv:37107:22
				csr_rdata_int = pmp_addr_rdata[14];
			12'h3bf:
				// Trace: design.sv:37108:22
				csr_rdata_int = pmp_addr_rdata[15];
			12'h7b0: begin
				// Trace: design.sv:37111:9
				csr_rdata_int = dcsr_q;
				// Trace: design.sv:37112:9
				illegal_csr = ~debug_mode_i;
			end
			12'h7b1: begin
				// Trace: design.sv:37115:9
				csr_rdata_int = depc_q;
				// Trace: design.sv:37116:9
				illegal_csr = ~debug_mode_i;
			end
			12'h7b2: begin
				// Trace: design.sv:37119:9
				csr_rdata_int = dscratch0_q;
				// Trace: design.sv:37120:9
				illegal_csr = ~debug_mode_i;
			end
			12'h7b3: begin
				// Trace: design.sv:37123:9
				csr_rdata_int = dscratch1_q;
				// Trace: design.sv:37124:9
				illegal_csr = ~debug_mode_i;
			end
			12'h320:
				// Trace: design.sv:37128:26
				csr_rdata_int = mcountinhibit;
			12'h323, 12'h324, 12'h325, 12'h326, 12'h327, 12'h328, 12'h329, 12'h32a, 12'h32b, 12'h32c, 12'h32d, 12'h32e, 12'h32f, 12'h330, 12'h331, 12'h332, 12'h333, 12'h334, 12'h335, 12'h336, 12'h337, 12'h338, 12'h339, 12'h33a, 12'h33b, 12'h33c, 12'h33d, 12'h33e, 12'h33f:
				// Trace: design.sv:37137:9
				csr_rdata_int = mhpmevent[mhpmcounter_idx];
			12'hb00, 12'hb02, 12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f:
				// Trace: design.sv:37150:9
				csr_rdata_int = mhpmcounter[mhpmcounter_idx][31:0];
			12'hb80, 12'hb82, 12'hb83, 12'hb84, 12'hb85, 12'hb86, 12'hb87, 12'hb88, 12'hb89, 12'hb8a, 12'hb8b, 12'hb8c, 12'hb8d, 12'hb8e, 12'hb8f, 12'hb90, 12'hb91, 12'hb92, 12'hb93, 12'hb94, 12'hb95, 12'hb96, 12'hb97, 12'hb98, 12'hb99, 12'hb9a, 12'hb9b, 12'hb9c, 12'hb9d, 12'hb9e, 12'hb9f:
				// Trace: design.sv:37163:9
				csr_rdata_int = mhpmcounter[mhpmcounter_idx][63:32];
			12'h7a0: begin
				// Trace: design.sv:37168:9
				csr_rdata_int = tselect_rdata;
				// Trace: design.sv:37169:9
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7a1: begin
				// Trace: design.sv:37172:9
				csr_rdata_int = tmatch_control_rdata;
				// Trace: design.sv:37173:9
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7a2: begin
				// Trace: design.sv:37176:9
				csr_rdata_int = tmatch_value_rdata;
				// Trace: design.sv:37177:9
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7a3: begin
				// Trace: design.sv:37180:9
				csr_rdata_int = 1'sb0;
				// Trace: design.sv:37181:9
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7a8: begin
				// Trace: design.sv:37184:9
				csr_rdata_int = 1'sb0;
				// Trace: design.sv:37185:9
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7aa: begin
				// Trace: design.sv:37188:9
				csr_rdata_int = 1'sb0;
				// Trace: design.sv:37189:9
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7c0:
				// Trace: design.sv:37194:9
				csr_rdata_int = {{24 {1'b0}}, cpuctrl_q};
			12'h7c1:
				// Trace: design.sv:37199:9
				csr_rdata_int = 1'sb0;
			default:
				// Trace: design.sv:37203:9
				illegal_csr = 1'b1;
		endcase
	end
	// Trace: design.sv:37209:3
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:37210:5
		exception_pc = pc_id_i;
		// Trace: design.sv:37212:5
		priv_lvl_d = priv_lvl_q;
		// Trace: design.sv:37213:5
		mstatus_en = 1'b0;
		// Trace: design.sv:37214:5
		mstatus_d = mstatus_q;
		// Trace: design.sv:37215:5
		mie_en = 1'b0;
		// Trace: design.sv:37216:5
		mscratch_en = 1'b0;
		// Trace: design.sv:37217:5
		mepc_en = 1'b0;
		// Trace: design.sv:37218:5
		mepc_d = {csr_wdata_int[31:1], 1'b0};
		// Trace: design.sv:37219:5
		mcause_en = 1'b0;
		// Trace: design.sv:37220:5
		mcause_d = {csr_wdata_int[31], csr_wdata_int[4:0]};
		// Trace: design.sv:37221:5
		mtval_en = 1'b0;
		// Trace: design.sv:37222:5
		mtval_d = csr_wdata_int;
		// Trace: design.sv:37223:5
		mtvec_en = csr_mtvec_init_i;
		// Trace: design.sv:37226:5
		mtvec_d = (csr_mtvec_init_i ? {boot_addr_i[31:8], 8'b00000001} : {csr_wdata_int[31:8], 8'b00000001});
		// Trace: design.sv:37228:5
		dcsr_en = 1'b0;
		// Trace: design.sv:37229:5
		dcsr_d = dcsr_q;
		// Trace: design.sv:37230:5
		depc_d = {csr_wdata_int[31:1], 1'b0};
		// Trace: design.sv:37231:5
		depc_en = 1'b0;
		// Trace: design.sv:37232:5
		dscratch0_en = 1'b0;
		// Trace: design.sv:37233:5
		dscratch1_en = 1'b0;
		// Trace: design.sv:37235:5
		mstack_en = 1'b0;
		// Trace: design.sv:37236:5
		mstack_d[2] = mstatus_q[4];
		// Trace: design.sv:37237:5
		mstack_d[1-:2] = mstatus_q[3-:2];
		// Trace: design.sv:37238:5
		mstack_epc_d = mepc_q;
		// Trace: design.sv:37239:5
		mstack_cause_d = mcause_q;
		// Trace: design.sv:37241:5
		mcountinhibit_we = 1'b0;
		// Trace: design.sv:37242:5
		mhpmcounter_we = 1'sb0;
		// Trace: design.sv:37243:5
		mhpmcounterh_we = 1'sb0;
		// Trace: design.sv:37245:5
		cpuctrl_we = 1'b0;
		// Trace: design.sv:37246:5
		cpuctrl_d = cpuctrl_q;
		// Trace: design.sv:37248:5
		double_fault_seen_o = 1'b0;
		// Trace: design.sv:37250:5
		if (csr_we_int)
			// Trace: design.sv:37251:7
			(* full_case, parallel_case *)
			case (csr_addr_i)
				12'h300: begin
					// Trace: design.sv:37254:11
					mstatus_en = 1'b1;
					// Trace: design.sv:37255:11
					mstatus_d = {csr_wdata_int[ibex_pkg_CSR_MSTATUS_MIE_BIT], csr_wdata_int[ibex_pkg_CSR_MSTATUS_MPIE_BIT], sv2v_cast_2(csr_wdata_int[ibex_pkg_CSR_MSTATUS_MPP_BIT_HIGH:ibex_pkg_CSR_MSTATUS_MPP_BIT_LOW]), csr_wdata_int[ibex_pkg_CSR_MSTATUS_MPRV_BIT], csr_wdata_int[ibex_pkg_CSR_MSTATUS_TW_BIT]};
					// Trace: design.sv:37263:11
					if ((mstatus_d[3-:2] != 2'b11) && (mstatus_d[3-:2] != 2'b00))
						// Trace: design.sv:37264:13
						mstatus_d[3-:2] = 2'b11;
				end
				12'h304:
					// Trace: design.sv:37269:18
					mie_en = 1'b1;
				12'h340:
					// Trace: design.sv:37271:23
					mscratch_en = 1'b1;
				12'h341:
					// Trace: design.sv:37274:19
					mepc_en = 1'b1;
				12'h342:
					// Trace: design.sv:37277:21
					mcause_en = 1'b1;
				12'h343:
					// Trace: design.sv:37280:20
					mtval_en = 1'b1;
				12'h305:
					// Trace: design.sv:37283:20
					mtvec_en = 1'b1;
				12'h7b0: begin
					// Trace: design.sv:37286:11
					dcsr_d = csr_wdata_int;
					// Trace: design.sv:37287:11
					dcsr_d[31-:4] = 4'd4;
					// Trace: design.sv:37289:11
					if ((dcsr_d[1-:2] != 2'b11) && (dcsr_d[1-:2] != 2'b00))
						// Trace: design.sv:37290:13
						dcsr_d[1-:2] = 2'b11;
					// Trace: design.sv:37294:11
					dcsr_d[8-:3] = dcsr_q[8-:3];
					// Trace: design.sv:37297:11
					dcsr_d[11] = 1'b0;
					// Trace: design.sv:37300:11
					dcsr_d[3] = 1'b0;
					// Trace: design.sv:37301:11
					dcsr_d[4] = 1'b0;
					// Trace: design.sv:37302:11
					dcsr_d[10] = 1'b0;
					// Trace: design.sv:37303:11
					dcsr_d[9] = 1'b0;
					// Trace: design.sv:37306:11
					dcsr_d[5] = 1'b0;
					// Trace: design.sv:37307:11
					dcsr_d[14] = 1'b0;
					// Trace: design.sv:37308:11
					dcsr_d[27-:12] = 12'h000;
					// Trace: design.sv:37309:11
					dcsr_en = 1'b1;
				end
				12'h7b1:
					// Trace: design.sv:37313:18
					depc_en = 1'b1;
				12'h7b2:
					// Trace: design.sv:37315:24
					dscratch0_en = 1'b1;
				12'h7b3:
					// Trace: design.sv:37316:24
					dscratch1_en = 1'b1;
				12'h320:
					// Trace: design.sv:37319:28
					mcountinhibit_we = 1'b1;
				12'hb00, 12'hb02, 12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f:
					// Trace: design.sv:37331:11
					mhpmcounter_we[mhpmcounter_idx] = 1'b1;
				12'hb80, 12'hb82, 12'hb83, 12'hb84, 12'hb85, 12'hb86, 12'hb87, 12'hb88, 12'hb89, 12'hb8a, 12'hb8b, 12'hb8c, 12'hb8d, 12'hb8e, 12'hb8f, 12'hb90, 12'hb91, 12'hb92, 12'hb93, 12'hb94, 12'hb95, 12'hb96, 12'hb97, 12'hb98, 12'hb99, 12'hb9a, 12'hb9b, 12'hb9c, 12'hb9d, 12'hb9e, 12'hb9f:
					// Trace: design.sv:37344:11
					mhpmcounterh_we[mhpmcounter_idx] = 1'b1;
				12'h7c0: begin
					// Trace: design.sv:37348:11
					cpuctrl_d = cpuctrl_wdata;
					// Trace: design.sv:37349:11
					cpuctrl_we = 1'b1;
				end
				default:
					;
			endcase
		(* full_case, parallel_case *)
		case (1'b1)
			csr_save_cause_i: begin
				// Trace: design.sv:37360:9
				(* full_case, parallel_case *)
				case (1'b1)
					csr_save_if_i:
						// Trace: design.sv:37362:13
						exception_pc = pc_if_i;
					csr_save_id_i:
						// Trace: design.sv:37365:13
						exception_pc = pc_id_i;
					csr_save_wb_i:
						// Trace: design.sv:37368:13
						exception_pc = pc_wb_i;
					default:
						;
				endcase
				// Trace: design.sv:37374:9
				priv_lvl_d = 2'b11;
				if (debug_csr_save_i) begin
					// Trace: design.sv:37379:11
					dcsr_d[1-:2] = priv_lvl_q;
					// Trace: design.sv:37380:11
					dcsr_d[8-:3] = debug_cause_i;
					// Trace: design.sv:37381:11
					dcsr_en = 1'b1;
					// Trace: design.sv:37382:11
					depc_d = exception_pc;
					// Trace: design.sv:37383:11
					depc_en = 1'b1;
				end
				else if (!debug_mode_i) begin
					// Trace: design.sv:37387:11
					mtval_en = 1'b1;
					// Trace: design.sv:37388:11
					mtval_d = csr_mtval_i;
					// Trace: design.sv:37389:11
					mstatus_en = 1'b1;
					// Trace: design.sv:37390:11
					mstatus_d[5] = 1'b0;
					// Trace: design.sv:37392:11
					mstatus_d[4] = mstatus_q[5];
					// Trace: design.sv:37393:11
					mstatus_d[3-:2] = priv_lvl_q;
					// Trace: design.sv:37394:11
					mepc_en = 1'b1;
					// Trace: design.sv:37395:11
					mepc_d = exception_pc;
					// Trace: design.sv:37396:11
					mcause_en = 1'b1;
					// Trace: design.sv:37397:11
					mcause_d = {csr_mcause_i};
					// Trace: design.sv:37399:11
					mstack_en = 1'b1;
					// Trace: design.sv:37401:11
					if (!mcause_d[5]) begin
						// Trace: design.sv:37404:13
						cpuctrl_we = 1'b1;
						// Trace: design.sv:37406:13
						cpuctrl_d[6] = 1'b1;
						// Trace: design.sv:37407:13
						if (cpuctrl_q[6]) begin
							// Trace: design.sv:37408:15
							double_fault_seen_o = 1'b1;
							// Trace: design.sv:37409:15
							cpuctrl_d[7] = 1'b1;
						end
					end
				end
			end
			csr_restore_dret_i:
				// Trace: design.sv:37416:9
				priv_lvl_d = dcsr_q[1-:2];
			csr_restore_mret_i: begin
				// Trace: design.sv:37420:9
				priv_lvl_d = mstatus_q[3-:2];
				// Trace: design.sv:37421:9
				mstatus_en = 1'b1;
				// Trace: design.sv:37422:9
				mstatus_d[5] = mstatus_q[4];
				// Trace: design.sv:37426:9
				cpuctrl_we = 1'b1;
				// Trace: design.sv:37427:9
				cpuctrl_d[6] = 1'b0;
				// Trace: design.sv:37429:9
				if (nmi_mode_i) begin
					// Trace: design.sv:37431:11
					mstatus_d[4] = mstack_q[2];
					// Trace: design.sv:37432:11
					mstatus_d[3-:2] = mstack_q[1-:2];
					// Trace: design.sv:37433:11
					mepc_en = 1'b1;
					// Trace: design.sv:37434:11
					mepc_d = mstack_epc_q;
					// Trace: design.sv:37435:11
					mcause_en = 1'b1;
					// Trace: design.sv:37436:11
					mcause_d = mstack_cause_q;
				end
				else begin
					// Trace: design.sv:37440:11
					mstatus_d[4] = 1'b1;
					// Trace: design.sv:37441:11
					mstatus_d[3-:2] = 2'b00;
				end
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:37450:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:37451:5
		if (!rst_ni)
			// Trace: design.sv:37452:7
			priv_lvl_q <= 2'b11;
		else
			// Trace: design.sv:37454:7
			priv_lvl_q <= priv_lvl_d;
	// Trace: design.sv:37459:3
	assign priv_mode_id_o = priv_lvl_q;
	// Trace: design.sv:37461:3
	assign priv_mode_lsu_o = (mstatus_q[1] ? mstatus_q[3-:2] : priv_lvl_q);
	// Trace: design.sv:37464:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:37465:5
		(* full_case, parallel_case *)
		case (csr_op_i)
			2'd1:
				// Trace: design.sv:37466:21
				csr_wdata_int = csr_wdata_i;
			2'd2:
				// Trace: design.sv:37467:21
				csr_wdata_int = csr_wdata_i | csr_rdata_o;
			2'd3:
				// Trace: design.sv:37468:21
				csr_wdata_int = ~csr_wdata_i & csr_rdata_o;
			2'd0:
				// Trace: design.sv:37469:21
				csr_wdata_int = csr_wdata_i;
			default:
				// Trace: design.sv:37470:21
				csr_wdata_int = csr_wdata_i;
		endcase
	end
	// Trace: design.sv:37474:3
	assign csr_wr = |{csr_op_i == 2'd1, csr_op_i == 2'd2, csr_op_i == 2'd3};
	// Trace: design.sv:37477:3
	assign csr_we_int = (csr_wr & csr_op_en_i) & ~illegal_csr_insn_o;
	// Trace: design.sv:37479:3
	assign csr_rdata_o = csr_rdata_int;
	// Trace: design.sv:37482:3
	assign csr_mepc_o = mepc_q;
	// Trace: design.sv:37483:3
	assign csr_depc_o = depc_q;
	// Trace: design.sv:37484:3
	assign csr_mtvec_o = mtvec_q;
	// Trace: design.sv:37486:3
	assign csr_mstatus_mie_o = mstatus_q[5];
	// Trace: design.sv:37487:3
	assign csr_mstatus_tw_o = mstatus_q[0];
	// Trace: design.sv:37488:3
	assign debug_single_step_o = dcsr_q[2];
	// Trace: design.sv:37489:3
	assign debug_ebreakm_o = dcsr_q[15];
	// Trace: design.sv:37490:3
	assign debug_ebreaku_o = dcsr_q[12];
	// Trace: design.sv:37494:3
	assign irqs_o = mip & mie_q;
	// Trace: design.sv:37495:3
	assign irq_pending_o = |irqs_o;
	// Trace: design.sv:37502:3
	localparam [5:0] MSTATUS_RST_VAL = 6'b010000;
	// Trace: design.sv:37507:3
	ibex_csr #(
		.Width(6),
		.ShadowCopy(ShadowCSR),
		.ResetValue({MSTATUS_RST_VAL})
	) u_mstatus_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({mstatus_d}),
		.wr_en_i(mstatus_en),
		.rd_data_o(mstatus_q),
		.rd_error_o(mstatus_err)
	);
	// Trace: design.sv:37521:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mepc_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mepc_d),
		.wr_en_i(mepc_en),
		.rd_data_o(mepc_q),
		.rd_error_o()
	);
	// Trace: design.sv:37535:3
	assign mie_d[17] = csr_wdata_int[ibex_pkg_CSR_MSIX_BIT];
	// Trace: design.sv:37536:3
	assign mie_d[16] = csr_wdata_int[ibex_pkg_CSR_MTIX_BIT];
	// Trace: design.sv:37537:3
	assign mie_d[15] = csr_wdata_int[ibex_pkg_CSR_MEIX_BIT];
	// Trace: design.sv:37538:3
	assign mie_d[14-:15] = csr_wdata_int[ibex_pkg_CSR_MFIX_BIT_HIGH:ibex_pkg_CSR_MFIX_BIT_LOW];
	// Trace: design.sv:37539:3
	ibex_csr #(
		.Width(18),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mie_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({mie_d}),
		.wr_en_i(mie_en),
		.rd_data_o(mie_q),
		.rd_error_o()
	);
	// Trace: design.sv:37553:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mscratch_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(csr_wdata_int),
		.wr_en_i(mscratch_en),
		.rd_data_o(mscratch_q),
		.rd_error_o()
	);
	// Trace: design.sv:37567:3
	ibex_csr #(
		.Width(6),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mcause_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mcause_d),
		.wr_en_i(mcause_en),
		.rd_data_o(mcause_q),
		.rd_error_o()
	);
	// Trace: design.sv:37581:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mtval_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mtval_d),
		.wr_en_i(mtval_en),
		.rd_data_o(mtval_q),
		.rd_error_o()
	);
	// Trace: design.sv:37595:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(ShadowCSR),
		.ResetValue(32'd1)
	) u_mtvec_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mtvec_d),
		.wr_en_i(mtvec_en),
		.rd_data_o(mtvec_q),
		.rd_error_o(mtvec_err)
	);
	// Trace: design.sv:37609:3
	localparam [31:0] DCSR_RESET_VAL = 32'h40000003;
	// Trace: design.sv:37615:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue({DCSR_RESET_VAL})
	) u_dcsr_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({dcsr_d}),
		.wr_en_i(dcsr_en),
		.rd_data_o(dcsr_q),
		.rd_error_o()
	);
	// Trace: design.sv:37629:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_depc_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(depc_d),
		.wr_en_i(depc_en),
		.rd_data_o(depc_q),
		.rd_error_o()
	);
	// Trace: design.sv:37643:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_dscratch0_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(csr_wdata_int),
		.wr_en_i(dscratch0_en),
		.rd_data_o(dscratch0_q),
		.rd_error_o()
	);
	// Trace: design.sv:37657:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_dscratch1_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(csr_wdata_int),
		.wr_en_i(dscratch1_en),
		.rd_data_o(dscratch1_q),
		.rd_error_o()
	);
	// Trace: design.sv:37671:3
	localparam [2:0] MSTACK_RESET_VAL = 3'b100;
	// Trace: design.sv:37672:3
	ibex_csr #(
		.Width(3),
		.ShadowCopy(1'b0),
		.ResetValue({MSTACK_RESET_VAL})
	) u_mstack_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({mstack_d}),
		.wr_en_i(mstack_en),
		.rd_data_o(mstack_q),
		.rd_error_o()
	);
	// Trace: design.sv:37686:3
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mstack_epc_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mstack_epc_d),
		.wr_en_i(mstack_en),
		.rd_data_o(mstack_epc_q),
		.rd_error_o()
	);
	// Trace: design.sv:37700:3
	ibex_csr #(
		.Width(6),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mstack_cause_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mstack_cause_d),
		.wr_en_i(mstack_en),
		.rd_data_o(mstack_cause_q),
		.rd_error_o()
	);
	// Trace: design.sv:37717:3
	localparam [11:0] ibex_pkg_CSR_OFF_PMP_ADDR = 12'h3b0;
	localparam [11:0] ibex_pkg_CSR_OFF_PMP_CFG = 12'h3a0;
	generate
		if (PMPEnable) begin : g_pmp_registers
			// Trace: ../src/openhwgroup.org_ip_cve2_0/rtl/ibex_pmp_reset_default.svh:12:1
			localparam [95:0] pmp_cfg_rst = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			// Trace: ../src/openhwgroup.org_ip_cve2_0/rtl/ibex_pmp_reset_default.svh:34:1
			localparam [543:0] pmp_addr_rst = 544'h0;
			// Trace: ../src/openhwgroup.org_ip_cve2_0/rtl/ibex_pmp_reset_default.svh:53:1
			localparam [2:0] pmp_mseccfg_rst = 3'b000;
			// Trace: design.sv:37725:5
			wire [2:0] pmp_mseccfg_q;
			wire [2:0] pmp_mseccfg_d;
			// Trace: design.sv:37726:5
			wire pmp_mseccfg_we;
			// Trace: design.sv:37727:5
			wire pmp_mseccfg_err;
			// Trace: design.sv:37728:5
			wire [5:0] pmp_cfg [0:PMPNumRegions - 1];
			// Trace: design.sv:37729:5
			wire [PMPNumRegions - 1:0] pmp_cfg_locked;
			// Trace: design.sv:37730:5
			reg [5:0] pmp_cfg_wdata [0:PMPNumRegions - 1];
			// Trace: design.sv:37731:5
			wire [PMPAddrWidth - 1:0] pmp_addr [0:PMPNumRegions - 1];
			// Trace: design.sv:37732:5
			wire [PMPNumRegions - 1:0] pmp_cfg_we;
			// Trace: design.sv:37733:5
			wire [PMPNumRegions - 1:0] pmp_cfg_err;
			// Trace: design.sv:37734:5
			wire [PMPNumRegions - 1:0] pmp_addr_we;
			// Trace: design.sv:37735:5
			wire [PMPNumRegions - 1:0] pmp_addr_err;
			// Trace: design.sv:37736:5
			wire any_pmp_entry_locked;
			genvar _gv_i_56;
			for (_gv_i_56 = 0; _gv_i_56 < ibex_pkg_PMP_MAX_REGIONS; _gv_i_56 = _gv_i_56 + 1) begin : g_exp_rd_data
				localparam i = _gv_i_56;
				if (i < PMPNumRegions) begin : g_implemented_regions
					// Trace: design.sv:37742:9
					assign pmp_cfg_rdata[i] = {pmp_cfg[i][5], 2'b00, pmp_cfg[i][4-:2], pmp_cfg[i][2], pmp_cfg[i][1], pmp_cfg[i][0]};
					if (PMPGranularity == 0) begin : g_pmp_g0
						// Trace: design.sv:37749:11
						wire [32:1] sv2v_tmp_2683A;
						assign sv2v_tmp_2683A = pmp_addr[i];
						always @(*) pmp_addr_rdata[i] = sv2v_tmp_2683A;
					end
					else if (PMPGranularity == 1) begin : g_pmp_g1
						// Trace: design.sv:37753:11
						always @(*) begin
							if (_sv2v_0)
								;
							// Trace: design.sv:37754:13
							pmp_addr_rdata[i] = pmp_addr[i];
							// Trace: design.sv:37755:13
							if ((pmp_cfg[i][4-:2] == 2'b00) || (pmp_cfg[i][4-:2] == 2'b01))
								// Trace: design.sv:37756:15
								pmp_addr_rdata[i][PMPGranularity - 1:0] = 1'sb0;
						end
					end
					else begin : g_pmp_g2
						// Trace: design.sv:37762:11
						always @(*) begin
							if (_sv2v_0)
								;
							// Trace: design.sv:37764:13
							pmp_addr_rdata[i] = {pmp_addr[i], {PMPGranularity - 1 {1'b1}}};
							// Trace: design.sv:37766:13
							if ((pmp_cfg[i][4-:2] == 2'b00) || (pmp_cfg[i][4-:2] == 2'b01))
								// Trace: design.sv:37768:15
								pmp_addr_rdata[i][PMPGranularity - 1:0] = 1'sb0;
						end
					end
				end
				else begin : g_other_regions
					// Trace: design.sv:37775:9
					assign pmp_cfg_rdata[i] = 1'sb0;
					// Trace: design.sv:37776:9
					wire [32:1] sv2v_tmp_D50E5;
					assign sv2v_tmp_D50E5 = 1'sb0;
					always @(*) pmp_addr_rdata[i] = sv2v_tmp_D50E5;
				end
			end
			genvar _gv_i_57;
			for (_gv_i_57 = 0; _gv_i_57 < PMPNumRegions; _gv_i_57 = _gv_i_57 + 1) begin : g_pmp_csrs
				localparam i = _gv_i_57;
				// Trace: design.sv:37785:7
				assign pmp_cfg_we[i] = (csr_we_int & ~pmp_cfg_locked[i]) & (csr_addr == (ibex_pkg_CSR_OFF_PMP_CFG + (i[11:0] >> 2)));
				// Trace: design.sv:37789:7
				wire [1:1] sv2v_tmp_8F287;
				assign sv2v_tmp_8F287 = csr_wdata_int[((i % 4) * ibex_pkg_PMP_CFG_W) + 7];
				always @(*) pmp_cfg_wdata[i][5] = sv2v_tmp_8F287;
				// Trace: design.sv:37791:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:37792:9
					(* full_case, parallel_case *)
					case (csr_wdata_int[((i % 4) * ibex_pkg_PMP_CFG_W) + 3+:2])
						2'b00:
							// Trace: design.sv:37793:21
							pmp_cfg_wdata[i][4-:2] = 2'b00;
						2'b01:
							// Trace: design.sv:37794:21
							pmp_cfg_wdata[i][4-:2] = 2'b01;
						2'b10:
							// Trace: design.sv:37795:21
							pmp_cfg_wdata[i][4-:2] = (PMPGranularity == 0 ? 2'b10 : 2'b00);
						2'b11:
							// Trace: design.sv:37797:21
							pmp_cfg_wdata[i][4-:2] = 2'b11;
						default:
							// Trace: design.sv:37798:21
							pmp_cfg_wdata[i][4-:2] = 2'b00;
					endcase
				end
				// Trace: design.sv:37801:7
				wire [1:1] sv2v_tmp_45785;
				assign sv2v_tmp_45785 = csr_wdata_int[((i % 4) * ibex_pkg_PMP_CFG_W) + 2];
				always @(*) pmp_cfg_wdata[i][2] = sv2v_tmp_45785;
				// Trace: design.sv:37804:7
				wire [1:1] sv2v_tmp_BB30C;
				assign sv2v_tmp_BB30C = (pmp_mseccfg_q[0] ? csr_wdata_int[((i % 4) * ibex_pkg_PMP_CFG_W) + 1] : &csr_wdata_int[(i % 4) * ibex_pkg_PMP_CFG_W+:2]);
				always @(*) pmp_cfg_wdata[i][1] = sv2v_tmp_BB30C;
				// Trace: design.sv:37806:7
				wire [1:1] sv2v_tmp_F1349;
				assign sv2v_tmp_F1349 = csr_wdata_int[(i % 4) * ibex_pkg_PMP_CFG_W];
				always @(*) pmp_cfg_wdata[i][0] = sv2v_tmp_F1349;
				// Trace: design.sv:37808:7
				ibex_csr #(
					.Width(6),
					.ShadowCopy(ShadowCSR),
					.ResetValue(pmp_cfg_rst[(15 - i) * 6+:6])
				) u_pmp_cfg_csr(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.wr_data_i({pmp_cfg_wdata[i]}),
					.wr_en_i(pmp_cfg_we[i]),
					.rd_data_o(pmp_cfg[i]),
					.rd_error_o(pmp_cfg_err[i])
				);
				// Trace: design.sv:37823:7
				assign pmp_cfg_locked[i] = pmp_cfg[i][5] & ~pmp_mseccfg_q[2];
				if (i < (PMPNumRegions - 1)) begin : g_lower
					// Trace: design.sv:37829:9
					assign pmp_addr_we[i] = ((csr_we_int & ~pmp_cfg_locked[i]) & (~pmp_cfg_locked[i + 1] | (pmp_cfg[i + 1][4-:2] != 2'b01))) & (csr_addr == (ibex_pkg_CSR_OFF_PMP_ADDR + i[11:0]));
				end
				else begin : g_upper
					// Trace: design.sv:37833:9
					assign pmp_addr_we[i] = (csr_we_int & ~pmp_cfg_locked[i]) & (csr_addr == (ibex_pkg_CSR_OFF_PMP_ADDR + i[11:0]));
				end
				// Trace: design.sv:37837:7
				ibex_csr #(
					.Width(PMPAddrWidth),
					.ShadowCopy(ShadowCSR),
					.ResetValue(pmp_addr_rst[((15 - i) * 34) + 33-:PMPAddrWidth])
				) u_pmp_addr_csr(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.wr_data_i(csr_wdata_int[31-:PMPAddrWidth]),
					.wr_en_i(pmp_addr_we[i]),
					.rd_data_o(pmp_addr[i]),
					.rd_error_o(pmp_addr_err[i])
				);
				// Trace: design.sv:37852:7
				assign csr_pmp_cfg_o[((PMPNumRegions - 1) - i) * 6+:6] = pmp_cfg[i];
				// Trace: design.sv:37853:7
				assign csr_pmp_addr_o[((PMPNumRegions - 1) - i) * 34+:34] = {pmp_addr_rdata[i], 2'b00};
			end
			// Trace: design.sv:37856:5
			assign pmp_mseccfg_we = csr_we_int & (csr_addr == 12'h747);
			// Trace: design.sv:37859:5
			assign pmp_mseccfg_d[0] = (pmp_mseccfg_q[0] ? 1'b1 : csr_wdata_int[ibex_pkg_CSR_MSECCFG_MML_BIT]);
			// Trace: design.sv:37860:5
			assign pmp_mseccfg_d[1] = (pmp_mseccfg_q[1] ? 1'b1 : csr_wdata_int[ibex_pkg_CSR_MSECCFG_MMWP_BIT]);
			// Trace: design.sv:37864:5
			assign any_pmp_entry_locked = |pmp_cfg_locked;
			// Trace: design.sv:37868:5
			assign pmp_mseccfg_d[2] = (any_pmp_entry_locked ? 1'b0 : csr_wdata_int[ibex_pkg_CSR_MSECCFG_RLB_BIT]);
			// Trace: design.sv:37870:5
			ibex_csr #(
				.Width(3),
				.ShadowCopy(ShadowCSR),
				.ResetValue(pmp_mseccfg_rst)
			) u_pmp_mseccfg(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.wr_data_i(pmp_mseccfg_d),
				.wr_en_i(pmp_mseccfg_we),
				.rd_data_o(pmp_mseccfg_q),
				.rd_error_o(pmp_mseccfg_err)
			);
			// Trace: design.sv:37883:5
			assign pmp_csr_err = (|pmp_cfg_err | (|pmp_addr_err)) | pmp_mseccfg_err;
			// Trace: design.sv:37884:5
			assign pmp_mseccfg = pmp_mseccfg_q;
		end
		else begin : g_no_pmp_tieoffs
			genvar _gv_i_58;
			for (_gv_i_58 = 0; _gv_i_58 < ibex_pkg_PMP_MAX_REGIONS; _gv_i_58 = _gv_i_58 + 1) begin : g_rdata
				localparam i = _gv_i_58;
				// Trace: design.sv:37889:7
				wire [32:1] sv2v_tmp_D50E5;
				assign sv2v_tmp_D50E5 = 1'sb0;
				always @(*) pmp_addr_rdata[i] = sv2v_tmp_D50E5;
				// Trace: design.sv:37890:7
				assign pmp_cfg_rdata[i] = 1'sb0;
			end
			genvar _gv_i_59;
			for (_gv_i_59 = 0; _gv_i_59 < PMPNumRegions; _gv_i_59 = _gv_i_59 + 1) begin : g_outputs
				localparam i = _gv_i_59;
				// Trace: design.sv:37893:7
				assign csr_pmp_cfg_o[((PMPNumRegions - 1) - i) * 6+:6] = 6'b000000;
				// Trace: design.sv:37894:7
				assign csr_pmp_addr_o[((PMPNumRegions - 1) - i) * 34+:34] = 1'sb0;
			end
			// Trace: design.sv:37896:5
			assign pmp_csr_err = 1'b0;
			// Trace: design.sv:37897:5
			assign pmp_mseccfg = 1'sb0;
		end
	endgenerate
	// Trace: design.sv:37900:3
	assign csr_pmp_mseccfg_o = pmp_mseccfg;
	// Trace: design.sv:37907:3
	always @(*) begin : mcountinhibit_update
		if (_sv2v_0)
			;
		// Trace: design.sv:37908:5
		if (mcountinhibit_we == 1'b1)
			// Trace: design.sv:37910:7
			mcountinhibit_d = {csr_wdata_int[MHPMCounterNum + 2:2], 1'b0, csr_wdata_int[0]};
		else
			// Trace: design.sv:37912:7
			mcountinhibit_d = mcountinhibit_q;
	end
	// Trace: design.sv:37917:3
	always @(*) begin : gen_mhpmcounter_incr
		if (_sv2v_0)
			;
		// Trace: design.sv:37920:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:37920:10
			reg [31:0] i;
			// Trace: design.sv:37920:10
			for (i = 0; i < 32; i = i + 1)
				begin : gen_mhpmcounter_incr_inactive
					// Trace: design.sv:37921:7
					mhpmcounter_incr[i] = 1'b0;
				end
		end
		// Trace: design.sv:37929:5
		mhpmcounter_incr[0] = 1'b1;
		// Trace: design.sv:37930:5
		mhpmcounter_incr[1] = 1'b0;
		// Trace: design.sv:37931:5
		mhpmcounter_incr[2] = instr_ret_i;
		// Trace: design.sv:37932:5
		mhpmcounter_incr[3] = dside_wait_i;
		// Trace: design.sv:37933:5
		mhpmcounter_incr[4] = iside_wait_i;
		// Trace: design.sv:37934:5
		mhpmcounter_incr[5] = mem_load_i;
		// Trace: design.sv:37935:5
		mhpmcounter_incr[6] = mem_store_i;
		// Trace: design.sv:37936:5
		mhpmcounter_incr[7] = jump_i;
		// Trace: design.sv:37937:5
		mhpmcounter_incr[8] = branch_i;
		// Trace: design.sv:37938:5
		mhpmcounter_incr[9] = branch_taken_i;
		// Trace: design.sv:37939:5
		mhpmcounter_incr[10] = instr_ret_compressed_i;
		// Trace: design.sv:37940:5
		mhpmcounter_incr[11] = mul_wait_i;
		// Trace: design.sv:37941:5
		mhpmcounter_incr[12] = div_wait_i;
	end
	// Trace: design.sv:37945:3
	always @(*) begin : gen_mhpmevent
		if (_sv2v_0)
			;
		// Trace: design.sv:37948:5
		begin : sv2v_autoblock_2
			// Trace: design.sv:37948:10
			reg signed [31:0] i;
			// Trace: design.sv:37948:10
			for (i = 0; i < 32; i = i + 1)
				begin : gen_mhpmevent_active
					// Trace: design.sv:37949:7
					mhpmevent[i] = 1'sb0;
					// Trace: design.sv:37950:7
					mhpmevent[i][i] = 1'b1;
				end
		end
		// Trace: design.sv:37954:5
		mhpmevent[1] = 1'sb0;
		begin : sv2v_autoblock_3
			// Trace: design.sv:37955:10
			reg [31:0] i;
			// Trace: design.sv:37955:10
			for (i = 3 + MHPMCounterNum; i < 32; i = i + 1)
				begin : gen_mhpmevent_inactive
					// Trace: design.sv:37956:7
					mhpmevent[i] = 1'sb0;
				end
		end
	end
	// Trace: design.sv:37961:3
	ibex_counter #(.CounterWidth(64)) mcycle_counter_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.counter_inc_i(mhpmcounter_incr[0] & ~mcountinhibit[0]),
		.counterh_we_i(mhpmcounterh_we[0]),
		.counter_we_i(mhpmcounter_we[0]),
		.counter_val_i(csr_wdata_int),
		.counter_val_o(mhpmcounter[0]),
		.counter_val_upd_o()
	);
	// Trace: design.sv:37976:3
	ibex_counter #(
		.CounterWidth(64),
		.ProvideValUpd(1)
	) minstret_counter_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.counter_inc_i(mhpmcounter_incr[2] & ~mcountinhibit[2]),
		.counterh_we_i(mhpmcounterh_we[2]),
		.counter_we_i(mhpmcounter_we[2]),
		.counter_val_i(csr_wdata_int),
		.counter_val_o(minstret_raw),
		.counter_val_upd_o(minstret_next)
	);
	// Trace: design.sv:37997:3
	assign mhpmcounter[2] = (instr_ret_spec_i & ~mcountinhibit[2] ? minstret_next : minstret_raw);
	// Trace: design.sv:38000:3
	assign mhpmcounter[1] = 1'sb0;
	// Trace: design.sv:38001:3
	assign unused_mhpmcounter_we_1 = mhpmcounter_we[1];
	// Trace: design.sv:38002:3
	assign unused_mhpmcounterh_we_1 = mhpmcounterh_we[1];
	// Trace: design.sv:38003:3
	assign unused_mhpmcounter_incr_1 = mhpmcounter_incr[1];
	// Trace: design.sv:38006:3
	genvar _gv_i_60;
	generate
		for (_gv_i_60 = 0; _gv_i_60 < 29; _gv_i_60 = _gv_i_60 + 1) begin : gen_cntrs
			localparam i = _gv_i_60;
			// Trace: design.sv:38007:5
			localparam signed [31:0] Cnt = i + 3;
			if (i < MHPMCounterNum) begin : gen_imp
				// Trace: design.sv:38010:7
				wire [63:0] mhpmcounter_raw;
				wire [63:0] mhpmcounter_next;
				// Trace: design.sv:38012:7
				ibex_counter #(
					.CounterWidth(MHPMCounterWidth),
					.ProvideValUpd(Cnt == 10)
				) mcounters_variable_i(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.counter_inc_i(mhpmcounter_incr[Cnt] & ~mcountinhibit[Cnt]),
					.counterh_we_i(mhpmcounterh_we[Cnt]),
					.counter_we_i(mhpmcounter_we[Cnt]),
					.counter_val_i(csr_wdata_int),
					.counter_val_o(mhpmcounter_raw),
					.counter_val_upd_o(mhpmcounter_next)
				);
				if (Cnt == 10) begin : gen_compressed_instr_cnt
					// Trace: design.sv:38029:9
					assign mhpmcounter[Cnt] = (instr_ret_compressed_spec_i & ~mcountinhibit[Cnt] ? mhpmcounter_next : mhpmcounter_raw);
				end
				else begin : gen_other_cnts
					// Trace: design.sv:38033:9
					wire [63:0] unused_mhpmcounter_next;
					// Trace: design.sv:38035:9
					assign mhpmcounter[Cnt] = mhpmcounter_raw;
					// Trace: design.sv:38036:9
					assign unused_mhpmcounter_next = mhpmcounter_next;
				end
			end
			else begin : gen_unimp
				// Trace: design.sv:38039:7
				assign mhpmcounter[Cnt] = 1'sb0;
				if (Cnt == 10) begin : gen_no_compressed_instr_cnt
					// Trace: design.sv:38042:9
					wire unused_instr_ret_compressed_spec_i;
					// Trace: design.sv:38043:9
					assign unused_instr_ret_compressed_spec_i = instr_ret_compressed_spec_i;
				end
			end
		end
	endgenerate
	// Trace: design.sv:38048:3
	generate
		if (MHPMCounterNum < 29) begin : g_mcountinhibit_reduced
			// Trace: design.sv:38049:5
			wire [(29 - MHPMCounterNum) - 1:0] unused_mhphcounter_we;
			// Trace: design.sv:38050:5
			wire [(29 - MHPMCounterNum) - 1:0] unused_mhphcounterh_we;
			// Trace: design.sv:38051:5
			wire [(29 - MHPMCounterNum) - 1:0] unused_mhphcounter_incr;
			// Trace: design.sv:38053:5
			assign mcountinhibit = {{29 - MHPMCounterNum {1'b1}}, mcountinhibit_q};
			// Trace: design.sv:38055:5
			assign unused_mhphcounter_we = mhpmcounter_we[31:MHPMCounterNum + 3];
			// Trace: design.sv:38056:5
			assign unused_mhphcounterh_we = mhpmcounterh_we[31:MHPMCounterNum + 3];
			// Trace: design.sv:38057:5
			assign unused_mhphcounter_incr = mhpmcounter_incr[31:MHPMCounterNum + 3];
		end
		else begin : g_mcountinhibit_full
			// Trace: design.sv:38059:5
			assign mcountinhibit = mcountinhibit_q;
		end
	endgenerate
	// Trace: design.sv:38062:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:38063:5
		if (!rst_ni)
			// Trace: design.sv:38064:7
			mcountinhibit_q <= 1'sb0;
		else
			// Trace: design.sv:38066:7
			mcountinhibit_q <= mcountinhibit_d;
	// Trace: design.sv:38074:3
	generate
		if (DbgTriggerEn) begin : gen_trigger_regs
			// Trace: design.sv:38075:5
			localparam [31:0] DbgHwNumLen = (DbgHwBreakNum > 1 ? $clog2(DbgHwBreakNum) : 1);
			// Trace: design.sv:38076:5
			localparam [31:0] MaxTselect = DbgHwBreakNum - 1;
			// Trace: design.sv:38079:5
			wire [DbgHwNumLen - 1:0] tselect_d;
			wire [DbgHwNumLen - 1:0] tselect_q;
			// Trace: design.sv:38080:5
			wire tmatch_control_d;
			// Trace: design.sv:38081:5
			wire [DbgHwBreakNum - 1:0] tmatch_control_q;
			// Trace: design.sv:38082:5
			wire [31:0] tmatch_value_d;
			// Trace: design.sv:38083:5
			wire [31:0] tmatch_value_q [0:DbgHwBreakNum - 1];
			// Trace: design.sv:38084:5
			wire selected_tmatch_control;
			// Trace: design.sv:38085:5
			wire [31:0] selected_tmatch_value;
			// Trace: design.sv:38088:5
			wire tselect_we;
			// Trace: design.sv:38089:5
			wire [DbgHwBreakNum - 1:0] tmatch_control_we;
			// Trace: design.sv:38090:5
			wire [DbgHwBreakNum - 1:0] tmatch_value_we;
			// Trace: design.sv:38092:5
			wire [DbgHwBreakNum - 1:0] trigger_match;
			// Trace: design.sv:38095:5
			assign tselect_we = (csr_we_int & debug_mode_i) & (csr_addr_i == 12'h7a0);
			genvar _gv_i_61;
			for (_gv_i_61 = 0; _gv_i_61 < DbgHwBreakNum; _gv_i_61 = _gv_i_61 + 1) begin : g_dbg_tmatch_we
				localparam i = _gv_i_61;
				// Trace: design.sv:38097:7
				assign tmatch_control_we[i] = (((i[DbgHwNumLen - 1:0] == tselect_q) & csr_we_int) & debug_mode_i) & (csr_addr_i == 12'h7a1);
				// Trace: design.sv:38099:7
				assign tmatch_value_we[i] = (((i[DbgHwNumLen - 1:0] == tselect_q) & csr_we_int) & debug_mode_i) & (csr_addr_i == 12'h7a2);
			end
			// Trace: design.sv:38105:5
			assign tselect_d = (csr_wdata_int < DbgHwBreakNum ? csr_wdata_int[DbgHwNumLen - 1:0] : MaxTselect[DbgHwNumLen - 1:0]);
			// Trace: design.sv:38109:5
			assign tmatch_control_d = csr_wdata_int[2];
			// Trace: design.sv:38110:5
			assign tmatch_value_d = csr_wdata_int[31:0];
			// Trace: design.sv:38113:5
			ibex_csr #(
				.Width(DbgHwNumLen),
				.ShadowCopy(1'b0),
				.ResetValue(1'sb0)
			) u_tselect_csr(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.wr_data_i(tselect_d),
				.wr_en_i(tselect_we),
				.rd_data_o(tselect_q),
				.rd_error_o()
			);
			genvar _gv_i_62;
			for (_gv_i_62 = 0; _gv_i_62 < DbgHwBreakNum; _gv_i_62 = _gv_i_62 + 1) begin : g_dbg_tmatch_reg
				localparam i = _gv_i_62;
				// Trace: design.sv:38127:7
				ibex_csr #(
					.Width(1),
					.ShadowCopy(1'b0),
					.ResetValue(1'sb0)
				) u_tmatch_control_csr(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.wr_data_i(tmatch_control_d),
					.wr_en_i(tmatch_control_we[i]),
					.rd_data_o(tmatch_control_q[i]),
					.rd_error_o()
				);
				// Trace: design.sv:38140:7
				ibex_csr #(
					.Width(32),
					.ShadowCopy(1'b0),
					.ResetValue(1'sb0)
				) u_tmatch_value_csr(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.wr_data_i(tmatch_value_d),
					.wr_en_i(tmatch_value_we[i]),
					.rd_data_o(tmatch_value_q[i]),
					.rd_error_o()
				);
			end
			// Trace: design.sv:38156:5
			localparam [31:0] TSelectRdataPadlen = (DbgHwNumLen >= 32 ? 0 : 32 - DbgHwNumLen);
			// Trace: design.sv:38157:5
			assign tselect_rdata = {{TSelectRdataPadlen {1'b0}}, tselect_q};
			if (DbgHwBreakNum > 1) begin : g_dbg_tmatch_multiple_select
				// Trace: design.sv:38160:7
				assign selected_tmatch_control = tmatch_control_q[tselect_q];
				// Trace: design.sv:38161:7
				assign selected_tmatch_value = tmatch_value_q[tselect_q];
			end
			else begin : g_dbg_tmatch_single_select
				// Trace: design.sv:38163:7
				assign selected_tmatch_control = tmatch_control_q[0];
				// Trace: design.sv:38164:7
				assign selected_tmatch_value = tmatch_value_q[0];
			end
			// Trace: design.sv:38168:5
			assign tmatch_control_rdata = {29'h05000209, selected_tmatch_control, 2'b00};
			// Trace: design.sv:38187:5
			assign tmatch_value_rdata = selected_tmatch_value;
			genvar _gv_i_63;
			for (_gv_i_63 = 0; _gv_i_63 < DbgHwBreakNum; _gv_i_63 = _gv_i_63 + 1) begin : g_dbg_trigger_match
				localparam i = _gv_i_63;
				// Trace: design.sv:38192:7
				assign trigger_match[i] = tmatch_control_q[i] & (pc_if_i[31:0] == tmatch_value_q[i]);
			end
			// Trace: design.sv:38194:5
			assign trigger_match_o = |trigger_match;
		end
		else begin : gen_no_trigger_regs
			// Trace: design.sv:38197:5
			assign tselect_rdata = 'b0;
			// Trace: design.sv:38198:5
			assign tmatch_control_rdata = 'b0;
			// Trace: design.sv:38199:5
			assign tmatch_value_rdata = 'b0;
			// Trace: design.sv:38200:5
			assign trigger_match_o = 'b0;
		end
	endgenerate
	// Trace: design.sv:38208:3
	assign cpuctrl_wdata_raw = csr_wdata_int[7:0];
	// Trace: design.sv:38211:3
	generate
		if (DataIndTiming) begin : gen_dit
			// Trace: design.sv:38213:5
			assign cpuctrl_wdata[1] = cpuctrl_wdata_raw[1];
		end
		else begin : gen_no_dit
			// Trace: design.sv:38217:5
			wire unused_dit;
			// Trace: design.sv:38218:5
			assign unused_dit = cpuctrl_wdata_raw[1];
			// Trace: design.sv:38221:5
			assign cpuctrl_wdata[1] = 1'b0;
		end
	endgenerate
	// Trace: design.sv:38224:3
	assign data_ind_timing_o = cpuctrl_q[1];
	// Trace: design.sv:38227:3
	generate
		if (DummyInstructions) begin : gen_dummy
			// Trace: design.sv:38229:5
			assign cpuctrl_wdata[2] = cpuctrl_wdata_raw[2];
			// Trace: design.sv:38230:5
			assign cpuctrl_wdata[5-:3] = cpuctrl_wdata_raw[5-:3];
			// Trace: design.sv:38233:5
			assign dummy_instr_seed_en_o = csr_we_int && (csr_addr == 12'h7c1);
			// Trace: design.sv:38234:5
			assign dummy_instr_seed_o = csr_wdata_int;
		end
		else begin : gen_no_dummy
			// Trace: design.sv:38238:5
			wire unused_dummy_en;
			// Trace: design.sv:38239:5
			wire [2:0] unused_dummy_mask;
			// Trace: design.sv:38240:5
			assign unused_dummy_en = cpuctrl_wdata_raw[2];
			// Trace: design.sv:38241:5
			assign unused_dummy_mask = cpuctrl_wdata_raw[5-:3];
			// Trace: design.sv:38244:5
			assign cpuctrl_wdata[2] = 1'b0;
			// Trace: design.sv:38245:5
			assign cpuctrl_wdata[5-:3] = 3'b000;
			// Trace: design.sv:38246:5
			assign dummy_instr_seed_en_o = 1'b0;
			// Trace: design.sv:38247:5
			assign dummy_instr_seed_o = 1'sb0;
		end
	endgenerate
	// Trace: design.sv:38250:3
	assign dummy_instr_en_o = cpuctrl_q[2];
	// Trace: design.sv:38251:3
	assign dummy_instr_mask_o = cpuctrl_q[5-:3];
	// Trace: design.sv:38254:3
	generate
		if (ICache) begin : gen_icache_enable
			// Trace: design.sv:38255:5
			assign cpuctrl_wdata[0] = cpuctrl_wdata_raw[0];
		end
		else begin : gen_no_icache
			// Trace: design.sv:38258:5
			wire unused_icen;
			// Trace: design.sv:38259:5
			assign unused_icen = cpuctrl_wdata_raw[0];
			// Trace: design.sv:38262:5
			assign cpuctrl_wdata[0] = 1'b0;
		end
	endgenerate
	// Trace: design.sv:38265:3
	assign cpuctrl_wdata[7] = cpuctrl_wdata_raw[7];
	// Trace: design.sv:38266:3
	assign cpuctrl_wdata[6] = cpuctrl_wdata_raw[6];
	// Trace: design.sv:38268:3
	assign icache_enable_o = cpuctrl_q[0];
	// Trace: design.sv:38270:3
	ibex_csr #(
		.Width(8),
		.ShadowCopy(ShadowCSR),
		.ResetValue(1'sb0)
	) u_cpuctrl_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({cpuctrl_d}),
		.wr_en_i(cpuctrl_we),
		.rd_data_o(cpuctrl_q),
		.rd_error_o(cpuctrl_err)
	);
	// Trace: design.sv:38283:3
	assign csr_shadow_err_o = ((mstatus_err | mtvec_err) | pmp_csr_err) | cpuctrl_err;
	initial _sv2v_0 = 0;
endmodule
module ibex_csr (
	clk_i,
	rst_ni,
	wr_data_i,
	wr_en_i,
	rd_data_o,
	rd_error_o
);
	// Trace: design.sv:38303:13
	parameter [31:0] Width = 32;
	// Trace: design.sv:38304:13
	parameter [0:0] ShadowCopy = 1'b0;
	// Trace: design.sv:38305:13
	parameter [Width - 1:0] ResetValue = 1'sb0;
	// Trace: design.sv:38307:3
	input wire clk_i;
	// Trace: design.sv:38308:3
	input wire rst_ni;
	// Trace: design.sv:38310:3
	input wire [Width - 1:0] wr_data_i;
	// Trace: design.sv:38311:3
	input wire wr_en_i;
	// Trace: design.sv:38312:3
	output wire [Width - 1:0] rd_data_o;
	// Trace: design.sv:38314:3
	output wire rd_error_o;
	// Trace: design.sv:38317:3
	reg [Width - 1:0] rdata_q;
	// Trace: design.sv:38319:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:38320:5
		if (!rst_ni)
			// Trace: design.sv:38321:7
			rdata_q <= ResetValue;
		else if (wr_en_i)
			// Trace: design.sv:38323:7
			rdata_q <= wr_data_i;
	// Trace: design.sv:38327:3
	assign rd_data_o = rdata_q;
	// Trace: design.sv:38329:3
	generate
		if (ShadowCopy) begin : gen_shadow
			// Trace: design.sv:38330:5
			reg [Width - 1:0] shadow_q;
			// Trace: design.sv:38332:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:38333:7
				if (!rst_ni)
					// Trace: design.sv:38334:9
					shadow_q <= ~ResetValue;
				else if (wr_en_i)
					// Trace: design.sv:38336:9
					shadow_q <= ~wr_data_i;
			// Trace: design.sv:38340:5
			assign rd_error_o = rdata_q != ~shadow_q;
		end
		else begin : gen_no_shadow
			// Trace: design.sv:38343:5
			assign rd_error_o = 1'b0;
		end
	endgenerate
endmodule
module ibex_counter (
	clk_i,
	rst_ni,
	counter_inc_i,
	counterh_we_i,
	counter_we_i,
	counter_val_i,
	counter_val_o,
	counter_val_upd_o
);
	reg _sv2v_0;
	// Trace: design.sv:38350:13
	parameter signed [31:0] CounterWidth = 32;
	// Trace: design.sv:38354:13
	parameter [0:0] ProvideValUpd = 0;
	// Trace: design.sv:38356:3
	input wire clk_i;
	// Trace: design.sv:38357:3
	input wire rst_ni;
	// Trace: design.sv:38359:3
	input wire counter_inc_i;
	// Trace: design.sv:38360:3
	input wire counterh_we_i;
	// Trace: design.sv:38361:3
	input wire counter_we_i;
	// Trace: design.sv:38362:3
	input wire [31:0] counter_val_i;
	// Trace: design.sv:38363:3
	output wire [63:0] counter_val_o;
	// Trace: design.sv:38364:3
	output wire [63:0] counter_val_upd_o;
	// Trace: design.sv:38367:3
	wire [63:0] counter;
	// Trace: design.sv:38368:3
	wire [CounterWidth - 1:0] counter_upd;
	// Trace: design.sv:38369:3
	reg [63:0] counter_load;
	// Trace: design.sv:38370:3
	reg we;
	// Trace: design.sv:38371:3
	reg [CounterWidth - 1:0] counter_d;
	// Trace: design.sv:38374:3
	assign counter_upd = counter[CounterWidth - 1:0] + {{CounterWidth - 1 {1'b0}}, 1'b1};
	// Trace: design.sv:38377:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:38379:5
		we = counter_we_i | counterh_we_i;
		// Trace: design.sv:38380:5
		counter_load[63:32] = counter[63:32];
		// Trace: design.sv:38381:5
		counter_load[31:0] = counter_val_i;
		// Trace: design.sv:38382:5
		if (counterh_we_i) begin
			// Trace: design.sv:38383:7
			counter_load[63:32] = counter_val_i;
			// Trace: design.sv:38384:7
			counter_load[31:0] = counter[31:0];
		end
		if (we)
			// Trace: design.sv:38389:7
			counter_d = counter_load[CounterWidth - 1:0];
		else if (counter_inc_i)
			// Trace: design.sv:38391:7
			counter_d = counter_upd[CounterWidth - 1:0];
		else
			// Trace: design.sv:38393:7
			counter_d = counter[CounterWidth - 1:0];
	end
	// Trace: design.sv:38405:3
	reg [CounterWidth - 1:0] counter_q;
	// Trace: design.sv:38411:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:38412:5
		if (!rst_ni)
			// Trace: design.sv:38413:7
			counter_q <= 1'sb0;
		else
			// Trace: design.sv:38415:7
			counter_q <= counter_d;
	// Trace: design.sv:38419:3
	generate
		if (CounterWidth < 64) begin : g_counter_narrow
			// Trace: design.sv:38420:5
			wire [63:CounterWidth] unused_counter_load;
			// Trace: design.sv:38422:5
			assign counter[CounterWidth - 1:0] = counter_q;
			// Trace: design.sv:38423:5
			assign counter[63:CounterWidth] = 1'sb0;
			if (ProvideValUpd) begin : g_counter_val_upd_o
				// Trace: design.sv:38426:7
				assign counter_val_upd_o[CounterWidth - 1:0] = counter_upd;
			end
			else begin : g_no_counter_val_upd_o
				// Trace: design.sv:38428:7
				assign counter_val_upd_o[CounterWidth - 1:0] = 1'sb0;
			end
			// Trace: design.sv:38430:5
			assign counter_val_upd_o[63:CounterWidth] = 1'sb0;
			// Trace: design.sv:38431:5
			assign unused_counter_load = counter_load[63:CounterWidth];
		end
		else begin : g_counter_full
			// Trace: design.sv:38433:5
			assign counter = counter_q;
			if (ProvideValUpd) begin : g_counter_val_upd_o
				// Trace: design.sv:38436:7
				assign counter_val_upd_o = counter_upd;
			end
			else begin : g_no_counter_val_upd_o
				// Trace: design.sv:38438:7
				assign counter_val_upd_o = 1'sb0;
			end
		end
	endgenerate
	// Trace: design.sv:38442:3
	assign counter_val_o = counter;
	initial _sv2v_0 = 0;
endmodule
module ibex_decoder (
	clk_i,
	rst_ni,
	illegal_insn_o,
	ebrk_insn_o,
	mret_insn_o,
	dret_insn_o,
	ecall_insn_o,
	wfi_insn_o,
	jump_set_o,
	branch_taken_i,
	icache_inval_o,
	instr_first_cycle_i,
	instr_rdata_i,
	instr_rdata_alu_i,
	illegal_c_insn_i,
	imm_a_mux_sel_o,
	imm_b_mux_sel_o,
	bt_a_mux_sel_o,
	bt_b_mux_sel_o,
	imm_i_type_o,
	imm_s_type_o,
	imm_b_type_o,
	imm_u_type_o,
	imm_j_type_o,
	zimm_rs1_type_o,
	rf_wdata_sel_o,
	rf_we_o,
	rf_raddr_a_o,
	rf_raddr_b_o,
	rf_waddr_o,
	rf_ren_a_o,
	rf_ren_b_o,
	alu_operator_o,
	alu_op_a_mux_sel_o,
	alu_op_b_mux_sel_o,
	alu_multicycle_o,
	mult_en_o,
	div_en_o,
	mult_sel_o,
	div_sel_o,
	multdiv_operator_o,
	multdiv_signed_mode_o,
	csr_access_o,
	csr_op_o,
	data_req_o,
	data_we_o,
	data_type_o,
	data_sign_extension_o,
	jump_in_dec_o,
	branch_in_dec_o
);
	reg _sv2v_0;
	// Trace: design.sv:38464:13
	parameter [0:0] RV32E = 0;
	// Trace: design.sv:38465:13
	// removed localparam type ibex_pkg_rv32m_e
	parameter integer RV32M = 32'sd2;
	// Trace: design.sv:38466:13
	// removed localparam type ibex_pkg_rv32b_e
	parameter integer RV32B = 32'sd0;
	// Trace: design.sv:38467:13
	parameter [0:0] BranchTargetALU = 0;
	// Trace: design.sv:38469:3
	input wire clk_i;
	// Trace: design.sv:38470:3
	input wire rst_ni;
	// Trace: design.sv:38473:3
	output wire illegal_insn_o;
	// Trace: design.sv:38474:3
	output reg ebrk_insn_o;
	// Trace: design.sv:38475:3
	output reg mret_insn_o;
	// Trace: design.sv:38477:3
	output reg dret_insn_o;
	// Trace: design.sv:38478:3
	output reg ecall_insn_o;
	// Trace: design.sv:38479:3
	output reg wfi_insn_o;
	// Trace: design.sv:38480:3
	output reg jump_set_o;
	// Trace: design.sv:38481:3
	input wire branch_taken_i;
	// Trace: design.sv:38482:3
	output reg icache_inval_o;
	// Trace: design.sv:38485:3
	input wire instr_first_cycle_i;
	// Trace: design.sv:38486:3
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:38487:3
	input wire [31:0] instr_rdata_alu_i;
	// Trace: design.sv:38490:3
	input wire illegal_c_insn_i;
	// Trace: design.sv:38493:3
	// removed localparam type ibex_pkg_imm_a_sel_e
	output reg imm_a_mux_sel_o;
	// Trace: design.sv:38494:3
	// removed localparam type ibex_pkg_imm_b_sel_e
	output reg [2:0] imm_b_mux_sel_o;
	// Trace: design.sv:38495:3
	// removed localparam type ibex_pkg_op_a_sel_e
	output reg [1:0] bt_a_mux_sel_o;
	// Trace: design.sv:38496:3
	output reg [2:0] bt_b_mux_sel_o;
	// Trace: design.sv:38497:3
	output wire [31:0] imm_i_type_o;
	// Trace: design.sv:38498:3
	output wire [31:0] imm_s_type_o;
	// Trace: design.sv:38499:3
	output wire [31:0] imm_b_type_o;
	// Trace: design.sv:38500:3
	output wire [31:0] imm_u_type_o;
	// Trace: design.sv:38501:3
	output wire [31:0] imm_j_type_o;
	// Trace: design.sv:38502:3
	output wire [31:0] zimm_rs1_type_o;
	// Trace: design.sv:38505:3
	// removed localparam type ibex_pkg_rf_wd_sel_e
	output reg rf_wdata_sel_o;
	// Trace: design.sv:38506:3
	output wire rf_we_o;
	// Trace: design.sv:38507:3
	output wire [4:0] rf_raddr_a_o;
	// Trace: design.sv:38508:3
	output wire [4:0] rf_raddr_b_o;
	// Trace: design.sv:38509:3
	output wire [4:0] rf_waddr_o;
	// Trace: design.sv:38510:3
	output reg rf_ren_a_o;
	// Trace: design.sv:38511:3
	output reg rf_ren_b_o;
	// Trace: design.sv:38514:3
	// removed localparam type ibex_pkg_alu_op_e
	output reg [6:0] alu_operator_o;
	// Trace: design.sv:38515:3
	output reg [1:0] alu_op_a_mux_sel_o;
	// Trace: design.sv:38517:3
	// removed localparam type ibex_pkg_op_b_sel_e
	output reg alu_op_b_mux_sel_o;
	// Trace: design.sv:38519:3
	output reg alu_multicycle_o;
	// Trace: design.sv:38522:3
	output wire mult_en_o;
	// Trace: design.sv:38523:3
	output wire div_en_o;
	// Trace: design.sv:38524:3
	output reg mult_sel_o;
	// Trace: design.sv:38525:3
	output reg div_sel_o;
	// Trace: design.sv:38527:3
	// removed localparam type ibex_pkg_md_op_e
	output reg [1:0] multdiv_operator_o;
	// Trace: design.sv:38528:3
	output reg [1:0] multdiv_signed_mode_o;
	// Trace: design.sv:38531:3
	output reg csr_access_o;
	// Trace: design.sv:38532:3
	// removed localparam type ibex_pkg_csr_op_e
	output reg [1:0] csr_op_o;
	// Trace: design.sv:38535:3
	output reg data_req_o;
	// Trace: design.sv:38536:3
	output reg data_we_o;
	// Trace: design.sv:38537:3
	output reg [1:0] data_type_o;
	// Trace: design.sv:38539:3
	output reg data_sign_extension_o;
	// Trace: design.sv:38543:3
	output reg jump_in_dec_o;
	// Trace: design.sv:38544:3
	output reg branch_in_dec_o;
	// Trace: design.sv:38547:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:38549:3
	reg illegal_insn;
	// Trace: design.sv:38550:3
	wire illegal_reg_rv32e;
	// Trace: design.sv:38551:3
	reg csr_illegal;
	// Trace: design.sv:38552:3
	reg rf_we;
	// Trace: design.sv:38554:3
	wire [31:0] instr;
	// Trace: design.sv:38555:3
	wire [31:0] instr_alu;
	// Trace: design.sv:38556:3
	wire [9:0] unused_instr_alu;
	// Trace: design.sv:38558:3
	wire [4:0] instr_rs1;
	// Trace: design.sv:38559:3
	wire [4:0] instr_rs2;
	// Trace: design.sv:38560:3
	wire [4:0] instr_rs3;
	// Trace: design.sv:38561:3
	wire [4:0] instr_rd;
	// Trace: design.sv:38563:3
	reg use_rs3_d;
	// Trace: design.sv:38564:3
	reg use_rs3_q;
	// Trace: design.sv:38566:3
	reg [1:0] csr_op;
	// Trace: design.sv:38568:3
	// removed localparam type ibex_pkg_opcode_e
	reg [6:0] opcode;
	// Trace: design.sv:38569:3
	reg [6:0] opcode_alu;
	// Trace: design.sv:38574:3
	assign instr = instr_rdata_i;
	// Trace: design.sv:38575:3
	assign instr_alu = instr_rdata_alu_i;
	// Trace: design.sv:38582:3
	assign imm_i_type_o = {{20 {instr[31]}}, instr[31:20]};
	// Trace: design.sv:38583:3
	assign imm_s_type_o = {{20 {instr[31]}}, instr[31:25], instr[11:7]};
	// Trace: design.sv:38584:3
	assign imm_b_type_o = {{19 {instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
	// Trace: design.sv:38585:3
	assign imm_u_type_o = {instr[31:12], 12'b000000000000};
	// Trace: design.sv:38586:3
	assign imm_j_type_o = {{12 {instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};
	// Trace: design.sv:38589:3
	assign zimm_rs1_type_o = {27'b000000000000000000000000000, instr_rs1};
	// Trace: design.sv:38591:3
	generate
		if (RV32B != 32'sd0) begin : gen_rs3_flop
			// Trace: design.sv:38593:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:38594:7
				if (!rst_ni)
					// Trace: design.sv:38595:9
					use_rs3_q <= 1'b0;
				else
					// Trace: design.sv:38597:9
					use_rs3_q <= use_rs3_d;
		end
		else begin : gen_no_rs3_flop
			// Trace: design.sv:38601:5
			wire unused_clk;
			// Trace: design.sv:38602:5
			wire unused_rst_n;
			// Trace: design.sv:38605:5
			assign unused_clk = clk_i;
			// Trace: design.sv:38606:5
			assign unused_rst_n = rst_ni;
			// Trace: design.sv:38609:5
			wire [1:1] sv2v_tmp_12378;
			assign sv2v_tmp_12378 = use_rs3_d;
			always @(*) use_rs3_q = sv2v_tmp_12378;
		end
	endgenerate
	// Trace: design.sv:38613:3
	assign instr_rs1 = instr[19:15];
	// Trace: design.sv:38614:3
	assign instr_rs2 = instr[24:20];
	// Trace: design.sv:38615:3
	assign instr_rs3 = instr[31:27];
	// Trace: design.sv:38616:3
	assign rf_raddr_a_o = (use_rs3_q & ~instr_first_cycle_i ? instr_rs3 : instr_rs1);
	// Trace: design.sv:38617:3
	assign rf_raddr_b_o = instr_rs2;
	// Trace: design.sv:38620:3
	assign instr_rd = instr[11:7];
	// Trace: design.sv:38621:3
	assign rf_waddr_o = instr_rd;
	// Trace: design.sv:38626:3
	generate
		if (RV32E) begin : gen_rv32e_reg_check_active
			// Trace: design.sv:38627:5
			assign illegal_reg_rv32e = ((rf_raddr_a_o[4] & (alu_op_a_mux_sel_o == 2'd0)) | (rf_raddr_b_o[4] & (alu_op_b_mux_sel_o == 1'd0))) | (rf_waddr_o[4] & rf_we);
		end
		else begin : gen_rv32e_reg_check_inactive
			// Trace: design.sv:38631:5
			assign illegal_reg_rv32e = 1'b0;
		end
	endgenerate
	// Trace: design.sv:38637:3
	always @(*) begin : csr_operand_check
		if (_sv2v_0)
			;
		// Trace: design.sv:38638:5
		csr_op_o = csr_op;
		// Trace: design.sv:38642:5
		if (((csr_op == 2'd2) || (csr_op == 2'd3)) && (instr_rs1 == {5 {1'sb0}}))
			// Trace: design.sv:38644:7
			csr_op_o = 2'd0;
	end
	// Trace: design.sv:38652:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:38653:5
		jump_in_dec_o = 1'b0;
		// Trace: design.sv:38654:5
		jump_set_o = 1'b0;
		// Trace: design.sv:38655:5
		branch_in_dec_o = 1'b0;
		// Trace: design.sv:38656:5
		icache_inval_o = 1'b0;
		// Trace: design.sv:38658:5
		multdiv_operator_o = 2'd0;
		// Trace: design.sv:38659:5
		multdiv_signed_mode_o = 2'b00;
		// Trace: design.sv:38661:5
		rf_wdata_sel_o = 1'd0;
		// Trace: design.sv:38662:5
		rf_we = 1'b0;
		// Trace: design.sv:38663:5
		rf_ren_a_o = 1'b0;
		// Trace: design.sv:38664:5
		rf_ren_b_o = 1'b0;
		// Trace: design.sv:38666:5
		csr_access_o = 1'b0;
		// Trace: design.sv:38667:5
		csr_illegal = 1'b0;
		// Trace: design.sv:38668:5
		csr_op = 2'd0;
		// Trace: design.sv:38670:5
		data_we_o = 1'b0;
		// Trace: design.sv:38671:5
		data_type_o = 2'b00;
		// Trace: design.sv:38672:5
		data_sign_extension_o = 1'b0;
		// Trace: design.sv:38673:5
		data_req_o = 1'b0;
		// Trace: design.sv:38675:5
		illegal_insn = 1'b0;
		// Trace: design.sv:38676:5
		ebrk_insn_o = 1'b0;
		// Trace: design.sv:38677:5
		mret_insn_o = 1'b0;
		// Trace: design.sv:38678:5
		dret_insn_o = 1'b0;
		// Trace: design.sv:38679:5
		ecall_insn_o = 1'b0;
		// Trace: design.sv:38680:5
		wfi_insn_o = 1'b0;
		// Trace: design.sv:38682:5
		opcode = instr[6:0];
		// Trace: design.sv:38684:5
		(* full_case, parallel_case *)
		case (opcode)
			7'h6f: begin
				// Trace: design.sv:38691:9
				jump_in_dec_o = 1'b1;
				// Trace: design.sv:38693:9
				if (instr_first_cycle_i) begin
					// Trace: design.sv:38695:11
					rf_we = BranchTargetALU;
					// Trace: design.sv:38696:11
					jump_set_o = 1'b1;
				end
				else
					// Trace: design.sv:38699:11
					rf_we = 1'b1;
			end
			7'h67: begin
				// Trace: design.sv:38704:9
				jump_in_dec_o = 1'b1;
				// Trace: design.sv:38706:9
				if (instr_first_cycle_i) begin
					// Trace: design.sv:38708:11
					rf_we = BranchTargetALU;
					// Trace: design.sv:38709:11
					jump_set_o = 1'b1;
				end
				else
					// Trace: design.sv:38712:11
					rf_we = 1'b1;
				if (instr[14:12] != 3'b000)
					// Trace: design.sv:38715:11
					illegal_insn = 1'b1;
				// Trace: design.sv:38718:9
				rf_ren_a_o = 1'b1;
			end
			7'h63: begin
				// Trace: design.sv:38722:9
				branch_in_dec_o = 1'b1;
				// Trace: design.sv:38724:9
				(* full_case, parallel_case *)
				case (instr[14:12])
					3'b000, 3'b001, 3'b100, 3'b101, 3'b110, 3'b111:
						// Trace: design.sv:38730:20
						illegal_insn = 1'b0;
					default:
						// Trace: design.sv:38731:20
						illegal_insn = 1'b1;
				endcase
				// Trace: design.sv:38734:9
				rf_ren_a_o = 1'b1;
				// Trace: design.sv:38735:9
				rf_ren_b_o = 1'b1;
			end
			7'h23: begin
				// Trace: design.sv:38743:9
				rf_ren_a_o = 1'b1;
				// Trace: design.sv:38744:9
				rf_ren_b_o = 1'b1;
				// Trace: design.sv:38745:9
				data_req_o = 1'b1;
				// Trace: design.sv:38746:9
				data_we_o = 1'b1;
				// Trace: design.sv:38748:9
				if (instr[14])
					// Trace: design.sv:38749:11
					illegal_insn = 1'b1;
				(* full_case, parallel_case *)
				case (instr[13:12])
					2'b00:
						// Trace: design.sv:38754:20
						data_type_o = 2'b10;
					2'b01:
						// Trace: design.sv:38755:20
						data_type_o = 2'b01;
					2'b10:
						// Trace: design.sv:38756:20
						data_type_o = 2'b00;
					default:
						// Trace: design.sv:38757:20
						illegal_insn = 1'b1;
				endcase
			end
			7'h03: begin
				// Trace: design.sv:38762:9
				rf_ren_a_o = 1'b1;
				// Trace: design.sv:38763:9
				data_req_o = 1'b1;
				// Trace: design.sv:38764:9
				data_type_o = 2'b00;
				// Trace: design.sv:38767:9
				data_sign_extension_o = ~instr[14];
				// Trace: design.sv:38770:9
				(* full_case, parallel_case *)
				case (instr[13:12])
					2'b00:
						// Trace: design.sv:38771:18
						data_type_o = 2'b10;
					2'b01:
						// Trace: design.sv:38772:18
						data_type_o = 2'b01;
					2'b10: begin
						// Trace: design.sv:38774:13
						data_type_o = 2'b00;
						// Trace: design.sv:38775:13
						if (instr[14])
							// Trace: design.sv:38776:15
							illegal_insn = 1'b1;
					end
					default:
						// Trace: design.sv:38780:13
						illegal_insn = 1'b1;
				endcase
			end
			7'h37:
				// Trace: design.sv:38790:9
				rf_we = 1'b1;
			7'h17:
				// Trace: design.sv:38794:9
				rf_we = 1'b1;
			7'h13: begin
				// Trace: design.sv:38798:9
				rf_ren_a_o = 1'b1;
				// Trace: design.sv:38799:9
				rf_we = 1'b1;
				// Trace: design.sv:38801:9
				(* full_case, parallel_case *)
				case (instr[14:12])
					3'b000, 3'b010, 3'b011, 3'b100, 3'b110, 3'b111:
						// Trace: design.sv:38807:19
						illegal_insn = 1'b0;
					3'b001:
						// Trace: design.sv:38810:13
						(* full_case, parallel_case *)
						case (instr[31:27])
							5'b00000:
								// Trace: design.sv:38811:26
								illegal_insn = (instr[26:25] == 2'b00 ? 1'b0 : 1'b1);
							5'b00100:
								// Trace: design.sv:38813:17
								illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
							5'b01001, 5'b00101, 5'b01101:
								// Trace: design.sv:38817:26
								illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
							5'b00001:
								// Trace: design.sv:38819:17
								if (instr[26] == 1'b0)
									// Trace: design.sv:38820:19
									illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
								else
									// Trace: design.sv:38822:19
									illegal_insn = 1'b1;
							5'b01100:
								// Trace: design.sv:38826:17
								(* full_case, parallel_case *)
								case (instr[26:20])
									7'b0000000, 7'b0000001, 7'b0000010, 7'b0000100, 7'b0000101:
										// Trace: design.sv:38831:32
										illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
									7'b0010000, 7'b0010001, 7'b0010010, 7'b0011000, 7'b0011001, 7'b0011010:
										// Trace: design.sv:38838:21
										illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
									default:
										// Trace: design.sv:38840:28
										illegal_insn = 1'b1;
								endcase
							default:
								// Trace: design.sv:38843:25
								illegal_insn = 1'b1;
						endcase
					3'b101:
						// Trace: design.sv:38848:13
						if (instr[26])
							// Trace: design.sv:38849:15
							illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
						else
							// Trace: design.sv:38851:15
							(* full_case, parallel_case *)
							case (instr[31:27])
								5'b00000, 5'b01000:
									// Trace: design.sv:38853:28
									illegal_insn = (instr[26:25] == 2'b00 ? 1'b0 : 1'b1);
								5'b00100:
									// Trace: design.sv:38856:19
									illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
								5'b01100, 5'b01001:
									// Trace: design.sv:38859:28
									illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
								5'b01101:
									// Trace: design.sv:38862:19
									if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
										// Trace: design.sv:38863:21
										illegal_insn = 1'b0;
									else if (RV32B == 32'sd1)
										// Trace: design.sv:38865:21
										illegal_insn = (instr[24:20] == 5'b11000 ? 1'b0 : 1'b1);
									else
										// Trace: design.sv:38867:21
										illegal_insn = 1'b1;
								5'b00101:
									// Trace: design.sv:38871:19
									if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
										// Trace: design.sv:38872:21
										illegal_insn = 1'b0;
									else if (instr[24:20] == 5'b00111)
										// Trace: design.sv:38874:21
										illegal_insn = (RV32B == 32'sd1 ? 1'b0 : 1'b1);
									else
										// Trace: design.sv:38876:21
										illegal_insn = 1'b1;
								5'b00001:
									// Trace: design.sv:38880:19
									if (instr[26] == 1'b0)
										// Trace: design.sv:38881:21
										illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
									else
										// Trace: design.sv:38883:21
										illegal_insn = 1'b1;
								default:
									// Trace: design.sv:38887:26
									illegal_insn = 1'b1;
							endcase
					default:
						// Trace: design.sv:38892:20
						illegal_insn = 1'b1;
				endcase
			end
			7'h33: begin
				// Trace: design.sv:38897:9
				rf_ren_a_o = 1'b1;
				// Trace: design.sv:38898:9
				rf_ren_b_o = 1'b1;
				// Trace: design.sv:38899:9
				rf_we = 1'b1;
				// Trace: design.sv:38900:9
				if ({instr[26], instr[13:12]} == 3'b101)
					// Trace: design.sv:38901:11
					illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
				else
					// Trace: design.sv:38903:11
					(* full_case, parallel_case *)
					case ({instr[31:25], instr[14:12]})
						10'b0000000000, 10'b0100000000, 10'b0000000010, 10'b0000000011, 10'b0000000100, 10'b0000000110, 10'b0000000111, 10'b0000000001, 10'b0000000101, 10'b0100000101:
							// Trace: design.sv:38914:36
							illegal_insn = 1'b0;
						10'b0010000010, 10'b0010000100, 10'b0010000110, 10'b0100000111, 10'b0100000110, 10'b0100000100, 10'b0110000001, 10'b0110000101, 10'b0000101100, 10'b0000101110, 10'b0000101101, 10'b0000101111, 10'b0000100100, 10'b0100100100, 10'b0000100111, 10'b0100100001, 10'b0010100001, 10'b0110100001, 10'b0100100101, 10'b0100100111:
							// Trace: design.sv:38939:36
							illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
						10'b0110100101, 10'b0010100101, 10'b0000100001, 10'b0000100101, 10'b0010100010, 10'b0010100100, 10'b0010100110, 10'b0010000001, 10'b0010000101, 10'b0000101001, 10'b0000101010, 10'b0000101011:
							// Trace: design.sv:38954:15
							illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
						10'b0100100110, 10'b0000100110:
							// Trace: design.sv:38958:36
							illegal_insn = (RV32B == 32'sd3 ? 1'b0 : 1'b1);
						10'b0000001000: begin
							// Trace: design.sv:38962:15
							multdiv_operator_o = 2'd0;
							// Trace: design.sv:38963:15
							multdiv_signed_mode_o = 2'b00;
							// Trace: design.sv:38964:15
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001001: begin
							// Trace: design.sv:38967:15
							multdiv_operator_o = 2'd1;
							// Trace: design.sv:38968:15
							multdiv_signed_mode_o = 2'b11;
							// Trace: design.sv:38969:15
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001010: begin
							// Trace: design.sv:38972:15
							multdiv_operator_o = 2'd1;
							// Trace: design.sv:38973:15
							multdiv_signed_mode_o = 2'b01;
							// Trace: design.sv:38974:15
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001011: begin
							// Trace: design.sv:38977:15
							multdiv_operator_o = 2'd1;
							// Trace: design.sv:38978:15
							multdiv_signed_mode_o = 2'b00;
							// Trace: design.sv:38979:15
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001100: begin
							// Trace: design.sv:38982:15
							multdiv_operator_o = 2'd2;
							// Trace: design.sv:38983:15
							multdiv_signed_mode_o = 2'b11;
							// Trace: design.sv:38984:15
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001101: begin
							// Trace: design.sv:38987:15
							multdiv_operator_o = 2'd2;
							// Trace: design.sv:38988:15
							multdiv_signed_mode_o = 2'b00;
							// Trace: design.sv:38989:15
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001110: begin
							// Trace: design.sv:38992:15
							multdiv_operator_o = 2'd3;
							// Trace: design.sv:38993:15
							multdiv_signed_mode_o = 2'b11;
							// Trace: design.sv:38994:15
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001111: begin
							// Trace: design.sv:38997:15
							multdiv_operator_o = 2'd3;
							// Trace: design.sv:38998:15
							multdiv_signed_mode_o = 2'b00;
							// Trace: design.sv:38999:15
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						default:
							// Trace: design.sv:39002:15
							illegal_insn = 1'b1;
					endcase
			end
			7'h0f:
				// Trace: design.sv:39013:9
				(* full_case, parallel_case *)
				case (instr[14:12])
					3'b000:
						// Trace: design.sv:39016:13
						rf_we = 1'b0;
					3'b001: begin
						// Trace: design.sv:39023:13
						jump_in_dec_o = 1'b1;
						// Trace: design.sv:39025:13
						rf_we = 1'b0;
						// Trace: design.sv:39027:13
						if (instr_first_cycle_i) begin
							// Trace: design.sv:39028:15
							jump_set_o = 1'b1;
							// Trace: design.sv:39029:15
							icache_inval_o = 1'b1;
						end
					end
					default:
						// Trace: design.sv:39033:13
						illegal_insn = 1'b1;
				endcase
			7'h73:
				// Trace: design.sv:39039:9
				if (instr[14:12] == 3'b000) begin
					// Trace: design.sv:39041:11
					(* full_case, parallel_case *)
					case (instr[31:20])
						12'h000:
							// Trace: design.sv:39044:15
							ecall_insn_o = 1'b1;
						12'h001:
							// Trace: design.sv:39048:15
							ebrk_insn_o = 1'b1;
						12'h302:
							// Trace: design.sv:39051:15
							mret_insn_o = 1'b1;
						12'h7b2:
							// Trace: design.sv:39054:15
							dret_insn_o = 1'b1;
						12'h105:
							// Trace: design.sv:39057:15
							wfi_insn_o = 1'b1;
						default:
							// Trace: design.sv:39060:15
							illegal_insn = 1'b1;
					endcase
					if ((instr_rs1 != 5'b00000) || (instr_rd != 5'b00000))
						// Trace: design.sv:39065:13
						illegal_insn = 1'b1;
				end
				else begin
					// Trace: design.sv:39069:11
					csr_access_o = 1'b1;
					// Trace: design.sv:39070:11
					rf_wdata_sel_o = 1'd1;
					// Trace: design.sv:39071:11
					rf_we = 1'b1;
					// Trace: design.sv:39073:11
					if (~instr[14])
						// Trace: design.sv:39074:13
						rf_ren_a_o = 1'b1;
					(* full_case, parallel_case *)
					case (instr[13:12])
						2'b01:
							// Trace: design.sv:39078:22
							csr_op = 2'd1;
						2'b10:
							// Trace: design.sv:39079:22
							csr_op = 2'd2;
						2'b11:
							// Trace: design.sv:39080:22
							csr_op = 2'd3;
						default:
							// Trace: design.sv:39081:22
							csr_illegal = 1'b1;
					endcase
					// Trace: design.sv:39084:11
					illegal_insn = csr_illegal;
				end
			default:
				// Trace: design.sv:39089:9
				illegal_insn = 1'b1;
		endcase
		if (illegal_c_insn_i)
			// Trace: design.sv:39095:7
			illegal_insn = 1'b1;
		if (illegal_insn) begin
			// Trace: design.sv:39104:7
			rf_we = 1'b0;
			// Trace: design.sv:39105:7
			data_req_o = 1'b0;
			// Trace: design.sv:39106:7
			data_we_o = 1'b0;
			// Trace: design.sv:39107:7
			jump_in_dec_o = 1'b0;
			// Trace: design.sv:39108:7
			jump_set_o = 1'b0;
			// Trace: design.sv:39109:7
			branch_in_dec_o = 1'b0;
			// Trace: design.sv:39110:7
			csr_access_o = 1'b0;
		end
	end
	// Trace: design.sv:39118:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:39119:5
		alu_operator_o = 7'd44;
		// Trace: design.sv:39120:5
		alu_op_a_mux_sel_o = 2'd3;
		// Trace: design.sv:39121:5
		alu_op_b_mux_sel_o = 1'd1;
		// Trace: design.sv:39123:5
		imm_a_mux_sel_o = 1'd1;
		// Trace: design.sv:39124:5
		imm_b_mux_sel_o = 3'd0;
		// Trace: design.sv:39126:5
		bt_a_mux_sel_o = 2'd2;
		// Trace: design.sv:39127:5
		bt_b_mux_sel_o = 3'd0;
		// Trace: design.sv:39130:5
		opcode_alu = instr_alu[6:0];
		// Trace: design.sv:39132:5
		use_rs3_d = 1'b0;
		// Trace: design.sv:39133:5
		alu_multicycle_o = 1'b0;
		// Trace: design.sv:39134:5
		mult_sel_o = 1'b0;
		// Trace: design.sv:39135:5
		div_sel_o = 1'b0;
		// Trace: design.sv:39137:5
		(* full_case, parallel_case *)
		case (opcode_alu)
			7'h6f: begin
				// Trace: design.sv:39144:9
				if (BranchTargetALU) begin
					// Trace: design.sv:39145:11
					bt_a_mux_sel_o = 2'd2;
					// Trace: design.sv:39146:11
					bt_b_mux_sel_o = 3'd4;
				end
				if (instr_first_cycle_i && !BranchTargetALU) begin
					// Trace: design.sv:39152:11
					alu_op_a_mux_sel_o = 2'd2;
					// Trace: design.sv:39153:11
					alu_op_b_mux_sel_o = 1'd1;
					// Trace: design.sv:39154:11
					imm_b_mux_sel_o = 3'd4;
					// Trace: design.sv:39155:11
					alu_operator_o = 7'd0;
				end
				else begin
					// Trace: design.sv:39158:11
					alu_op_a_mux_sel_o = 2'd2;
					// Trace: design.sv:39159:11
					alu_op_b_mux_sel_o = 1'd1;
					// Trace: design.sv:39160:11
					imm_b_mux_sel_o = 3'd5;
					// Trace: design.sv:39161:11
					alu_operator_o = 7'd0;
				end
			end
			7'h67: begin
				// Trace: design.sv:39166:9
				if (BranchTargetALU) begin
					// Trace: design.sv:39167:11
					bt_a_mux_sel_o = 2'd0;
					// Trace: design.sv:39168:11
					bt_b_mux_sel_o = 3'd0;
				end
				if (instr_first_cycle_i && !BranchTargetALU) begin
					// Trace: design.sv:39174:11
					alu_op_a_mux_sel_o = 2'd0;
					// Trace: design.sv:39175:11
					alu_op_b_mux_sel_o = 1'd1;
					// Trace: design.sv:39176:11
					imm_b_mux_sel_o = 3'd0;
					// Trace: design.sv:39177:11
					alu_operator_o = 7'd0;
				end
				else begin
					// Trace: design.sv:39180:11
					alu_op_a_mux_sel_o = 2'd2;
					// Trace: design.sv:39181:11
					alu_op_b_mux_sel_o = 1'd1;
					// Trace: design.sv:39182:11
					imm_b_mux_sel_o = 3'd5;
					// Trace: design.sv:39183:11
					alu_operator_o = 7'd0;
				end
			end
			7'h63: begin
				// Trace: design.sv:39189:9
				(* full_case, parallel_case *)
				case (instr_alu[14:12])
					3'b000:
						// Trace: design.sv:39190:20
						alu_operator_o = 7'd29;
					3'b001:
						// Trace: design.sv:39191:20
						alu_operator_o = 7'd30;
					3'b100:
						// Trace: design.sv:39192:20
						alu_operator_o = 7'd25;
					3'b101:
						// Trace: design.sv:39193:20
						alu_operator_o = 7'd27;
					3'b110:
						// Trace: design.sv:39194:20
						alu_operator_o = 7'd26;
					3'b111:
						// Trace: design.sv:39195:20
						alu_operator_o = 7'd28;
					default:
						;
				endcase
				if (BranchTargetALU) begin
					// Trace: design.sv:39200:11
					bt_a_mux_sel_o = 2'd2;
					// Trace: design.sv:39202:11
					bt_b_mux_sel_o = (branch_taken_i ? 3'd2 : 3'd5);
				end
				if (instr_first_cycle_i) begin
					// Trace: design.sv:39209:11
					alu_op_a_mux_sel_o = 2'd0;
					// Trace: design.sv:39210:11
					alu_op_b_mux_sel_o = 1'd0;
				end
				else if (!BranchTargetALU) begin
					// Trace: design.sv:39213:11
					alu_op_a_mux_sel_o = 2'd2;
					// Trace: design.sv:39214:11
					alu_op_b_mux_sel_o = 1'd1;
					// Trace: design.sv:39216:11
					imm_b_mux_sel_o = (branch_taken_i ? 3'd2 : 3'd5);
					// Trace: design.sv:39217:11
					alu_operator_o = 7'd0;
				end
			end
			7'h23: begin
				// Trace: design.sv:39226:9
				alu_op_a_mux_sel_o = 2'd0;
				// Trace: design.sv:39227:9
				alu_op_b_mux_sel_o = 1'd0;
				// Trace: design.sv:39228:9
				alu_operator_o = 7'd0;
				// Trace: design.sv:39230:9
				if (!instr_alu[14]) begin
					// Trace: design.sv:39232:11
					imm_b_mux_sel_o = 3'd1;
					// Trace: design.sv:39233:11
					alu_op_b_mux_sel_o = 1'd1;
				end
			end
			7'h03: begin
				// Trace: design.sv:39238:9
				alu_op_a_mux_sel_o = 2'd0;
				// Trace: design.sv:39241:9
				alu_operator_o = 7'd0;
				// Trace: design.sv:39242:9
				alu_op_b_mux_sel_o = 1'd1;
				// Trace: design.sv:39243:9
				imm_b_mux_sel_o = 3'd0;
			end
			7'h37: begin
				// Trace: design.sv:39251:9
				alu_op_a_mux_sel_o = 2'd3;
				// Trace: design.sv:39252:9
				alu_op_b_mux_sel_o = 1'd1;
				// Trace: design.sv:39253:9
				imm_a_mux_sel_o = 1'd1;
				// Trace: design.sv:39254:9
				imm_b_mux_sel_o = 3'd3;
				// Trace: design.sv:39255:9
				alu_operator_o = 7'd0;
			end
			7'h17: begin
				// Trace: design.sv:39259:9
				alu_op_a_mux_sel_o = 2'd2;
				// Trace: design.sv:39260:9
				alu_op_b_mux_sel_o = 1'd1;
				// Trace: design.sv:39261:9
				imm_b_mux_sel_o = 3'd3;
				// Trace: design.sv:39262:9
				alu_operator_o = 7'd0;
			end
			7'h13: begin
				// Trace: design.sv:39266:9
				alu_op_a_mux_sel_o = 2'd0;
				// Trace: design.sv:39267:9
				alu_op_b_mux_sel_o = 1'd1;
				// Trace: design.sv:39268:9
				imm_b_mux_sel_o = 3'd0;
				// Trace: design.sv:39270:9
				(* full_case, parallel_case *)
				case (instr_alu[14:12])
					3'b000:
						// Trace: design.sv:39271:19
						alu_operator_o = 7'd0;
					3'b010:
						// Trace: design.sv:39272:19
						alu_operator_o = 7'd43;
					3'b011:
						// Trace: design.sv:39273:19
						alu_operator_o = 7'd44;
					3'b100:
						// Trace: design.sv:39274:19
						alu_operator_o = 7'd2;
					3'b110:
						// Trace: design.sv:39275:19
						alu_operator_o = 7'd3;
					3'b111:
						// Trace: design.sv:39276:19
						alu_operator_o = 7'd4;
					3'b001:
						// Trace: design.sv:39279:13
						if (RV32B != 32'sd0)
							// Trace: design.sv:39280:15
							(* full_case, parallel_case *)
							case (instr_alu[31:27])
								5'b00000:
									// Trace: design.sv:39281:28
									alu_operator_o = 7'd10;
								5'b00100:
									// Trace: design.sv:39284:19
									if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
										// Trace: design.sv:39284:71
										alu_operator_o = 7'd12;
								5'b01001:
									// Trace: design.sv:39286:28
									alu_operator_o = 7'd50;
								5'b00101:
									// Trace: design.sv:39287:28
									alu_operator_o = 7'd49;
								5'b01101:
									// Trace: design.sv:39288:28
									alu_operator_o = 7'd51;
								5'b00001:
									if (instr_alu[26] == 0)
										// Trace: design.sv:39290:52
										alu_operator_o = 7'd17;
								5'b01100:
									// Trace: design.sv:39292:19
									(* full_case, parallel_case *)
									case (instr_alu[26:20])
										7'b0000000:
											// Trace: design.sv:39293:34
											alu_operator_o = 7'd40;
										7'b0000001:
											// Trace: design.sv:39294:34
											alu_operator_o = 7'd41;
										7'b0000010:
											// Trace: design.sv:39295:34
											alu_operator_o = 7'd42;
										7'b0000100:
											// Trace: design.sv:39296:34
											alu_operator_o = 7'd38;
										7'b0000101:
											// Trace: design.sv:39297:34
											alu_operator_o = 7'd39;
										7'b0010000:
											// Trace: design.sv:39299:23
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												// Trace: design.sv:39300:25
												alu_operator_o = 7'd59;
												// Trace: design.sv:39301:25
												alu_multicycle_o = 1'b1;
											end
										7'b0010001:
											// Trace: design.sv:39305:23
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												// Trace: design.sv:39306:25
												alu_operator_o = 7'd61;
												// Trace: design.sv:39307:25
												alu_multicycle_o = 1'b1;
											end
										7'b0010010:
											// Trace: design.sv:39311:23
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												// Trace: design.sv:39312:25
												alu_operator_o = 7'd63;
												// Trace: design.sv:39313:25
												alu_multicycle_o = 1'b1;
											end
										7'b0011000:
											// Trace: design.sv:39317:23
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												// Trace: design.sv:39318:25
												alu_operator_o = 7'd60;
												// Trace: design.sv:39319:25
												alu_multicycle_o = 1'b1;
											end
										7'b0011001:
											// Trace: design.sv:39323:23
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												// Trace: design.sv:39324:25
												alu_operator_o = 7'd62;
												// Trace: design.sv:39325:25
												alu_multicycle_o = 1'b1;
											end
										7'b0011010:
											// Trace: design.sv:39329:23
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												// Trace: design.sv:39330:25
												alu_operator_o = 7'd64;
												// Trace: design.sv:39331:25
												alu_multicycle_o = 1'b1;
											end
										default:
											;
									endcase
								default:
									;
							endcase
						else
							// Trace: design.sv:39341:15
							alu_operator_o = 7'd10;
					3'b101:
						// Trace: design.sv:39346:13
						if (RV32B != 32'sd0) begin
							begin
								// Trace: design.sv:39347:15
								if (instr_alu[26] == 1'b1) begin
									// Trace: design.sv:39348:17
									alu_operator_o = 7'd48;
									// Trace: design.sv:39349:17
									alu_multicycle_o = 1'b1;
									// Trace: design.sv:39350:17
									if (instr_first_cycle_i)
										// Trace: design.sv:39351:19
										use_rs3_d = 1'b1;
									else
										// Trace: design.sv:39353:19
										use_rs3_d = 1'b0;
								end
								else
									// Trace: design.sv:39356:17
									(* full_case, parallel_case *)
									case (instr_alu[31:27])
										5'b00000:
											// Trace: design.sv:39357:30
											alu_operator_o = 7'd9;
										5'b01000:
											// Trace: design.sv:39358:30
											alu_operator_o = 7'd8;
										5'b00100:
											// Trace: design.sv:39361:21
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
												// Trace: design.sv:39361:73
												alu_operator_o = 7'd11;
										5'b01001:
											// Trace: design.sv:39363:30
											alu_operator_o = 7'd52;
										5'b01100: begin
											// Trace: design.sv:39365:21
											alu_operator_o = 7'd13;
											// Trace: design.sv:39366:21
											alu_multicycle_o = 1'b1;
										end
										5'b01101:
											// Trace: design.sv:39368:30
											alu_operator_o = 7'd15;
										5'b00101:
											// Trace: design.sv:39369:30
											alu_operator_o = 7'd16;
										5'b00001:
											// Trace: design.sv:39372:21
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												begin
													// Trace: design.sv:39373:23
													if (instr_alu[26] == 1'b0)
														// Trace: design.sv:39373:50
														alu_operator_o = 7'd18;
												end
											end
										default:
											;
									endcase
							end
						end
						else
							// Trace: design.sv:39381:15
							if (instr_alu[31:27] == 5'b00000)
								// Trace: design.sv:39382:17
								alu_operator_o = 7'd9;
							else if (instr_alu[31:27] == 5'b01000)
								// Trace: design.sv:39384:17
								alu_operator_o = 7'd8;
					default:
						;
				endcase
			end
			7'h33: begin
				// Trace: design.sv:39394:9
				alu_op_a_mux_sel_o = 2'd0;
				// Trace: design.sv:39395:9
				alu_op_b_mux_sel_o = 1'd0;
				// Trace: design.sv:39397:9
				if (instr_alu[26]) begin
					begin
						// Trace: design.sv:39398:11
						if (RV32B != 32'sd0)
							// Trace: design.sv:39399:13
							(* full_case, parallel_case *)
							case ({instr_alu[26:25], instr_alu[14:12]})
								5'b11001: begin
									// Trace: design.sv:39401:17
									alu_operator_o = 7'd46;
									// Trace: design.sv:39402:17
									alu_multicycle_o = 1'b1;
									// Trace: design.sv:39403:17
									if (instr_first_cycle_i)
										// Trace: design.sv:39404:19
										use_rs3_d = 1'b1;
									else
										// Trace: design.sv:39406:19
										use_rs3_d = 1'b0;
								end
								5'b11101: begin
									// Trace: design.sv:39410:17
									alu_operator_o = 7'd45;
									// Trace: design.sv:39411:17
									alu_multicycle_o = 1'b1;
									// Trace: design.sv:39412:17
									if (instr_first_cycle_i)
										// Trace: design.sv:39413:19
										use_rs3_d = 1'b1;
									else
										// Trace: design.sv:39415:19
										use_rs3_d = 1'b0;
								end
								5'b10001: begin
									// Trace: design.sv:39419:17
									alu_operator_o = 7'd47;
									// Trace: design.sv:39420:17
									alu_multicycle_o = 1'b1;
									// Trace: design.sv:39421:17
									if (instr_first_cycle_i)
										// Trace: design.sv:39422:19
										use_rs3_d = 1'b1;
									else
										// Trace: design.sv:39424:19
										use_rs3_d = 1'b0;
								end
								5'b10101: begin
									// Trace: design.sv:39428:17
									alu_operator_o = 7'd48;
									// Trace: design.sv:39429:17
									alu_multicycle_o = 1'b1;
									// Trace: design.sv:39430:17
									if (instr_first_cycle_i)
										// Trace: design.sv:39431:19
										use_rs3_d = 1'b1;
									else
										// Trace: design.sv:39433:19
										use_rs3_d = 1'b0;
								end
								default:
									;
							endcase
					end
				end
				else
					// Trace: design.sv:39440:11
					(* full_case, parallel_case *)
					case ({instr_alu[31:25], instr_alu[14:12]})
						10'b0000000000:
							// Trace: design.sv:39442:36
							alu_operator_o = 7'd0;
						10'b0100000000:
							// Trace: design.sv:39443:36
							alu_operator_o = 7'd1;
						10'b0000000010:
							// Trace: design.sv:39444:36
							alu_operator_o = 7'd43;
						10'b0000000011:
							// Trace: design.sv:39445:36
							alu_operator_o = 7'd44;
						10'b0000000100:
							// Trace: design.sv:39446:36
							alu_operator_o = 7'd2;
						10'b0000000110:
							// Trace: design.sv:39447:36
							alu_operator_o = 7'd3;
						10'b0000000111:
							// Trace: design.sv:39448:36
							alu_operator_o = 7'd4;
						10'b0000000001:
							// Trace: design.sv:39449:36
							alu_operator_o = 7'd10;
						10'b0000000101:
							// Trace: design.sv:39450:36
							alu_operator_o = 7'd9;
						10'b0100000101:
							// Trace: design.sv:39451:36
							alu_operator_o = 7'd8;
						10'b0110000001:
							// Trace: design.sv:39455:15
							if (RV32B != 32'sd0) begin
								// Trace: design.sv:39456:17
								alu_operator_o = 7'd14;
								// Trace: design.sv:39457:17
								alu_multicycle_o = 1'b1;
							end
						10'b0110000101:
							// Trace: design.sv:39461:15
							if (RV32B != 32'sd0) begin
								// Trace: design.sv:39462:17
								alu_operator_o = 7'd13;
								// Trace: design.sv:39463:17
								alu_multicycle_o = 1'b1;
							end
						10'b0000101100:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39467:60
								alu_operator_o = 7'd31;
						10'b0000101110:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39468:60
								alu_operator_o = 7'd33;
						10'b0000101101:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39469:60
								alu_operator_o = 7'd32;
						10'b0000101111:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39470:60
								alu_operator_o = 7'd34;
						10'b0000100100:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39472:60
								alu_operator_o = 7'd35;
						10'b0100100100:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39473:60
								alu_operator_o = 7'd36;
						10'b0000100111:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39474:60
								alu_operator_o = 7'd37;
						10'b0100000100:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39476:60
								alu_operator_o = 7'd5;
						10'b0100000110:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39477:60
								alu_operator_o = 7'd6;
						10'b0100000111:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39478:60
								alu_operator_o = 7'd7;
						10'b0010000010:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39481:60
								alu_operator_o = 7'd22;
						10'b0010000100:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39482:60
								alu_operator_o = 7'd23;
						10'b0010000110:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39483:60
								alu_operator_o = 7'd24;
						10'b0100100001:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39486:60
								alu_operator_o = 7'd50;
						10'b0010100001:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39487:60
								alu_operator_o = 7'd49;
						10'b0110100001:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39488:60
								alu_operator_o = 7'd51;
						10'b0100100101:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39489:60
								alu_operator_o = 7'd52;
						10'b0100100111:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39492:60
								alu_operator_o = 7'd55;
						10'b0110100101:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39495:60
								alu_operator_o = 7'd15;
						10'b0010100101:
							if (RV32B != 32'sd0)
								// Trace: design.sv:39496:60
								alu_operator_o = 7'd16;
						10'b0000100001:
							// Trace: design.sv:39498:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39498:67
								alu_operator_o = 7'd17;
						10'b0000100101:
							// Trace: design.sv:39501:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39501:67
								alu_operator_o = 7'd18;
						10'b0010100010:
							// Trace: design.sv:39504:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39504:67
								alu_operator_o = 7'd19;
						10'b0010100100:
							// Trace: design.sv:39507:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39507:67
								alu_operator_o = 7'd20;
						10'b0010100110:
							// Trace: design.sv:39510:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39510:67
								alu_operator_o = 7'd21;
						10'b0010000001:
							// Trace: design.sv:39513:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39513:67
								alu_operator_o = 7'd12;
						10'b0010000101:
							// Trace: design.sv:39516:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39516:67
								alu_operator_o = 7'd11;
						10'b0000101001:
							// Trace: design.sv:39521:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39521:67
								alu_operator_o = 7'd56;
						10'b0000101010:
							// Trace: design.sv:39524:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39524:67
								alu_operator_o = 7'd57;
						10'b0000101011:
							// Trace: design.sv:39527:15
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								// Trace: design.sv:39527:67
								alu_operator_o = 7'd58;
						10'b0100100110:
							// Trace: design.sv:39532:15
							if (RV32B == 32'sd3) begin
								// Trace: design.sv:39533:17
								alu_operator_o = 7'd54;
								// Trace: design.sv:39534:17
								alu_multicycle_o = 1'b1;
							end
						10'b0000100110:
							// Trace: design.sv:39538:15
							if (RV32B == 32'sd3) begin
								// Trace: design.sv:39539:17
								alu_operator_o = 7'd53;
								// Trace: design.sv:39540:17
								alu_multicycle_o = 1'b1;
							end
						10'b0000001000: begin
							// Trace: design.sv:39546:15
							alu_operator_o = 7'd0;
							// Trace: design.sv:39547:15
							mult_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001001: begin
							// Trace: design.sv:39550:15
							alu_operator_o = 7'd0;
							// Trace: design.sv:39551:15
							mult_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001010: begin
							// Trace: design.sv:39554:15
							alu_operator_o = 7'd0;
							// Trace: design.sv:39555:15
							mult_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001011: begin
							// Trace: design.sv:39558:15
							alu_operator_o = 7'd0;
							// Trace: design.sv:39559:15
							mult_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001100: begin
							// Trace: design.sv:39562:15
							alu_operator_o = 7'd0;
							// Trace: design.sv:39563:15
							div_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001101: begin
							// Trace: design.sv:39566:15
							alu_operator_o = 7'd0;
							// Trace: design.sv:39567:15
							div_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001110: begin
							// Trace: design.sv:39570:15
							alu_operator_o = 7'd0;
							// Trace: design.sv:39571:15
							div_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001111: begin
							// Trace: design.sv:39574:15
							alu_operator_o = 7'd0;
							// Trace: design.sv:39575:15
							div_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						default:
							;
					endcase
			end
			7'h0f:
				// Trace: design.sv:39588:9
				(* full_case, parallel_case *)
				case (instr_alu[14:12])
					3'b000: begin
						// Trace: design.sv:39591:13
						alu_operator_o = 7'd0;
						// Trace: design.sv:39592:13
						alu_op_a_mux_sel_o = 2'd0;
						// Trace: design.sv:39593:13
						alu_op_b_mux_sel_o = 1'd1;
					end
					3'b001:
						// Trace: design.sv:39597:13
						if (BranchTargetALU) begin
							// Trace: design.sv:39598:15
							bt_a_mux_sel_o = 2'd2;
							// Trace: design.sv:39599:15
							bt_b_mux_sel_o = 3'd5;
						end
						else begin
							// Trace: design.sv:39601:15
							alu_op_a_mux_sel_o = 2'd2;
							// Trace: design.sv:39602:15
							alu_op_b_mux_sel_o = 1'd1;
							// Trace: design.sv:39603:15
							imm_b_mux_sel_o = 3'd5;
							// Trace: design.sv:39604:15
							alu_operator_o = 7'd0;
						end
					default:
						;
				endcase
			7'h73:
				// Trace: design.sv:39612:9
				if (instr_alu[14:12] == 3'b000) begin
					// Trace: design.sv:39614:11
					alu_op_a_mux_sel_o = 2'd0;
					// Trace: design.sv:39615:11
					alu_op_b_mux_sel_o = 1'd1;
				end
				else begin
					// Trace: design.sv:39618:11
					alu_op_b_mux_sel_o = 1'd1;
					// Trace: design.sv:39619:11
					imm_a_mux_sel_o = 1'd0;
					// Trace: design.sv:39620:11
					imm_b_mux_sel_o = 3'd0;
					// Trace: design.sv:39622:11
					if (instr_alu[14])
						// Trace: design.sv:39624:13
						alu_op_a_mux_sel_o = 2'd3;
					else
						// Trace: design.sv:39626:13
						alu_op_a_mux_sel_o = 2'd0;
				end
			default:
				;
		endcase
	end
	// Trace: design.sv:39636:3
	assign mult_en_o = (illegal_insn ? 1'b0 : mult_sel_o);
	// Trace: design.sv:39637:3
	assign div_en_o = (illegal_insn ? 1'b0 : div_sel_o);
	// Trace: design.sv:39641:3
	assign illegal_insn_o = illegal_insn | illegal_reg_rv32e;
	// Trace: design.sv:39644:3
	assign rf_we_o = rf_we & ~illegal_reg_rv32e;
	// Trace: design.sv:39647:3
	assign unused_instr_alu = {instr_alu[19:15], instr_alu[11:7]};
	initial _sv2v_0 = 0;
endmodule
module ibex_ex_block (
	clk_i,
	rst_ni,
	alu_operator_i,
	alu_operand_a_i,
	alu_operand_b_i,
	alu_instr_first_cycle_i,
	bt_a_operand_i,
	bt_b_operand_i,
	multdiv_operator_i,
	mult_en_i,
	div_en_i,
	mult_sel_i,
	div_sel_i,
	multdiv_signed_mode_i,
	multdiv_operand_a_i,
	multdiv_operand_b_i,
	multdiv_ready_id_i,
	data_ind_timing_i,
	imd_val_we_o,
	imd_val_d_o,
	imd_val_q_i,
	alu_adder_result_ex_o,
	result_ex_o,
	branch_target_o,
	branch_decision_o,
	ex_valid_o
);
	// Trace: design.sv:39668:13
	// removed localparam type ibex_pkg_rv32m_e
	parameter integer RV32M = 32'sd2;
	// Trace: design.sv:39669:13
	// removed localparam type ibex_pkg_rv32b_e
	parameter integer RV32B = 32'sd0;
	// Trace: design.sv:39670:13
	parameter [0:0] BranchTargetALU = 0;
	// Trace: design.sv:39672:3
	input wire clk_i;
	// Trace: design.sv:39673:3
	input wire rst_ni;
	// Trace: design.sv:39676:3
	// removed localparam type ibex_pkg_alu_op_e
	input wire [6:0] alu_operator_i;
	// Trace: design.sv:39677:3
	input wire [31:0] alu_operand_a_i;
	// Trace: design.sv:39678:3
	input wire [31:0] alu_operand_b_i;
	// Trace: design.sv:39679:3
	input wire alu_instr_first_cycle_i;
	// Trace: design.sv:39683:3
	input wire [31:0] bt_a_operand_i;
	// Trace: design.sv:39684:3
	input wire [31:0] bt_b_operand_i;
	// Trace: design.sv:39687:3
	// removed localparam type ibex_pkg_md_op_e
	input wire [1:0] multdiv_operator_i;
	// Trace: design.sv:39688:3
	input wire mult_en_i;
	// Trace: design.sv:39689:3
	input wire div_en_i;
	// Trace: design.sv:39690:3
	input wire mult_sel_i;
	// Trace: design.sv:39691:3
	input wire div_sel_i;
	// Trace: design.sv:39692:3
	input wire [1:0] multdiv_signed_mode_i;
	// Trace: design.sv:39693:3
	input wire [31:0] multdiv_operand_a_i;
	// Trace: design.sv:39694:3
	input wire [31:0] multdiv_operand_b_i;
	// Trace: design.sv:39695:3
	input wire multdiv_ready_id_i;
	// Trace: design.sv:39696:3
	input wire data_ind_timing_i;
	// Trace: design.sv:39699:3
	output wire [1:0] imd_val_we_o;
	// Trace: design.sv:39700:3
	output wire [67:0] imd_val_d_o;
	// Trace: design.sv:39701:3
	input wire [67:0] imd_val_q_i;
	// Trace: design.sv:39704:3
	output wire [31:0] alu_adder_result_ex_o;
	// Trace: design.sv:39705:3
	output wire [31:0] result_ex_o;
	// Trace: design.sv:39706:3
	output wire [31:0] branch_target_o;
	// Trace: design.sv:39707:3
	output wire branch_decision_o;
	// Trace: design.sv:39709:3
	output wire ex_valid_o;
	// Trace: design.sv:39712:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:39714:3
	wire [31:0] alu_result;
	wire [31:0] multdiv_result;
	// Trace: design.sv:39716:3
	wire [32:0] multdiv_alu_operand_b;
	wire [32:0] multdiv_alu_operand_a;
	// Trace: design.sv:39717:3
	wire [33:0] alu_adder_result_ext;
	// Trace: design.sv:39718:3
	wire alu_cmp_result;
	wire alu_is_equal_result;
	// Trace: design.sv:39719:3
	wire multdiv_valid;
	// Trace: design.sv:39720:3
	wire multdiv_sel;
	// Trace: design.sv:39721:3
	wire [63:0] alu_imd_val_q;
	// Trace: design.sv:39722:3
	wire [63:0] alu_imd_val_d;
	// Trace: design.sv:39723:3
	wire [1:0] alu_imd_val_we;
	// Trace: design.sv:39724:3
	wire [67:0] multdiv_imd_val_d;
	// Trace: design.sv:39725:3
	wire [1:0] multdiv_imd_val_we;
	// Trace: design.sv:39732:3
	generate
		if (RV32M != 32'sd0) begin : gen_multdiv_m
			// Trace: design.sv:39733:5
			assign multdiv_sel = mult_sel_i | div_sel_i;
		end
		else begin : gen_multdiv_no_m
			// Trace: design.sv:39735:5
			assign multdiv_sel = 1'b0;
		end
	endgenerate
	// Trace: design.sv:39739:3
	assign imd_val_d_o[34+:34] = (multdiv_sel ? multdiv_imd_val_d[34+:34] : {2'b00, alu_imd_val_d[32+:32]});
	// Trace: design.sv:39740:3
	assign imd_val_d_o[0+:34] = (multdiv_sel ? multdiv_imd_val_d[0+:34] : {2'b00, alu_imd_val_d[0+:32]});
	// Trace: design.sv:39741:3
	assign imd_val_we_o = (multdiv_sel ? multdiv_imd_val_we : alu_imd_val_we);
	// Trace: design.sv:39743:3
	assign alu_imd_val_q = {imd_val_q_i[65-:32], imd_val_q_i[31-:32]};
	// Trace: design.sv:39745:3
	assign result_ex_o = (multdiv_sel ? multdiv_result : alu_result);
	// Trace: design.sv:39748:3
	assign branch_decision_o = alu_cmp_result;
	// Trace: design.sv:39750:3
	generate
		if (BranchTargetALU) begin : g_branch_target_alu
			// Trace: design.sv:39751:5
			wire [32:0] bt_alu_result;
			// Trace: design.sv:39752:5
			wire unused_bt_carry;
			// Trace: design.sv:39754:5
			assign bt_alu_result = bt_a_operand_i + bt_b_operand_i;
			// Trace: design.sv:39756:5
			assign unused_bt_carry = bt_alu_result[32];
			// Trace: design.sv:39757:5
			assign branch_target_o = bt_alu_result[31:0];
		end
		else begin : g_no_branch_target_alu
			// Trace: design.sv:39760:5
			wire [31:0] unused_bt_a_operand;
			wire [31:0] unused_bt_b_operand;
			// Trace: design.sv:39762:5
			assign unused_bt_a_operand = bt_a_operand_i;
			// Trace: design.sv:39763:5
			assign unused_bt_b_operand = bt_b_operand_i;
			// Trace: design.sv:39765:5
			assign branch_target_o = alu_adder_result_ex_o;
		end
	endgenerate
	// Trace: design.sv:39772:3
	ibex_alu #(.RV32B(RV32B)) alu_i(
		.operator_i(alu_operator_i),
		.operand_a_i(alu_operand_a_i),
		.operand_b_i(alu_operand_b_i),
		.instr_first_cycle_i(alu_instr_first_cycle_i),
		.imd_val_q_i(alu_imd_val_q),
		.imd_val_we_o(alu_imd_val_we),
		.imd_val_d_o(alu_imd_val_d),
		.multdiv_operand_a_i(multdiv_alu_operand_a),
		.multdiv_operand_b_i(multdiv_alu_operand_b),
		.multdiv_sel_i(multdiv_sel),
		.adder_result_o(alu_adder_result_ex_o),
		.adder_result_ext_o(alu_adder_result_ext),
		.result_o(alu_result),
		.comparison_result_o(alu_cmp_result),
		.is_equal_result_o(alu_is_equal_result)
	);
	// Trace: design.sv:39796:3
	generate
		if (RV32M == 32'sd1) begin : gen_multdiv_slow
			// Trace: design.sv:39797:5
			ibex_multdiv_slow multdiv_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.mult_en_i(mult_en_i),
				.div_en_i(div_en_i),
				.mult_sel_i(mult_sel_i),
				.div_sel_i(div_sel_i),
				.operator_i(multdiv_operator_i),
				.signed_mode_i(multdiv_signed_mode_i),
				.op_a_i(multdiv_operand_a_i),
				.op_b_i(multdiv_operand_b_i),
				.alu_adder_ext_i(alu_adder_result_ext),
				.alu_adder_i(alu_adder_result_ex_o),
				.equal_to_zero_i(alu_is_equal_result),
				.data_ind_timing_i(data_ind_timing_i),
				.valid_o(multdiv_valid),
				.alu_operand_a_o(multdiv_alu_operand_a),
				.alu_operand_b_o(multdiv_alu_operand_b),
				.imd_val_q_i(imd_val_q_i),
				.imd_val_d_o(multdiv_imd_val_d),
				.imd_val_we_o(multdiv_imd_val_we),
				.multdiv_ready_id_i(multdiv_ready_id_i),
				.multdiv_result_o(multdiv_result)
			);
		end
		else if ((RV32M == 32'sd2) || (RV32M == 32'sd3)) begin : gen_multdiv_fast
			// Trace: design.sv:39822:5
			ibex_multdiv_fast #(.RV32M(RV32M)) multdiv_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.mult_en_i(mult_en_i),
				.div_en_i(div_en_i),
				.mult_sel_i(mult_sel_i),
				.div_sel_i(div_sel_i),
				.operator_i(multdiv_operator_i),
				.signed_mode_i(multdiv_signed_mode_i),
				.op_a_i(multdiv_operand_a_i),
				.op_b_i(multdiv_operand_b_i),
				.alu_operand_a_o(multdiv_alu_operand_a),
				.alu_operand_b_o(multdiv_alu_operand_b),
				.alu_adder_ext_i(alu_adder_result_ext),
				.alu_adder_i(alu_adder_result_ex_o),
				.equal_to_zero_i(alu_is_equal_result),
				.data_ind_timing_i(data_ind_timing_i),
				.imd_val_q_i(imd_val_q_i),
				.imd_val_d_o(multdiv_imd_val_d),
				.imd_val_we_o(multdiv_imd_val_we),
				.multdiv_ready_id_i(multdiv_ready_id_i),
				.valid_o(multdiv_valid),
				.multdiv_result_o(multdiv_result)
			);
		end
	endgenerate
	// Trace: design.sv:39853:3
	assign ex_valid_o = (multdiv_sel ? multdiv_valid : ~(|alu_imd_val_we));
endmodule
module ibex_fetch_fifo (
	clk_i,
	rst_ni,
	clear_i,
	busy_o,
	in_valid_i,
	in_addr_i,
	in_rdata_i,
	in_err_i,
	out_valid_o,
	out_ready_i,
	out_addr_o,
	out_rdata_o,
	out_err_o,
	out_err_plus2_o
);
	reg _sv2v_0;
	// Trace: design.sv:39871:13
	parameter [31:0] NUM_REQS = 2;
	// Trace: design.sv:39872:13
	parameter [0:0] ResetAll = 1'b0;
	// Trace: design.sv:39874:3
	input wire clk_i;
	// Trace: design.sv:39875:3
	input wire rst_ni;
	// Trace: design.sv:39878:3
	input wire clear_i;
	// Trace: design.sv:39879:3
	output wire [NUM_REQS - 1:0] busy_o;
	// Trace: design.sv:39882:3
	input wire in_valid_i;
	// Trace: design.sv:39883:3
	input wire [31:0] in_addr_i;
	// Trace: design.sv:39884:3
	input wire [31:0] in_rdata_i;
	// Trace: design.sv:39885:3
	input wire in_err_i;
	// Trace: design.sv:39888:3
	output reg out_valid_o;
	// Trace: design.sv:39889:3
	input wire out_ready_i;
	// Trace: design.sv:39890:3
	output wire [31:0] out_addr_o;
	// Trace: design.sv:39891:3
	output reg [31:0] out_rdata_o;
	// Trace: design.sv:39892:3
	output reg out_err_o;
	// Trace: design.sv:39893:3
	output reg out_err_plus2_o;
	// Trace: design.sv:39896:3
	localparam [31:0] DEPTH = NUM_REQS + 1;
	// Trace: design.sv:39899:3
	wire [(DEPTH * 32) - 1:0] rdata_d;
	reg [(DEPTH * 32) - 1:0] rdata_q;
	// Trace: design.sv:39900:3
	wire [DEPTH - 1:0] err_d;
	reg [DEPTH - 1:0] err_q;
	// Trace: design.sv:39901:3
	wire [DEPTH - 1:0] valid_d;
	reg [DEPTH - 1:0] valid_q;
	// Trace: design.sv:39902:3
	wire [DEPTH - 1:0] lowest_free_entry;
	// Trace: design.sv:39903:3
	wire [DEPTH - 1:0] valid_pushed;
	wire [DEPTH - 1:0] valid_popped;
	// Trace: design.sv:39904:3
	wire [DEPTH - 1:0] entry_en;
	// Trace: design.sv:39906:3
	wire pop_fifo;
	// Trace: design.sv:39907:3
	wire [31:0] rdata;
	wire [31:0] rdata_unaligned;
	// Trace: design.sv:39908:3
	wire err;
	wire err_unaligned;
	wire err_plus2;
	// Trace: design.sv:39909:3
	wire valid;
	wire valid_unaligned;
	// Trace: design.sv:39911:3
	wire aligned_is_compressed;
	wire unaligned_is_compressed;
	// Trace: design.sv:39913:3
	wire addr_incr_two;
	// Trace: design.sv:39914:3
	wire [31:1] instr_addr_next;
	// Trace: design.sv:39915:3
	wire [31:1] instr_addr_d;
	reg [31:1] instr_addr_q;
	// Trace: design.sv:39916:3
	wire instr_addr_en;
	// Trace: design.sv:39917:3
	wire unused_addr_in;
	// Trace: design.sv:39923:3
	assign rdata = (valid_q[0] ? rdata_q[0+:32] : in_rdata_i);
	// Trace: design.sv:39924:3
	assign err = (valid_q[0] ? err_q[0] : in_err_i);
	// Trace: design.sv:39925:3
	assign valid = valid_q[0] | in_valid_i;
	// Trace: design.sv:39939:3
	assign rdata_unaligned = (valid_q[1] ? {rdata_q[47-:16], rdata[31:16]} : {in_rdata_i[15:0], rdata[31:16]});
	// Trace: design.sv:39947:3
	assign err_unaligned = (valid_q[1] ? (err_q[1] & ~unaligned_is_compressed) | err_q[0] : (valid_q[0] & err_q[0]) | (in_err_i & (~valid_q[0] | ~unaligned_is_compressed)));
	// Trace: design.sv:39953:3
	assign err_plus2 = (valid_q[1] ? err_q[1] & ~err_q[0] : (in_err_i & valid_q[0]) & ~err_q[0]);
	// Trace: design.sv:39957:3
	assign valid_unaligned = (valid_q[1] ? 1'b1 : valid_q[0] & in_valid_i);
	// Trace: design.sv:39961:3
	assign unaligned_is_compressed = (rdata[17:16] != 2'b11) & ~err;
	// Trace: design.sv:39962:3
	assign aligned_is_compressed = (rdata[1:0] != 2'b11) & ~err;
	// Trace: design.sv:39968:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:39969:5
		if (out_addr_o[1]) begin
			// Trace: design.sv:39971:7
			out_rdata_o = rdata_unaligned;
			// Trace: design.sv:39972:7
			out_err_o = err_unaligned;
			// Trace: design.sv:39973:7
			out_err_plus2_o = err_plus2;
			// Trace: design.sv:39975:7
			if (unaligned_is_compressed)
				// Trace: design.sv:39976:9
				out_valid_o = valid;
			else
				// Trace: design.sv:39978:9
				out_valid_o = valid_unaligned;
		end
		else begin
			// Trace: design.sv:39982:7
			out_rdata_o = rdata;
			// Trace: design.sv:39983:7
			out_err_o = err;
			// Trace: design.sv:39984:7
			out_err_plus2_o = 1'b0;
			// Trace: design.sv:39985:7
			out_valid_o = valid;
		end
	end
	// Trace: design.sv:39994:3
	assign instr_addr_en = clear_i | (out_ready_i & out_valid_o);
	// Trace: design.sv:39997:3
	assign addr_incr_two = (instr_addr_q[1] ? unaligned_is_compressed : aligned_is_compressed);
	// Trace: design.sv:40000:3
	assign instr_addr_next = instr_addr_q[31:1] + {29'd0, ~addr_incr_two, addr_incr_two};
	// Trace: design.sv:40004:3
	assign instr_addr_d = (clear_i ? in_addr_i[31:1] : instr_addr_next);
	// Trace: design.sv:40007:3
	generate
		if (ResetAll) begin : g_instr_addr_ra
			// Trace: design.sv:40008:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:40009:7
				if (!rst_ni)
					// Trace: design.sv:40010:9
					instr_addr_q <= 1'sb0;
				else if (instr_addr_en)
					// Trace: design.sv:40012:9
					instr_addr_q <= instr_addr_d;
		end
		else begin : g_instr_addr_nr
			// Trace: design.sv:40016:5
			always @(posedge clk_i)
				// Trace: design.sv:40017:7
				if (instr_addr_en)
					// Trace: design.sv:40018:9
					instr_addr_q <= instr_addr_d;
		end
	endgenerate
	// Trace: design.sv:40024:3
	assign out_addr_o = {instr_addr_q, 1'b0};
	// Trace: design.sv:40027:3
	assign unused_addr_in = in_addr_i[0];
	// Trace: design.sv:40036:3
	assign busy_o = valid_q[DEPTH - 1:DEPTH - NUM_REQS];
	// Trace: design.sv:40043:3
	assign pop_fifo = (out_ready_i & out_valid_o) & (~aligned_is_compressed | out_addr_o[1]);
	// Trace: design.sv:40045:3
	genvar _gv_i_64;
	generate
		for (_gv_i_64 = 0; _gv_i_64 < (DEPTH - 1); _gv_i_64 = _gv_i_64 + 1) begin : g_fifo_next
			localparam i = _gv_i_64;
			if (i == 0) begin : g_ent0
				// Trace: design.sv:40048:7
				assign lowest_free_entry[i] = ~valid_q[i];
			end
			else begin : g_ent_others
				// Trace: design.sv:40050:7
				assign lowest_free_entry[i] = ~valid_q[i] & valid_q[i - 1];
			end
			// Trace: design.sv:40054:5
			assign valid_pushed[i] = (in_valid_i & lowest_free_entry[i]) | valid_q[i];
			// Trace: design.sv:40057:5
			assign valid_popped[i] = (pop_fifo ? valid_pushed[i + 1] : valid_pushed[i]);
			// Trace: design.sv:40059:5
			assign valid_d[i] = valid_popped[i] & ~clear_i;
			// Trace: design.sv:40062:5
			assign entry_en[i] = (valid_pushed[i + 1] & pop_fifo) | ((in_valid_i & lowest_free_entry[i]) & ~pop_fifo);
			// Trace: design.sv:40067:5
			assign rdata_d[i * 32+:32] = (valid_q[i + 1] ? rdata_q[(i + 1) * 32+:32] : in_rdata_i);
			// Trace: design.sv:40068:5
			assign err_d[i] = (valid_q[i + 1] ? err_q[i + 1] : in_err_i);
		end
	endgenerate
	// Trace: design.sv:40071:3
	assign lowest_free_entry[DEPTH - 1] = ~valid_q[DEPTH - 1] & valid_q[DEPTH - 2];
	// Trace: design.sv:40072:3
	assign valid_pushed[DEPTH - 1] = valid_q[DEPTH - 1] | (in_valid_i & lowest_free_entry[DEPTH - 1]);
	// Trace: design.sv:40073:3
	assign valid_popped[DEPTH - 1] = (pop_fifo ? 1'b0 : valid_pushed[DEPTH - 1]);
	// Trace: design.sv:40074:3
	assign valid_d[DEPTH - 1] = valid_popped[DEPTH - 1] & ~clear_i;
	// Trace: design.sv:40075:3
	assign entry_en[DEPTH - 1] = in_valid_i & lowest_free_entry[DEPTH - 1];
	// Trace: design.sv:40076:3
	assign rdata_d[(DEPTH - 1) * 32+:32] = in_rdata_i;
	// Trace: design.sv:40077:3
	assign err_d[DEPTH - 1] = in_err_i;
	// Trace: design.sv:40083:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:40084:5
		if (!rst_ni)
			// Trace: design.sv:40085:7
			valid_q <= 1'sb0;
		else
			// Trace: design.sv:40087:7
			valid_q <= valid_d;
	// Trace: design.sv:40091:3
	genvar _gv_i_65;
	generate
		for (_gv_i_65 = 0; _gv_i_65 < DEPTH; _gv_i_65 = _gv_i_65 + 1) begin : g_fifo_regs
			localparam i = _gv_i_65;
			if (ResetAll) begin : g_rdata_ra
				// Trace: design.sv:40093:7
				always @(posedge clk_i or negedge rst_ni)
					// Trace: design.sv:40094:9
					if (!rst_ni) begin
						// Trace: design.sv:40095:11
						rdata_q[i * 32+:32] <= 1'sb0;
						// Trace: design.sv:40096:11
						err_q[i] <= 1'sb0;
					end
					else if (entry_en[i]) begin
						// Trace: design.sv:40098:11
						rdata_q[i * 32+:32] <= rdata_d[i * 32+:32];
						// Trace: design.sv:40099:11
						err_q[i] <= err_d[i];
					end
			end
			else begin : g_rdata_nr
				// Trace: design.sv:40103:7
				always @(posedge clk_i)
					// Trace: design.sv:40104:9
					if (entry_en[i]) begin
						// Trace: design.sv:40105:11
						rdata_q[i * 32+:32] <= rdata_d[i * 32+:32];
						// Trace: design.sv:40106:11
						err_q[i] <= err_d[i];
					end
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module ibex_id_stage (
	clk_i,
	rst_ni,
	ctrl_busy_o,
	illegal_insn_o,
	instr_valid_i,
	instr_rdata_i,
	instr_rdata_alu_i,
	instr_rdata_c_i,
	instr_is_compressed_i,
	instr_bp_taken_i,
	instr_req_o,
	instr_first_cycle_id_o,
	instr_valid_clear_o,
	id_in_ready_o,
	icache_inval_o,
	branch_decision_i,
	pc_set_o,
	pc_mux_o,
	nt_branch_mispredict_o,
	nt_branch_addr_o,
	exc_pc_mux_o,
	exc_cause_o,
	illegal_c_insn_i,
	instr_fetch_err_i,
	instr_fetch_err_plus2_i,
	pc_id_i,
	ex_valid_i,
	lsu_resp_valid_i,
	alu_operator_ex_o,
	alu_operand_a_ex_o,
	alu_operand_b_ex_o,
	imd_val_we_ex_i,
	imd_val_d_ex_i,
	imd_val_q_ex_o,
	bt_a_operand_o,
	bt_b_operand_o,
	mult_en_ex_o,
	div_en_ex_o,
	mult_sel_ex_o,
	div_sel_ex_o,
	multdiv_operator_ex_o,
	multdiv_signed_mode_ex_o,
	multdiv_operand_a_ex_o,
	multdiv_operand_b_ex_o,
	multdiv_ready_id_o,
	csr_access_o,
	csr_op_o,
	csr_op_en_o,
	csr_save_if_o,
	csr_save_id_o,
	csr_save_wb_o,
	csr_restore_mret_id_o,
	csr_restore_dret_id_o,
	csr_save_cause_o,
	csr_mtval_o,
	priv_mode_i,
	csr_mstatus_tw_i,
	illegal_csr_insn_i,
	data_ind_timing_i,
	lsu_req_o,
	lsu_we_o,
	lsu_type_o,
	lsu_sign_ext_o,
	lsu_wdata_o,
	lsu_req_done_i,
	lsu_addr_incr_req_i,
	lsu_addr_last_i,
	csr_mstatus_mie_i,
	irq_pending_i,
	irqs_i,
	irq_nm_i,
	nmi_mode_o,
	lsu_load_err_i,
	lsu_store_err_i,
	debug_mode_o,
	debug_cause_o,
	debug_csr_save_o,
	debug_req_i,
	debug_single_step_i,
	debug_ebreakm_i,
	debug_ebreaku_i,
	trigger_match_i,
	wake_from_sleep_o,
	result_ex_i,
	csr_rdata_i,
	rf_raddr_a_o,
	rf_rdata_a_i,
	rf_raddr_b_o,
	rf_rdata_b_i,
	rf_ren_a_o,
	rf_ren_b_o,
	rf_waddr_id_o,
	rf_wdata_id_o,
	rf_we_id_o,
	rf_rd_a_wb_match_o,
	rf_rd_b_wb_match_o,
	rf_waddr_wb_i,
	rf_wdata_fwd_wb_i,
	rf_write_wb_i,
	en_wb_o,
	instr_type_wb_o,
	instr_perf_count_id_o,
	ready_wb_i,
	outstanding_load_wb_i,
	outstanding_store_wb_i,
	perf_jump_o,
	perf_branch_o,
	perf_tbranch_o,
	perf_dside_wait_o,
	perf_mul_wait_o,
	perf_div_wait_o,
	instr_id_done_o
);
	reg _sv2v_0;
	// Trace: design.sv:40145:13
	parameter [0:0] RV32E = 0;
	// Trace: design.sv:40146:13
	// removed localparam type ibex_pkg_rv32m_e
	parameter integer RV32M = 32'sd2;
	// Trace: design.sv:40147:13
	// removed localparam type ibex_pkg_rv32b_e
	parameter integer RV32B = 32'sd0;
	// Trace: design.sv:40148:13
	parameter [0:0] DataIndTiming = 1'b0;
	// Trace: design.sv:40149:13
	parameter [0:0] BranchTargetALU = 0;
	// Trace: design.sv:40150:13
	parameter [0:0] WritebackStage = 0;
	// Trace: design.sv:40151:13
	parameter [0:0] BranchPredictor = 0;
	// Trace: design.sv:40153:3
	input wire clk_i;
	// Trace: design.sv:40154:3
	input wire rst_ni;
	// Trace: design.sv:40156:3
	output wire ctrl_busy_o;
	// Trace: design.sv:40157:3
	output wire illegal_insn_o;
	// Trace: design.sv:40160:3
	input wire instr_valid_i;
	// Trace: design.sv:40161:3
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:40162:3
	input wire [31:0] instr_rdata_alu_i;
	// Trace: design.sv:40163:3
	input wire [15:0] instr_rdata_c_i;
	// Trace: design.sv:40164:3
	input wire instr_is_compressed_i;
	// Trace: design.sv:40165:3
	input wire instr_bp_taken_i;
	// Trace: design.sv:40166:3
	output wire instr_req_o;
	// Trace: design.sv:40167:3
	output wire instr_first_cycle_id_o;
	// Trace: design.sv:40168:3
	output wire instr_valid_clear_o;
	// Trace: design.sv:40169:3
	output wire id_in_ready_o;
	// Trace: design.sv:40170:3
	output wire icache_inval_o;
	// Trace: design.sv:40173:3
	input wire branch_decision_i;
	// Trace: design.sv:40176:3
	output wire pc_set_o;
	// Trace: design.sv:40177:3
	// removed localparam type ibex_pkg_pc_sel_e
	output wire [2:0] pc_mux_o;
	// Trace: design.sv:40178:3
	output wire nt_branch_mispredict_o;
	// Trace: design.sv:40179:3
	output wire [31:0] nt_branch_addr_o;
	// Trace: design.sv:40180:3
	// removed localparam type ibex_pkg_exc_pc_sel_e
	output wire [1:0] exc_pc_mux_o;
	// Trace: design.sv:40181:3
	// removed localparam type ibex_pkg_exc_cause_e
	output wire [5:0] exc_cause_o;
	// Trace: design.sv:40183:3
	input wire illegal_c_insn_i;
	// Trace: design.sv:40184:3
	input wire instr_fetch_err_i;
	// Trace: design.sv:40185:3
	input wire instr_fetch_err_plus2_i;
	// Trace: design.sv:40187:3
	input wire [31:0] pc_id_i;
	// Trace: design.sv:40190:3
	input wire ex_valid_i;
	// Trace: design.sv:40191:3
	input wire lsu_resp_valid_i;
	// Trace: design.sv:40193:3
	// removed localparam type ibex_pkg_alu_op_e
	output wire [6:0] alu_operator_ex_o;
	// Trace: design.sv:40194:3
	output wire [31:0] alu_operand_a_ex_o;
	// Trace: design.sv:40195:3
	output wire [31:0] alu_operand_b_ex_o;
	// Trace: design.sv:40198:3
	input wire [1:0] imd_val_we_ex_i;
	// Trace: design.sv:40199:3
	input wire [67:0] imd_val_d_ex_i;
	// Trace: design.sv:40200:3
	output wire [67:0] imd_val_q_ex_o;
	// Trace: design.sv:40203:3
	output reg [31:0] bt_a_operand_o;
	// Trace: design.sv:40204:3
	output reg [31:0] bt_b_operand_o;
	// Trace: design.sv:40207:3
	output wire mult_en_ex_o;
	// Trace: design.sv:40208:3
	output wire div_en_ex_o;
	// Trace: design.sv:40209:3
	output wire mult_sel_ex_o;
	// Trace: design.sv:40210:3
	output wire div_sel_ex_o;
	// Trace: design.sv:40211:3
	// removed localparam type ibex_pkg_md_op_e
	output wire [1:0] multdiv_operator_ex_o;
	// Trace: design.sv:40212:3
	output wire [1:0] multdiv_signed_mode_ex_o;
	// Trace: design.sv:40213:3
	output wire [31:0] multdiv_operand_a_ex_o;
	// Trace: design.sv:40214:3
	output wire [31:0] multdiv_operand_b_ex_o;
	// Trace: design.sv:40215:3
	output wire multdiv_ready_id_o;
	// Trace: design.sv:40218:3
	output wire csr_access_o;
	// Trace: design.sv:40219:3
	// removed localparam type ibex_pkg_csr_op_e
	output wire [1:0] csr_op_o;
	// Trace: design.sv:40220:3
	output wire csr_op_en_o;
	// Trace: design.sv:40221:3
	output wire csr_save_if_o;
	// Trace: design.sv:40222:3
	output wire csr_save_id_o;
	// Trace: design.sv:40223:3
	output wire csr_save_wb_o;
	// Trace: design.sv:40224:3
	output wire csr_restore_mret_id_o;
	// Trace: design.sv:40225:3
	output wire csr_restore_dret_id_o;
	// Trace: design.sv:40226:3
	output wire csr_save_cause_o;
	// Trace: design.sv:40227:3
	output wire [31:0] csr_mtval_o;
	// Trace: design.sv:40228:3
	// removed localparam type ibex_pkg_priv_lvl_e
	input wire [1:0] priv_mode_i;
	// Trace: design.sv:40229:3
	input wire csr_mstatus_tw_i;
	// Trace: design.sv:40230:3
	input wire illegal_csr_insn_i;
	// Trace: design.sv:40231:3
	input wire data_ind_timing_i;
	// Trace: design.sv:40234:3
	output wire lsu_req_o;
	// Trace: design.sv:40235:3
	output wire lsu_we_o;
	// Trace: design.sv:40236:3
	output wire [1:0] lsu_type_o;
	// Trace: design.sv:40237:3
	output wire lsu_sign_ext_o;
	// Trace: design.sv:40238:3
	output wire [31:0] lsu_wdata_o;
	// Trace: design.sv:40240:3
	input wire lsu_req_done_i;
	// Trace: design.sv:40245:3
	input wire lsu_addr_incr_req_i;
	// Trace: design.sv:40246:3
	input wire [31:0] lsu_addr_last_i;
	// Trace: design.sv:40249:3
	input wire csr_mstatus_mie_i;
	// Trace: design.sv:40250:3
	input wire irq_pending_i;
	// Trace: design.sv:40251:3
	// removed localparam type ibex_pkg_irqs_t
	input wire [17:0] irqs_i;
	// Trace: design.sv:40252:3
	input wire irq_nm_i;
	// Trace: design.sv:40253:3
	output wire nmi_mode_o;
	// Trace: design.sv:40255:3
	input wire lsu_load_err_i;
	// Trace: design.sv:40256:3
	input wire lsu_store_err_i;
	// Trace: design.sv:40259:3
	output wire debug_mode_o;
	// Trace: design.sv:40260:3
	// removed localparam type ibex_pkg_dbg_cause_e
	output wire [2:0] debug_cause_o;
	// Trace: design.sv:40261:3
	output wire debug_csr_save_o;
	// Trace: design.sv:40262:3
	input wire debug_req_i;
	// Trace: design.sv:40263:3
	input wire debug_single_step_i;
	// Trace: design.sv:40264:3
	input wire debug_ebreakm_i;
	// Trace: design.sv:40265:3
	input wire debug_ebreaku_i;
	// Trace: design.sv:40266:3
	input wire trigger_match_i;
	// Trace: design.sv:40269:3
	output wire wake_from_sleep_o;
	// Trace: design.sv:40272:3
	input wire [31:0] result_ex_i;
	// Trace: design.sv:40273:3
	input wire [31:0] csr_rdata_i;
	// Trace: design.sv:40276:3
	output wire [4:0] rf_raddr_a_o;
	// Trace: design.sv:40277:3
	input wire [31:0] rf_rdata_a_i;
	// Trace: design.sv:40278:3
	output wire [4:0] rf_raddr_b_o;
	// Trace: design.sv:40279:3
	input wire [31:0] rf_rdata_b_i;
	// Trace: design.sv:40280:3
	output wire rf_ren_a_o;
	// Trace: design.sv:40281:3
	output wire rf_ren_b_o;
	// Trace: design.sv:40284:3
	output wire [4:0] rf_waddr_id_o;
	// Trace: design.sv:40285:3
	output reg [31:0] rf_wdata_id_o;
	// Trace: design.sv:40286:3
	output wire rf_we_id_o;
	// Trace: design.sv:40287:3
	output wire rf_rd_a_wb_match_o;
	// Trace: design.sv:40288:3
	output wire rf_rd_b_wb_match_o;
	// Trace: design.sv:40291:3
	input wire [4:0] rf_waddr_wb_i;
	// Trace: design.sv:40292:3
	input wire [31:0] rf_wdata_fwd_wb_i;
	// Trace: design.sv:40293:3
	input wire rf_write_wb_i;
	// Trace: design.sv:40295:3
	output wire en_wb_o;
	// Trace: design.sv:40296:3
	// removed localparam type ibex_pkg_wb_instr_type_e
	output wire [1:0] instr_type_wb_o;
	// Trace: design.sv:40297:3
	output wire instr_perf_count_id_o;
	// Trace: design.sv:40298:3
	input wire ready_wb_i;
	// Trace: design.sv:40299:3
	input wire outstanding_load_wb_i;
	// Trace: design.sv:40300:3
	input wire outstanding_store_wb_i;
	// Trace: design.sv:40303:3
	output wire perf_jump_o;
	// Trace: design.sv:40304:3
	output reg perf_branch_o;
	// Trace: design.sv:40305:3
	output wire perf_tbranch_o;
	// Trace: design.sv:40306:3
	output wire perf_dside_wait_o;
	// Trace: design.sv:40308:3
	output wire perf_mul_wait_o;
	// Trace: design.sv:40309:3
	output wire perf_div_wait_o;
	// Trace: design.sv:40310:3
	output wire instr_id_done_o;
	// Trace: design.sv:40313:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:40316:3
	wire illegal_insn_dec;
	// Trace: design.sv:40317:3
	wire ebrk_insn;
	// Trace: design.sv:40318:3
	wire mret_insn_dec;
	// Trace: design.sv:40319:3
	wire dret_insn_dec;
	// Trace: design.sv:40320:3
	wire ecall_insn_dec;
	// Trace: design.sv:40321:3
	wire wfi_insn_dec;
	// Trace: design.sv:40323:3
	wire wb_exception;
	// Trace: design.sv:40324:3
	wire id_exception;
	// Trace: design.sv:40326:3
	wire branch_in_dec;
	// Trace: design.sv:40327:3
	wire branch_set;
	wire branch_set_raw;
	reg branch_set_raw_d;
	// Trace: design.sv:40328:3
	reg branch_jump_set_done_q;
	wire branch_jump_set_done_d;
	// Trace: design.sv:40329:3
	reg branch_not_set;
	// Trace: design.sv:40330:3
	wire branch_taken;
	// Trace: design.sv:40331:3
	wire jump_in_dec;
	// Trace: design.sv:40332:3
	wire jump_set_dec;
	// Trace: design.sv:40333:3
	wire jump_set;
	reg jump_set_raw;
	// Trace: design.sv:40335:3
	wire instr_first_cycle;
	// Trace: design.sv:40336:3
	wire instr_executing_spec;
	// Trace: design.sv:40337:3
	wire instr_executing;
	// Trace: design.sv:40338:3
	wire instr_done;
	// Trace: design.sv:40339:3
	wire controller_run;
	// Trace: design.sv:40340:3
	wire stall_ld_hz;
	// Trace: design.sv:40341:3
	wire stall_mem;
	// Trace: design.sv:40342:3
	reg stall_multdiv;
	// Trace: design.sv:40343:3
	reg stall_branch;
	// Trace: design.sv:40344:3
	reg stall_jump;
	// Trace: design.sv:40345:3
	wire stall_id;
	// Trace: design.sv:40346:3
	wire stall_wb;
	// Trace: design.sv:40347:3
	wire flush_id;
	// Trace: design.sv:40348:3
	wire multicycle_done;
	// Trace: design.sv:40351:3
	wire [31:0] imm_i_type;
	// Trace: design.sv:40352:3
	wire [31:0] imm_s_type;
	// Trace: design.sv:40353:3
	wire [31:0] imm_b_type;
	// Trace: design.sv:40354:3
	wire [31:0] imm_u_type;
	// Trace: design.sv:40355:3
	wire [31:0] imm_j_type;
	// Trace: design.sv:40356:3
	wire [31:0] zimm_rs1_type;
	// Trace: design.sv:40358:3
	wire [31:0] imm_a;
	// Trace: design.sv:40359:3
	reg [31:0] imm_b;
	// Trace: design.sv:40363:3
	// removed localparam type ibex_pkg_rf_wd_sel_e
	wire rf_wdata_sel;
	// Trace: design.sv:40364:3
	wire rf_we_dec;
	reg rf_we_raw;
	// Trace: design.sv:40365:3
	wire rf_ren_a;
	wire rf_ren_b;
	// Trace: design.sv:40366:3
	wire rf_ren_a_dec;
	wire rf_ren_b_dec;
	// Trace: design.sv:40369:3
	assign rf_ren_a = ((instr_valid_i & ~instr_fetch_err_i) & ~illegal_insn_o) & rf_ren_a_dec;
	// Trace: design.sv:40370:3
	assign rf_ren_b = ((instr_valid_i & ~instr_fetch_err_i) & ~illegal_insn_o) & rf_ren_b_dec;
	// Trace: design.sv:40372:3
	assign rf_ren_a_o = rf_ren_a;
	// Trace: design.sv:40373:3
	assign rf_ren_b_o = rf_ren_b;
	// Trace: design.sv:40375:3
	wire [31:0] rf_rdata_a_fwd;
	// Trace: design.sv:40376:3
	wire [31:0] rf_rdata_b_fwd;
	// Trace: design.sv:40379:3
	wire [6:0] alu_operator;
	// Trace: design.sv:40380:3
	// removed localparam type ibex_pkg_op_a_sel_e
	wire [1:0] alu_op_a_mux_sel;
	wire [1:0] alu_op_a_mux_sel_dec;
	// Trace: design.sv:40381:3
	// removed localparam type ibex_pkg_op_b_sel_e
	wire alu_op_b_mux_sel;
	wire alu_op_b_mux_sel_dec;
	// Trace: design.sv:40382:3
	wire alu_multicycle_dec;
	// Trace: design.sv:40383:3
	reg stall_alu;
	// Trace: design.sv:40385:3
	reg [67:0] imd_val_q;
	// Trace: design.sv:40387:3
	wire [1:0] bt_a_mux_sel;
	// Trace: design.sv:40388:3
	// removed localparam type ibex_pkg_imm_b_sel_e
	wire [2:0] bt_b_mux_sel;
	// Trace: design.sv:40390:3
	// removed localparam type ibex_pkg_imm_a_sel_e
	wire imm_a_mux_sel;
	// Trace: design.sv:40391:3
	wire [2:0] imm_b_mux_sel;
	wire [2:0] imm_b_mux_sel_dec;
	// Trace: design.sv:40394:3
	wire mult_en_id;
	wire mult_en_dec;
	// Trace: design.sv:40395:3
	wire div_en_id;
	wire div_en_dec;
	// Trace: design.sv:40396:3
	wire multdiv_en_dec;
	// Trace: design.sv:40397:3
	wire [1:0] multdiv_operator;
	// Trace: design.sv:40398:3
	wire [1:0] multdiv_signed_mode;
	// Trace: design.sv:40401:3
	wire lsu_we;
	// Trace: design.sv:40402:3
	wire [1:0] lsu_type;
	// Trace: design.sv:40403:3
	wire lsu_sign_ext;
	// Trace: design.sv:40404:3
	wire lsu_req;
	wire lsu_req_dec;
	// Trace: design.sv:40405:3
	wire data_req_allowed;
	// Trace: design.sv:40408:3
	reg csr_pipe_flush;
	// Trace: design.sv:40410:3
	reg [31:0] alu_operand_a;
	// Trace: design.sv:40411:3
	wire [31:0] alu_operand_b;
	// Trace: design.sv:40418:3
	assign alu_op_a_mux_sel = (lsu_addr_incr_req_i ? 2'd1 : alu_op_a_mux_sel_dec);
	// Trace: design.sv:40419:3
	assign alu_op_b_mux_sel = (lsu_addr_incr_req_i ? 1'd1 : alu_op_b_mux_sel_dec);
	// Trace: design.sv:40420:3
	assign imm_b_mux_sel = (lsu_addr_incr_req_i ? 3'd6 : imm_b_mux_sel_dec);
	// Trace: design.sv:40427:3
	assign imm_a = (imm_a_mux_sel == 1'd0 ? zimm_rs1_type : {32 {1'sb0}});
	// Trace: design.sv:40430:3
	always @(*) begin : alu_operand_a_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:40431:5
		(* full_case, parallel_case *)
		case (alu_op_a_mux_sel)
			2'd0:
				// Trace: design.sv:40432:20
				alu_operand_a = rf_rdata_a_fwd;
			2'd1:
				// Trace: design.sv:40433:20
				alu_operand_a = lsu_addr_last_i;
			2'd2:
				// Trace: design.sv:40434:20
				alu_operand_a = pc_id_i;
			2'd3:
				// Trace: design.sv:40435:20
				alu_operand_a = imm_a;
			default:
				// Trace: design.sv:40436:20
				alu_operand_a = pc_id_i;
		endcase
	end
	// Trace: design.sv:40440:3
	generate
		if (BranchTargetALU) begin : g_btalu_muxes
			// Trace: design.sv:40442:5
			always @(*) begin : bt_operand_a_mux
				if (_sv2v_0)
					;
				// Trace: design.sv:40443:7
				(* full_case, parallel_case *)
				case (bt_a_mux_sel)
					2'd0:
						// Trace: design.sv:40444:22
						bt_a_operand_o = rf_rdata_a_fwd;
					2'd2:
						// Trace: design.sv:40445:22
						bt_a_operand_o = pc_id_i;
					default:
						// Trace: design.sv:40446:22
						bt_a_operand_o = pc_id_i;
				endcase
			end
			// Trace: design.sv:40451:5
			always @(*) begin : bt_immediate_b_mux
				if (_sv2v_0)
					;
				// Trace: design.sv:40452:7
				(* full_case, parallel_case *)
				case (bt_b_mux_sel)
					3'd0:
						// Trace: design.sv:40453:26
						bt_b_operand_o = imm_i_type;
					3'd2:
						// Trace: design.sv:40454:26
						bt_b_operand_o = imm_b_type;
					3'd4:
						// Trace: design.sv:40455:26
						bt_b_operand_o = imm_j_type;
					3'd5:
						// Trace: design.sv:40456:26
						bt_b_operand_o = (instr_is_compressed_i ? 32'h00000002 : 32'h00000004);
					default:
						// Trace: design.sv:40457:26
						bt_b_operand_o = (instr_is_compressed_i ? 32'h00000002 : 32'h00000004);
				endcase
			end
			// Trace: design.sv:40462:5
			always @(*) begin : immediate_b_mux
				if (_sv2v_0)
					;
				// Trace: design.sv:40463:7
				(* full_case, parallel_case *)
				case (imm_b_mux_sel)
					3'd0:
						// Trace: design.sv:40464:26
						imm_b = imm_i_type;
					3'd1:
						// Trace: design.sv:40465:26
						imm_b = imm_s_type;
					3'd3:
						// Trace: design.sv:40466:26
						imm_b = imm_u_type;
					3'd5:
						// Trace: design.sv:40467:26
						imm_b = (instr_is_compressed_i ? 32'h00000002 : 32'h00000004);
					3'd6:
						// Trace: design.sv:40468:26
						imm_b = 32'h00000004;
					default:
						// Trace: design.sv:40469:26
						imm_b = 32'h00000004;
				endcase
			end
		end
		else begin : g_nobtalu
			// Trace: design.sv:40479:5
			wire [1:0] unused_a_mux_sel;
			// Trace: design.sv:40480:5
			wire [2:0] unused_b_mux_sel;
			// Trace: design.sv:40482:5
			assign unused_a_mux_sel = bt_a_mux_sel;
			// Trace: design.sv:40483:5
			assign unused_b_mux_sel = bt_b_mux_sel;
			// Trace: design.sv:40484:5
			wire [32:1] sv2v_tmp_1FCCD;
			assign sv2v_tmp_1FCCD = 1'sb0;
			always @(*) bt_a_operand_o = sv2v_tmp_1FCCD;
			// Trace: design.sv:40485:5
			wire [32:1] sv2v_tmp_B876E;
			assign sv2v_tmp_B876E = 1'sb0;
			always @(*) bt_b_operand_o = sv2v_tmp_B876E;
			// Trace: design.sv:40488:5
			always @(*) begin : immediate_b_mux
				if (_sv2v_0)
					;
				// Trace: design.sv:40489:7
				(* full_case, parallel_case *)
				case (imm_b_mux_sel)
					3'd0:
						// Trace: design.sv:40490:26
						imm_b = imm_i_type;
					3'd1:
						// Trace: design.sv:40491:26
						imm_b = imm_s_type;
					3'd2:
						// Trace: design.sv:40492:26
						imm_b = imm_b_type;
					3'd3:
						// Trace: design.sv:40493:26
						imm_b = imm_u_type;
					3'd4:
						// Trace: design.sv:40494:26
						imm_b = imm_j_type;
					3'd5:
						// Trace: design.sv:40495:26
						imm_b = (instr_is_compressed_i ? 32'h00000002 : 32'h00000004);
					3'd6:
						// Trace: design.sv:40496:26
						imm_b = 32'h00000004;
					default:
						// Trace: design.sv:40497:26
						imm_b = 32'h00000004;
				endcase
			end
		end
	endgenerate
	// Trace: design.sv:40511:3
	assign alu_operand_b = (alu_op_b_mux_sel == 1'd1 ? imm_b : rf_rdata_b_fwd);
	// Trace: design.sv:40517:3
	genvar _gv_i_66;
	generate
		for (_gv_i_66 = 0; _gv_i_66 < 2; _gv_i_66 = _gv_i_66 + 1) begin : gen_intermediate_val_reg
			localparam i = _gv_i_66;
			// Trace: design.sv:40518:5
			always @(posedge clk_i or negedge rst_ni) begin : intermediate_val_reg
				// Trace: design.sv:40519:7
				if (!rst_ni)
					// Trace: design.sv:40520:9
					imd_val_q[(1 - i) * 34+:34] <= 1'sb0;
				else if (imd_val_we_ex_i[i])
					// Trace: design.sv:40522:9
					imd_val_q[(1 - i) * 34+:34] <= imd_val_d_ex_i[(1 - i) * 34+:34];
			end
		end
	endgenerate
	// Trace: design.sv:40527:3
	assign imd_val_q_ex_o = imd_val_q;
	// Trace: design.sv:40534:3
	assign rf_we_id_o = (rf_we_raw & instr_executing) & ~illegal_csr_insn_i;
	// Trace: design.sv:40537:3
	always @(*) begin : rf_wdata_id_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:40538:5
		(* full_case, parallel_case *)
		case (rf_wdata_sel)
			1'd0:
				// Trace: design.sv:40539:18
				rf_wdata_id_o = result_ex_i;
			1'd1:
				// Trace: design.sv:40540:18
				rf_wdata_id_o = csr_rdata_i;
			default:
				// Trace: design.sv:40541:18
				rf_wdata_id_o = result_ex_i;
		endcase
	end
	// Trace: design.sv:40549:3
	ibex_decoder #(
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU)
	) decoder_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.illegal_insn_o(illegal_insn_dec),
		.ebrk_insn_o(ebrk_insn),
		.mret_insn_o(mret_insn_dec),
		.dret_insn_o(dret_insn_dec),
		.ecall_insn_o(ecall_insn_dec),
		.wfi_insn_o(wfi_insn_dec),
		.jump_set_o(jump_set_dec),
		.branch_taken_i(branch_taken),
		.icache_inval_o(icache_inval_o),
		.instr_first_cycle_i(instr_first_cycle),
		.instr_rdata_i(instr_rdata_i),
		.instr_rdata_alu_i(instr_rdata_alu_i),
		.illegal_c_insn_i(illegal_c_insn_i),
		.imm_a_mux_sel_o(imm_a_mux_sel),
		.imm_b_mux_sel_o(imm_b_mux_sel_dec),
		.bt_a_mux_sel_o(bt_a_mux_sel),
		.bt_b_mux_sel_o(bt_b_mux_sel),
		.imm_i_type_o(imm_i_type),
		.imm_s_type_o(imm_s_type),
		.imm_b_type_o(imm_b_type),
		.imm_u_type_o(imm_u_type),
		.imm_j_type_o(imm_j_type),
		.zimm_rs1_type_o(zimm_rs1_type),
		.rf_wdata_sel_o(rf_wdata_sel),
		.rf_we_o(rf_we_dec),
		.rf_raddr_a_o(rf_raddr_a_o),
		.rf_raddr_b_o(rf_raddr_b_o),
		.rf_waddr_o(rf_waddr_id_o),
		.rf_ren_a_o(rf_ren_a_dec),
		.rf_ren_b_o(rf_ren_b_dec),
		.alu_operator_o(alu_operator),
		.alu_op_a_mux_sel_o(alu_op_a_mux_sel_dec),
		.alu_op_b_mux_sel_o(alu_op_b_mux_sel_dec),
		.alu_multicycle_o(alu_multicycle_dec),
		.mult_en_o(mult_en_dec),
		.div_en_o(div_en_dec),
		.mult_sel_o(mult_sel_ex_o),
		.div_sel_o(div_sel_ex_o),
		.multdiv_operator_o(multdiv_operator),
		.multdiv_signed_mode_o(multdiv_signed_mode),
		.csr_access_o(csr_access_o),
		.csr_op_o(csr_op_o),
		.data_req_o(lsu_req_dec),
		.data_we_o(lsu_we),
		.data_type_o(lsu_type),
		.data_sign_extension_o(lsu_sign_ext),
		.jump_in_dec_o(jump_in_dec),
		.branch_in_dec_o(branch_in_dec)
	);
	// Trace: design.sv:40630:3
	// removed localparam type ibex_pkg_csr_num_e
	always @(*) begin : csr_pipeline_flushes
		if (_sv2v_0)
			;
		// Trace: design.sv:40631:5
		csr_pipe_flush = 1'b0;
		// Trace: design.sv:40638:5
		if ((csr_op_en_o == 1'b1) && ((csr_op_o == 2'd1) || (csr_op_o == 2'd2))) begin
			begin
				// Trace: design.sv:40639:7
				if ((instr_rdata_i[31:20] == 12'h300) || (instr_rdata_i[31:20] == 12'h304))
					// Trace: design.sv:40641:9
					csr_pipe_flush = 1'b1;
			end
		end
		else if ((csr_op_en_o == 1'b1) && (csr_op_o != 2'd0)) begin
			begin
				// Trace: design.sv:40644:7
				if ((((instr_rdata_i[31:20] == 12'h7b0) || (instr_rdata_i[31:20] == 12'h7b1)) || (instr_rdata_i[31:20] == 12'h7b2)) || (instr_rdata_i[31:20] == 12'h7b3))
					// Trace: design.sv:40648:9
					csr_pipe_flush = 1'b1;
			end
		end
	end
	// Trace: design.sv:40657:3
	assign illegal_insn_o = instr_valid_i & (illegal_insn_dec | illegal_csr_insn_i);
	// Trace: design.sv:40659:3
	ibex_controller #(
		.WritebackStage(WritebackStage),
		.BranchPredictor(BranchPredictor)
	) controller_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.ctrl_busy_o(ctrl_busy_o),
		.illegal_insn_i(illegal_insn_o),
		.ecall_insn_i(ecall_insn_dec),
		.mret_insn_i(mret_insn_dec),
		.dret_insn_i(dret_insn_dec),
		.wfi_insn_i(wfi_insn_dec),
		.ebrk_insn_i(ebrk_insn),
		.csr_pipe_flush_i(csr_pipe_flush),
		.instr_valid_i(instr_valid_i),
		.instr_i(instr_rdata_i),
		.instr_compressed_i(instr_rdata_c_i),
		.instr_is_compressed_i(instr_is_compressed_i),
		.instr_bp_taken_i(instr_bp_taken_i),
		.instr_fetch_err_i(instr_fetch_err_i),
		.instr_fetch_err_plus2_i(instr_fetch_err_plus2_i),
		.pc_id_i(pc_id_i),
		.instr_valid_clear_o(instr_valid_clear_o),
		.id_in_ready_o(id_in_ready_o),
		.controller_run_o(controller_run),
		.instr_req_o(instr_req_o),
		.pc_set_o(pc_set_o),
		.pc_mux_o(pc_mux_o),
		.nt_branch_mispredict_o(nt_branch_mispredict_o),
		.exc_pc_mux_o(exc_pc_mux_o),
		.exc_cause_o(exc_cause_o),
		.lsu_addr_last_i(lsu_addr_last_i),
		.load_err_i(lsu_load_err_i),
		.store_err_i(lsu_store_err_i),
		.wb_exception_o(wb_exception),
		.id_exception_o(id_exception),
		.branch_set_i(branch_set),
		.branch_not_set_i(branch_not_set),
		.jump_set_i(jump_set),
		.csr_mstatus_mie_i(csr_mstatus_mie_i),
		.irq_pending_i(irq_pending_i),
		.irqs_i(irqs_i),
		.irq_nm_i(irq_nm_i),
		.nmi_mode_o(nmi_mode_o),
		.csr_save_if_o(csr_save_if_o),
		.csr_save_id_o(csr_save_id_o),
		.csr_save_wb_o(csr_save_wb_o),
		.csr_restore_mret_id_o(csr_restore_mret_id_o),
		.csr_restore_dret_id_o(csr_restore_dret_id_o),
		.csr_save_cause_o(csr_save_cause_o),
		.csr_mtval_o(csr_mtval_o),
		.priv_mode_i(priv_mode_i),
		.csr_mstatus_tw_i(csr_mstatus_tw_i),
		.debug_mode_o(debug_mode_o),
		.debug_cause_o(debug_cause_o),
		.debug_csr_save_o(debug_csr_save_o),
		.debug_req_i(debug_req_i),
		.debug_single_step_i(debug_single_step_i),
		.debug_ebreakm_i(debug_ebreakm_i),
		.debug_ebreaku_i(debug_ebreaku_i),
		.trigger_match_i(trigger_match_i),
		.wake_from_sleep_o(wake_from_sleep_o),
		.stall_id_i(stall_id),
		.stall_wb_i(stall_wb),
		.flush_id_o(flush_id),
		.ready_wb_i(ready_wb_i),
		.perf_jump_o(perf_jump_o),
		.perf_tbranch_o(perf_tbranch_o)
	);
	// Trace: design.sv:40753:3
	assign multdiv_en_dec = mult_en_dec | div_en_dec;
	// Trace: design.sv:40755:3
	assign lsu_req = (instr_executing ? data_req_allowed & lsu_req_dec : 1'b0);
	// Trace: design.sv:40756:3
	assign mult_en_id = (instr_executing ? mult_en_dec : 1'b0);
	// Trace: design.sv:40757:3
	assign div_en_id = (instr_executing ? div_en_dec : 1'b0);
	// Trace: design.sv:40759:3
	assign lsu_req_o = lsu_req;
	// Trace: design.sv:40760:3
	assign lsu_we_o = lsu_we;
	// Trace: design.sv:40761:3
	assign lsu_type_o = lsu_type;
	// Trace: design.sv:40762:3
	assign lsu_sign_ext_o = lsu_sign_ext;
	// Trace: design.sv:40763:3
	assign lsu_wdata_o = rf_rdata_b_fwd;
	// Trace: design.sv:40768:3
	assign csr_op_en_o = (csr_access_o & instr_executing) & instr_id_done_o;
	// Trace: design.sv:40770:3
	assign alu_operator_ex_o = alu_operator;
	// Trace: design.sv:40771:3
	assign alu_operand_a_ex_o = alu_operand_a;
	// Trace: design.sv:40772:3
	assign alu_operand_b_ex_o = alu_operand_b;
	// Trace: design.sv:40774:3
	assign mult_en_ex_o = mult_en_id;
	// Trace: design.sv:40775:3
	assign div_en_ex_o = div_en_id;
	// Trace: design.sv:40777:3
	assign multdiv_operator_ex_o = multdiv_operator;
	// Trace: design.sv:40778:3
	assign multdiv_signed_mode_ex_o = multdiv_signed_mode;
	// Trace: design.sv:40779:3
	assign multdiv_operand_a_ex_o = rf_rdata_a_fwd;
	// Trace: design.sv:40780:3
	assign multdiv_operand_b_ex_o = rf_rdata_b_fwd;
	// Trace: design.sv:40786:3
	generate
		if (BranchTargetALU && !DataIndTiming) begin : g_branch_set_direct
			// Trace: design.sv:40789:5
			assign branch_set_raw = branch_set_raw_d;
		end
		else begin : g_branch_set_flop
			// Trace: design.sv:40794:5
			reg branch_set_raw_q;
			// Trace: design.sv:40796:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:40797:7
				if (!rst_ni)
					// Trace: design.sv:40798:9
					branch_set_raw_q <= 1'b0;
				else
					// Trace: design.sv:40800:9
					branch_set_raw_q <= branch_set_raw_d;
			// Trace: design.sv:40807:5
			assign branch_set_raw = (BranchTargetALU && !data_ind_timing_i ? branch_set_raw_d : branch_set_raw_q);
		end
	endgenerate
	// Trace: design.sv:40813:3
	assign branch_jump_set_done_d = ((branch_set_raw | jump_set_raw) | branch_jump_set_done_q) & ~instr_valid_clear_o;
	// Trace: design.sv:40816:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:40817:5
		if (!rst_ni)
			// Trace: design.sv:40818:7
			branch_jump_set_done_q <= 1'b0;
		else
			// Trace: design.sv:40820:7
			branch_jump_set_done_q <= branch_jump_set_done_d;
	// Trace: design.sv:40831:3
	assign jump_set = jump_set_raw & ~branch_jump_set_done_q;
	// Trace: design.sv:40832:3
	assign branch_set = branch_set_raw & ~branch_jump_set_done_q;
	// Trace: design.sv:40836:3
	generate
		if (DataIndTiming) begin : g_sec_branch_taken
			// Trace: design.sv:40838:5
			reg branch_taken_q;
			// Trace: design.sv:40840:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:40841:7
				if (!rst_ni)
					// Trace: design.sv:40842:9
					branch_taken_q <= 1'b0;
				else
					// Trace: design.sv:40844:9
					branch_taken_q <= branch_decision_i;
			// Trace: design.sv:40848:5
			assign branch_taken = ~data_ind_timing_i | branch_taken_q;
		end
		else begin : g_nosec_branch_taken
			// Trace: design.sv:40854:5
			assign branch_taken = 1'b1;
		end
	endgenerate
	// Trace: design.sv:40868:3
	generate
		if (BranchPredictor) begin : g_calc_nt_addr
			// Trace: design.sv:40869:5
			assign nt_branch_addr_o = pc_id_i + (instr_is_compressed_i ? 32'd2 : 32'd4);
		end
		else begin : g_n_calc_nt_addr
			// Trace: design.sv:40871:5
			assign nt_branch_addr_o = 32'd0;
		end
	endgenerate
	// Trace: design.sv:40878:3
	// removed localparam type id_fsm_e
	// Trace: design.sv:40879:3
	reg id_fsm_q;
	reg id_fsm_d;
	// Trace: design.sv:40881:3
	always @(posedge clk_i or negedge rst_ni) begin : id_pipeline_reg
		// Trace: design.sv:40882:5
		if (!rst_ni)
			// Trace: design.sv:40883:7
			id_fsm_q <= 1'd0;
		else if (instr_executing)
			// Trace: design.sv:40885:7
			id_fsm_q <= id_fsm_d;
	end
	// Trace: design.sv:40894:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:40895:5
		id_fsm_d = id_fsm_q;
		// Trace: design.sv:40896:5
		rf_we_raw = rf_we_dec;
		// Trace: design.sv:40897:5
		stall_multdiv = 1'b0;
		// Trace: design.sv:40898:5
		stall_jump = 1'b0;
		// Trace: design.sv:40899:5
		stall_branch = 1'b0;
		// Trace: design.sv:40900:5
		stall_alu = 1'b0;
		// Trace: design.sv:40901:5
		branch_set_raw_d = 1'b0;
		// Trace: design.sv:40902:5
		branch_not_set = 1'b0;
		// Trace: design.sv:40903:5
		jump_set_raw = 1'b0;
		// Trace: design.sv:40904:5
		perf_branch_o = 1'b0;
		// Trace: design.sv:40906:5
		if (instr_executing_spec)
			// Trace: design.sv:40907:7
			(* full_case, parallel_case *)
			case (id_fsm_q)
				1'd0:
					// Trace: design.sv:40909:11
					(* full_case, parallel_case *)
					case (1'b1)
						lsu_req_dec:
							// Trace: design.sv:40911:15
							if (!WritebackStage)
								// Trace: design.sv:40913:17
								id_fsm_d = 1'd1;
							else
								// Trace: design.sv:40915:17
								if (~lsu_req_done_i)
									// Trace: design.sv:40916:19
									id_fsm_d = 1'd1;
						multdiv_en_dec:
							// Trace: design.sv:40922:15
							if (~ex_valid_i) begin
								// Trace: design.sv:40925:17
								id_fsm_d = 1'd1;
								// Trace: design.sv:40926:17
								rf_we_raw = 1'b0;
								// Trace: design.sv:40927:17
								stall_multdiv = 1'b1;
							end
						branch_in_dec: begin
							// Trace: design.sv:40935:15
							id_fsm_d = (data_ind_timing_i || (!BranchTargetALU && branch_decision_i) ? 1'd1 : 1'd0);
							// Trace: design.sv:40937:15
							stall_branch = (~BranchTargetALU & branch_decision_i) | data_ind_timing_i;
							// Trace: design.sv:40938:15
							branch_set_raw_d = branch_decision_i | data_ind_timing_i;
							// Trace: design.sv:40940:15
							if (BranchPredictor)
								// Trace: design.sv:40941:17
								branch_not_set = ~branch_decision_i;
							// Trace: design.sv:40944:15
							perf_branch_o = 1'b1;
						end
						jump_in_dec: begin
							// Trace: design.sv:40949:15
							id_fsm_d = (BranchTargetALU ? 1'd0 : 1'd1);
							// Trace: design.sv:40950:15
							stall_jump = ~BranchTargetALU;
							// Trace: design.sv:40951:15
							jump_set_raw = jump_set_dec;
						end
						alu_multicycle_dec: begin
							// Trace: design.sv:40954:15
							stall_alu = 1'b1;
							// Trace: design.sv:40955:15
							id_fsm_d = 1'd1;
							// Trace: design.sv:40956:15
							rf_we_raw = 1'b0;
						end
						default:
							// Trace: design.sv:40959:15
							id_fsm_d = 1'd0;
					endcase
				1'd1: begin
					// Trace: design.sv:40965:11
					if (multdiv_en_dec)
						// Trace: design.sv:40966:13
						rf_we_raw = rf_we_dec & ex_valid_i;
					if (multicycle_done & ready_wb_i)
						// Trace: design.sv:40970:13
						id_fsm_d = 1'd0;
					else begin
						// Trace: design.sv:40972:13
						stall_multdiv = multdiv_en_dec;
						// Trace: design.sv:40973:13
						stall_branch = branch_in_dec;
						// Trace: design.sv:40974:13
						stall_jump = jump_in_dec;
					end
				end
				default:
					// Trace: design.sv:40979:11
					id_fsm_d = 1'd0;
			endcase
	end
	// Trace: design.sv:40986:3
	assign multdiv_ready_id_o = ready_wb_i;
	// Trace: design.sv:40993:3
	assign stall_id = ((((stall_ld_hz | stall_mem) | stall_multdiv) | stall_jump) | stall_branch) | stall_alu;
	// Trace: design.sv:41002:3
	assign instr_done = (~stall_id & ~flush_id) & instr_executing;
	// Trace: design.sv:41006:3
	assign instr_first_cycle = instr_valid_i & (id_fsm_q == 1'd0);
	// Trace: design.sv:41009:3
	assign instr_first_cycle_id_o = instr_first_cycle;
	// Trace: design.sv:41011:3
	generate
		if (WritebackStage) begin : gen_stall_mem
			// Trace: design.sv:41013:5
			wire rf_rd_a_wb_match;
			// Trace: design.sv:41014:5
			wire rf_rd_b_wb_match;
			// Trace: design.sv:41016:5
			wire rf_rd_a_hz;
			// Trace: design.sv:41017:5
			wire rf_rd_b_hz;
			// Trace: design.sv:41019:5
			wire outstanding_memory_access;
			// Trace: design.sv:41021:5
			wire instr_kill;
			// Trace: design.sv:41023:5
			assign multicycle_done = (lsu_req_dec ? ~stall_mem : ex_valid_i);
			// Trace: design.sv:41026:5
			assign outstanding_memory_access = (outstanding_load_wb_i | outstanding_store_wb_i) & ~lsu_resp_valid_i;
			// Trace: design.sv:41030:5
			assign data_req_allowed = ~outstanding_memory_access;
			// Trace: design.sv:41040:5
			assign instr_kill = ((instr_fetch_err_i | wb_exception) | id_exception) | ~controller_run;
			// Trace: design.sv:41061:5
			assign instr_executing_spec = ((instr_valid_i & ~instr_fetch_err_i) & controller_run) & ~stall_ld_hz;
			// Trace: design.sv:41066:5
			assign instr_executing = ((instr_valid_i & ~instr_kill) & ~stall_ld_hz) & ~outstanding_memory_access;
			// Trace: design.sv:41084:5
			assign stall_mem = instr_valid_i & (outstanding_memory_access | (lsu_req_dec & ~lsu_req_done_i));
			// Trace: design.sv:41092:5
			assign rf_rd_a_wb_match = (rf_waddr_wb_i == rf_raddr_a_o) & |rf_raddr_a_o;
			// Trace: design.sv:41093:5
			assign rf_rd_b_wb_match = (rf_waddr_wb_i == rf_raddr_b_o) & |rf_raddr_b_o;
			// Trace: design.sv:41095:5
			assign rf_rd_a_wb_match_o = rf_rd_a_wb_match;
			// Trace: design.sv:41096:5
			assign rf_rd_b_wb_match_o = rf_rd_b_wb_match;
			// Trace: design.sv:41100:5
			assign rf_rd_a_hz = rf_rd_a_wb_match & rf_ren_a;
			// Trace: design.sv:41101:5
			assign rf_rd_b_hz = rf_rd_b_wb_match & rf_ren_b;
			// Trace: design.sv:41106:5
			assign rf_rdata_a_fwd = (rf_rd_a_wb_match & rf_write_wb_i ? rf_wdata_fwd_wb_i : rf_rdata_a_i);
			// Trace: design.sv:41107:5
			assign rf_rdata_b_fwd = (rf_rd_b_wb_match & rf_write_wb_i ? rf_wdata_fwd_wb_i : rf_rdata_b_i);
			// Trace: design.sv:41109:5
			assign stall_ld_hz = outstanding_load_wb_i & (rf_rd_a_hz | rf_rd_b_hz);
			// Trace: design.sv:41111:5
			assign instr_type_wb_o = (~lsu_req_dec ? 2'd2 : (lsu_we ? 2'd1 : 2'd0));
			// Trace: design.sv:41115:5
			assign instr_id_done_o = en_wb_o & ready_wb_i;
			// Trace: design.sv:41118:5
			assign stall_wb = en_wb_o & ~ready_wb_i;
			// Trace: design.sv:41120:5
			assign perf_dside_wait_o = (instr_valid_i & ~instr_kill) & (outstanding_memory_access | stall_ld_hz);
		end
		else begin : gen_no_stall_mem
			// Trace: design.sv:41124:5
			assign multicycle_done = (lsu_req_dec ? lsu_resp_valid_i : ex_valid_i);
			// Trace: design.sv:41126:5
			assign data_req_allowed = instr_first_cycle;
			// Trace: design.sv:41130:5
			assign stall_mem = instr_valid_i & (lsu_req_dec & (~lsu_resp_valid_i | instr_first_cycle));
			// Trace: design.sv:41133:5
			assign stall_ld_hz = 1'b0;
			// Trace: design.sv:41136:5
			assign instr_executing_spec = (instr_valid_i & ~instr_fetch_err_i) & controller_run;
			// Trace: design.sv:41137:5
			assign instr_executing = instr_executing_spec;
			// Trace: design.sv:41144:5
			assign rf_rdata_a_fwd = rf_rdata_a_i;
			// Trace: design.sv:41145:5
			assign rf_rdata_b_fwd = rf_rdata_b_i;
			// Trace: design.sv:41147:5
			assign rf_rd_a_wb_match_o = 1'b0;
			// Trace: design.sv:41148:5
			assign rf_rd_b_wb_match_o = 1'b0;
			// Trace: design.sv:41153:5
			wire unused_data_req_done_ex;
			// Trace: design.sv:41154:5
			wire [4:0] unused_rf_waddr_wb;
			// Trace: design.sv:41155:5
			wire unused_rf_write_wb;
			// Trace: design.sv:41156:5
			wire unused_outstanding_load_wb;
			// Trace: design.sv:41157:5
			wire unused_outstanding_store_wb;
			// Trace: design.sv:41158:5
			wire unused_wb_exception;
			// Trace: design.sv:41159:5
			wire [31:0] unused_rf_wdata_fwd_wb;
			// Trace: design.sv:41160:5
			wire unused_id_exception;
			// Trace: design.sv:41162:5
			assign unused_data_req_done_ex = lsu_req_done_i;
			// Trace: design.sv:41163:5
			assign unused_rf_waddr_wb = rf_waddr_wb_i;
			// Trace: design.sv:41164:5
			assign unused_rf_write_wb = rf_write_wb_i;
			// Trace: design.sv:41165:5
			assign unused_outstanding_load_wb = outstanding_load_wb_i;
			// Trace: design.sv:41166:5
			assign unused_outstanding_store_wb = outstanding_store_wb_i;
			// Trace: design.sv:41167:5
			assign unused_wb_exception = wb_exception;
			// Trace: design.sv:41168:5
			assign unused_rf_wdata_fwd_wb = rf_wdata_fwd_wb_i;
			// Trace: design.sv:41169:5
			assign unused_id_exception = id_exception;
			// Trace: design.sv:41171:5
			assign instr_type_wb_o = 2'd2;
			// Trace: design.sv:41172:5
			assign stall_wb = 1'b0;
			// Trace: design.sv:41174:5
			assign perf_dside_wait_o = (instr_executing & lsu_req_dec) & ~lsu_resp_valid_i;
			// Trace: design.sv:41176:5
			assign instr_id_done_o = instr_done;
		end
	endgenerate
	// Trace: design.sv:41181:3
	assign instr_perf_count_id_o = (((~ebrk_insn & ~ecall_insn_dec) & ~illegal_insn_dec) & ~illegal_csr_insn_i) & ~instr_fetch_err_i;
	// Trace: design.sv:41186:3
	assign en_wb_o = instr_done;
	// Trace: design.sv:41188:3
	assign perf_mul_wait_o = stall_multdiv & mult_en_dec;
	// Trace: design.sv:41189:3
	assign perf_div_wait_o = stall_multdiv & div_en_dec;
	initial _sv2v_0 = 0;
endmodule
module ibex_if_stage (
	clk_i,
	rst_ni,
	boot_addr_i,
	req_i,
	instr_req_o,
	instr_addr_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_rdata_i,
	instr_err_i,
	ic_tag_req_o,
	ic_tag_write_o,
	ic_tag_addr_o,
	ic_tag_wdata_o,
	ic_tag_rdata_i,
	ic_data_req_o,
	ic_data_write_o,
	ic_data_addr_o,
	ic_data_wdata_o,
	ic_data_rdata_i,
	ic_scr_key_valid_i,
	instr_valid_id_o,
	instr_new_id_o,
	instr_rdata_id_o,
	instr_rdata_alu_id_o,
	instr_rdata_c_id_o,
	instr_is_compressed_id_o,
	instr_bp_taken_o,
	instr_fetch_err_o,
	instr_fetch_err_plus2_o,
	illegal_c_insn_id_o,
	dummy_instr_id_o,
	pc_if_o,
	pc_id_o,
	pmp_err_if_i,
	pmp_err_if_plus2_i,
	instr_valid_clear_i,
	pc_set_i,
	pc_mux_i,
	nt_branch_mispredict_i,
	nt_branch_addr_i,
	exc_pc_mux_i,
	exc_cause,
	dummy_instr_en_i,
	dummy_instr_mask_i,
	dummy_instr_seed_en_i,
	dummy_instr_seed_i,
	icache_enable_i,
	icache_inval_i,
	icache_ecc_error_o,
	branch_target_ex_i,
	csr_mepc_i,
	csr_depc_i,
	csr_mtvec_i,
	csr_mtvec_init_o,
	id_in_ready_i,
	pc_mismatch_alert_o,
	if_busy_o
);
	reg _sv2v_0;
	// removed import ibex_pkg::*;
	// Trace: design.sv:41269:13
	parameter [31:0] DmHaltAddr = 32'h1a110800;
	// Trace: design.sv:41270:13
	parameter [31:0] DmExceptionAddr = 32'h1a110808;
	// Trace: design.sv:41271:13
	parameter [0:0] DummyInstructions = 1'b0;
	// Trace: design.sv:41272:13
	parameter [0:0] ICache = 1'b0;
	// Trace: design.sv:41273:13
	parameter [0:0] ICacheECC = 1'b0;
	// Trace: design.sv:41274:13
	localparam [31:0] ibex_pkg_BUS_SIZE = 32;
	parameter [31:0] BusSizeECC = ibex_pkg_BUS_SIZE;
	// Trace: design.sv:41275:13
	localparam [31:0] ibex_pkg_ADDR_W = 32;
	localparam [31:0] ibex_pkg_IC_LINE_SIZE = 64;
	localparam [31:0] ibex_pkg_IC_LINE_BYTES = 8;
	localparam [31:0] ibex_pkg_IC_NUM_WAYS = 2;
	localparam [31:0] ibex_pkg_IC_SIZE_BYTES = 4096;
	localparam [31:0] ibex_pkg_IC_NUM_LINES = (ibex_pkg_IC_SIZE_BYTES / ibex_pkg_IC_NUM_WAYS) / ibex_pkg_IC_LINE_BYTES;
	localparam [31:0] ibex_pkg_IC_INDEX_W = $clog2(ibex_pkg_IC_NUM_LINES);
	localparam [31:0] ibex_pkg_IC_LINE_W = 3;
	localparam [31:0] ibex_pkg_IC_TAG_SIZE = ((ibex_pkg_ADDR_W - ibex_pkg_IC_INDEX_W) - ibex_pkg_IC_LINE_W) + 1;
	parameter [31:0] TagSizeECC = ibex_pkg_IC_TAG_SIZE;
	// Trace: design.sv:41276:13
	parameter [31:0] LineSizeECC = ibex_pkg_IC_LINE_SIZE;
	// Trace: design.sv:41277:13
	parameter [0:0] PCIncrCheck = 1'b0;
	// Trace: design.sv:41278:13
	parameter [0:0] ResetAll = 1'b0;
	// Trace: design.sv:41279:13
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	// removed localparam type ibex_pkg_lfsr_seed_t
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	// Trace: design.sv:41280:13
	// removed localparam type ibex_pkg_lfsr_perm_t
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	// Trace: design.sv:41281:13
	parameter [0:0] BranchPredictor = 1'b0;
	// Trace: design.sv:41283:3
	input wire clk_i;
	// Trace: design.sv:41284:3
	input wire rst_ni;
	// Trace: design.sv:41286:3
	input wire [31:0] boot_addr_i;
	// Trace: design.sv:41287:3
	input wire req_i;
	// Trace: design.sv:41290:3
	output wire instr_req_o;
	// Trace: design.sv:41291:3
	output wire [31:0] instr_addr_o;
	// Trace: design.sv:41292:3
	input wire instr_gnt_i;
	// Trace: design.sv:41293:3
	input wire instr_rvalid_i;
	// Trace: design.sv:41294:3
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:41295:3
	input wire instr_err_i;
	// Trace: design.sv:41298:3
	output wire [1:0] ic_tag_req_o;
	// Trace: design.sv:41299:3
	output wire ic_tag_write_o;
	// Trace: design.sv:41300:3
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr_o;
	// Trace: design.sv:41301:3
	output wire [TagSizeECC - 1:0] ic_tag_wdata_o;
	// Trace: design.sv:41302:3
	input wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata_i;
	// Trace: design.sv:41303:3
	output wire [1:0] ic_data_req_o;
	// Trace: design.sv:41304:3
	output wire ic_data_write_o;
	// Trace: design.sv:41305:3
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr_o;
	// Trace: design.sv:41306:3
	output wire [LineSizeECC - 1:0] ic_data_wdata_o;
	// Trace: design.sv:41307:3
	input wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata_i;
	// Trace: design.sv:41308:3
	input wire ic_scr_key_valid_i;
	// Trace: design.sv:41311:3
	output wire instr_valid_id_o;
	// Trace: design.sv:41312:3
	output wire instr_new_id_o;
	// Trace: design.sv:41313:3
	output reg [31:0] instr_rdata_id_o;
	// Trace: design.sv:41314:3
	output reg [31:0] instr_rdata_alu_id_o;
	// Trace: design.sv:41316:3
	output reg [15:0] instr_rdata_c_id_o;
	// Trace: design.sv:41319:3
	output reg instr_is_compressed_id_o;
	// Trace: design.sv:41321:3
	output wire instr_bp_taken_o;
	// Trace: design.sv:41323:3
	output reg instr_fetch_err_o;
	// Trace: design.sv:41324:3
	output reg instr_fetch_err_plus2_o;
	// Trace: design.sv:41325:3
	output reg illegal_c_insn_id_o;
	// Trace: design.sv:41327:3
	output reg dummy_instr_id_o;
	// Trace: design.sv:41328:3
	output wire [31:0] pc_if_o;
	// Trace: design.sv:41329:3
	output reg [31:0] pc_id_o;
	// Trace: design.sv:41330:3
	input wire pmp_err_if_i;
	// Trace: design.sv:41331:3
	input wire pmp_err_if_plus2_i;
	// Trace: design.sv:41334:3
	input wire instr_valid_clear_i;
	// Trace: design.sv:41335:3
	input wire pc_set_i;
	// Trace: design.sv:41336:3
	// removed localparam type ibex_pkg_pc_sel_e
	input wire [2:0] pc_mux_i;
	// Trace: design.sv:41337:3
	input wire nt_branch_mispredict_i;
	// Trace: design.sv:41339:3
	input wire [31:0] nt_branch_addr_i;
	// Trace: design.sv:41340:3
	// removed localparam type ibex_pkg_exc_pc_sel_e
	input wire [1:0] exc_pc_mux_i;
	// Trace: design.sv:41341:3
	// removed localparam type ibex_pkg_exc_cause_e
	input wire [5:0] exc_cause;
	// Trace: design.sv:41343:3
	input wire dummy_instr_en_i;
	// Trace: design.sv:41344:3
	input wire [2:0] dummy_instr_mask_i;
	// Trace: design.sv:41345:3
	input wire dummy_instr_seed_en_i;
	// Trace: design.sv:41346:3
	input wire [31:0] dummy_instr_seed_i;
	// Trace: design.sv:41347:3
	input wire icache_enable_i;
	// Trace: design.sv:41348:3
	input wire icache_inval_i;
	// Trace: design.sv:41349:3
	output wire icache_ecc_error_o;
	// Trace: design.sv:41352:3
	input wire [31:0] branch_target_ex_i;
	// Trace: design.sv:41355:3
	input wire [31:0] csr_mepc_i;
	// Trace: design.sv:41357:3
	input wire [31:0] csr_depc_i;
	// Trace: design.sv:41359:3
	input wire [31:0] csr_mtvec_i;
	// Trace: design.sv:41360:3
	output wire csr_mtvec_init_o;
	// Trace: design.sv:41363:3
	input wire id_in_ready_i;
	// Trace: design.sv:41366:3
	output wire pc_mismatch_alert_o;
	// Trace: design.sv:41367:3
	output wire if_busy_o;
	// Trace: design.sv:41370:3
	wire instr_valid_id_d;
	reg instr_valid_id_q;
	// Trace: design.sv:41371:3
	wire instr_new_id_d;
	reg instr_new_id_q;
	// Trace: design.sv:41374:3
	wire prefetch_busy;
	// Trace: design.sv:41375:3
	wire branch_req;
	// Trace: design.sv:41376:3
	reg [31:0] fetch_addr_n;
	// Trace: design.sv:41377:3
	wire unused_fetch_addr_n0;
	// Trace: design.sv:41379:3
	wire fetch_valid;
	// Trace: design.sv:41380:3
	wire fetch_ready;
	// Trace: design.sv:41381:3
	wire [31:0] fetch_rdata;
	// Trace: design.sv:41382:3
	wire [31:0] fetch_addr;
	// Trace: design.sv:41383:3
	wire fetch_err;
	// Trace: design.sv:41384:3
	wire fetch_err_plus2;
	// Trace: design.sv:41386:3
	wire [31:0] instr_decompressed;
	// Trace: design.sv:41387:3
	wire illegal_c_insn;
	// Trace: design.sv:41388:3
	wire instr_is_compressed;
	// Trace: design.sv:41390:3
	wire if_instr_valid;
	// Trace: design.sv:41391:3
	wire [31:0] if_instr_rdata;
	// Trace: design.sv:41392:3
	wire [31:0] if_instr_addr;
	// Trace: design.sv:41393:3
	wire if_instr_bus_err;
	// Trace: design.sv:41394:3
	wire if_instr_pmp_err;
	// Trace: design.sv:41395:3
	wire if_instr_err;
	// Trace: design.sv:41396:3
	wire if_instr_err_plus2;
	// Trace: design.sv:41398:3
	reg [31:0] exc_pc;
	// Trace: design.sv:41400:3
	wire [5:0] irq_id;
	// Trace: design.sv:41401:3
	wire unused_irq_bit;
	// Trace: design.sv:41403:3
	wire if_id_pipe_reg_we;
	// Trace: design.sv:41406:3
	wire stall_dummy_instr;
	// Trace: design.sv:41407:3
	wire [31:0] instr_out;
	// Trace: design.sv:41408:3
	wire instr_is_compressed_out;
	// Trace: design.sv:41409:3
	wire illegal_c_instr_out;
	// Trace: design.sv:41410:3
	wire instr_err_out;
	// Trace: design.sv:41412:3
	wire predict_branch_taken;
	// Trace: design.sv:41413:3
	wire [31:0] predict_branch_pc;
	// Trace: design.sv:41415:3
	wire [2:0] pc_mux_internal;
	// Trace: design.sv:41417:3
	wire [7:0] unused_boot_addr;
	// Trace: design.sv:41418:3
	wire [7:0] unused_csr_mtvec;
	// Trace: design.sv:41420:3
	assign unused_boot_addr = boot_addr_i[7:0];
	// Trace: design.sv:41421:3
	assign unused_csr_mtvec = csr_mtvec_i[7:0];
	// Trace: design.sv:41424:3
	assign irq_id = {exc_cause};
	// Trace: design.sv:41425:3
	assign unused_irq_bit = irq_id[5];
	// Trace: design.sv:41428:3
	always @(*) begin : exc_pc_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:41429:5
		(* full_case, parallel_case *)
		case (exc_pc_mux_i)
			2'd0:
				// Trace: design.sv:41430:23
				exc_pc = {csr_mtvec_i[31:8], 8'h00};
			2'd1:
				// Trace: design.sv:41431:23
				exc_pc = {csr_mtvec_i[31:8], 1'b0, irq_id[4:0], 2'b00};
			2'd2:
				// Trace: design.sv:41432:23
				exc_pc = DmHaltAddr;
			2'd3:
				// Trace: design.sv:41433:23
				exc_pc = DmExceptionAddr;
			default:
				// Trace: design.sv:41434:23
				exc_pc = {csr_mtvec_i[31:8], 8'h00};
		endcase
	end
	// Trace: design.sv:41440:3
	assign pc_mux_internal = ((BranchPredictor && predict_branch_taken) && !pc_set_i ? 3'd5 : pc_mux_i);
	// Trace: design.sv:41444:3
	always @(*) begin : fetch_addr_mux
		if (_sv2v_0)
			;
		// Trace: design.sv:41445:5
		(* full_case, parallel_case *)
		case (pc_mux_internal)
			3'd0:
				// Trace: design.sv:41446:16
				fetch_addr_n = {boot_addr_i[31:8], 8'h00};
			3'd1:
				// Trace: design.sv:41447:16
				fetch_addr_n = branch_target_ex_i;
			3'd2:
				// Trace: design.sv:41448:16
				fetch_addr_n = exc_pc;
			3'd3:
				// Trace: design.sv:41449:16
				fetch_addr_n = csr_mepc_i;
			3'd4:
				// Trace: design.sv:41450:16
				fetch_addr_n = csr_depc_i;
			3'd5:
				// Trace: design.sv:41453:16
				fetch_addr_n = (BranchPredictor ? predict_branch_pc : {boot_addr_i[31:8], 8'h00});
			default:
				// Trace: design.sv:41454:16
				fetch_addr_n = {boot_addr_i[31:8], 8'h00};
		endcase
	end
	// Trace: design.sv:41459:3
	assign csr_mtvec_init_o = (pc_mux_i == 3'd0) & pc_set_i;
	// Trace: design.sv:41461:3
	generate
		if (ICache) begin : gen_icache
			// Trace: design.sv:41463:5
			ibex_icache #(
				.ICacheECC(ICacheECC),
				.ResetAll(ResetAll),
				.BusSizeECC(BusSizeECC),
				.TagSizeECC(TagSizeECC),
				.LineSizeECC(LineSizeECC)
			) icache_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(req_i),
				.branch_i(branch_req),
				.branch_mispredict_i(nt_branch_mispredict_i),
				.mispredict_addr_i(nt_branch_addr_i),
				.addr_i({fetch_addr_n[31:1], 1'b0}),
				.ready_i(fetch_ready),
				.valid_o(fetch_valid),
				.rdata_o(fetch_rdata),
				.addr_o(fetch_addr),
				.err_o(fetch_err),
				.err_plus2_o(fetch_err_plus2),
				.instr_req_o(instr_req_o),
				.instr_addr_o(instr_addr_o),
				.instr_gnt_i(instr_gnt_i),
				.instr_rvalid_i(instr_rvalid_i),
				.instr_rdata_i(instr_rdata_i),
				.instr_err_i(instr_err_i),
				.ic_tag_req_o(ic_tag_req_o),
				.ic_tag_write_o(ic_tag_write_o),
				.ic_tag_addr_o(ic_tag_addr_o),
				.ic_tag_wdata_o(ic_tag_wdata_o),
				.ic_tag_rdata_i(ic_tag_rdata_i),
				.ic_data_req_o(ic_data_req_o),
				.ic_data_write_o(ic_data_write_o),
				.ic_data_addr_o(ic_data_addr_o),
				.ic_data_wdata_o(ic_data_wdata_o),
				.ic_data_rdata_i(ic_data_rdata_i),
				.ic_scr_key_valid_i(ic_scr_key_valid_i),
				.icache_enable_i(icache_enable_i),
				.icache_inval_i(icache_inval_i),
				.busy_o(prefetch_busy),
				.ecc_error_o(icache_ecc_error_o)
			);
		end
		else begin : gen_prefetch_buffer
			// Trace: design.sv:41513:5
			ibex_prefetch_buffer #(.ResetAll(ResetAll)) prefetch_buffer_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(req_i),
				.branch_i(branch_req),
				.branch_mispredict_i(nt_branch_mispredict_i),
				.mispredict_addr_i(nt_branch_addr_i),
				.addr_i({fetch_addr_n[31:1], 1'b0}),
				.ready_i(fetch_ready),
				.valid_o(fetch_valid),
				.rdata_o(fetch_rdata),
				.addr_o(fetch_addr),
				.err_o(fetch_err),
				.err_plus2_o(fetch_err_plus2),
				.instr_req_o(instr_req_o),
				.instr_addr_o(instr_addr_o),
				.instr_gnt_i(instr_gnt_i),
				.instr_rvalid_i(instr_rvalid_i),
				.instr_rdata_i(instr_rdata_i),
				.instr_err_i(instr_err_i),
				.busy_o(prefetch_busy)
			);
			// Trace: design.sv:41543:5
			wire unused_icen;
			wire unused_icinv;
			wire unused_scr_key_valid;
			// Trace: design.sv:41544:5
			wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] unused_tag_ram_input;
			// Trace: design.sv:41545:5
			wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] unused_data_ram_input;
			// Trace: design.sv:41546:5
			assign unused_icen = icache_enable_i;
			// Trace: design.sv:41547:5
			assign unused_icinv = icache_inval_i;
			// Trace: design.sv:41548:5
			assign unused_tag_ram_input = ic_tag_rdata_i;
			// Trace: design.sv:41549:5
			assign unused_data_ram_input = ic_data_rdata_i;
			// Trace: design.sv:41550:5
			assign unused_scr_key_valid = ic_scr_key_valid_i;
			// Trace: design.sv:41551:5
			assign ic_tag_req_o = 'b0;
			// Trace: design.sv:41552:5
			assign ic_tag_write_o = 'b0;
			// Trace: design.sv:41553:5
			assign ic_tag_addr_o = 'b0;
			// Trace: design.sv:41554:5
			assign ic_tag_wdata_o = 'b0;
			// Trace: design.sv:41555:5
			assign ic_data_req_o = 'b0;
			// Trace: design.sv:41556:5
			assign ic_data_write_o = 'b0;
			// Trace: design.sv:41557:5
			assign ic_data_addr_o = 'b0;
			// Trace: design.sv:41558:5
			assign ic_data_wdata_o = 'b0;
			// Trace: design.sv:41559:5
			assign icache_ecc_error_o = 'b0;
		end
	endgenerate
	// Trace: design.sv:41578:3
	assign unused_fetch_addr_n0 = fetch_addr_n[0];
	// Trace: design.sv:41580:3
	assign branch_req = pc_set_i | predict_branch_taken;
	// Trace: design.sv:41582:3
	assign pc_if_o = if_instr_addr;
	// Trace: design.sv:41583:3
	assign if_busy_o = prefetch_busy;
	// Trace: design.sv:41588:3
	assign if_instr_pmp_err = pmp_err_if_i | ((if_instr_addr[2] & ~instr_is_compressed) & pmp_err_if_plus2_i);
	// Trace: design.sv:41592:3
	assign if_instr_err = if_instr_bus_err | if_instr_pmp_err;
	// Trace: design.sv:41595:3
	assign if_instr_err_plus2 = (((if_instr_addr[2] & ~instr_is_compressed) & pmp_err_if_plus2_i) | fetch_err_plus2) & ~pmp_err_if_i;
	// Trace: design.sv:41603:3
	ibex_compressed_decoder compressed_decoder_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.valid_i(fetch_valid & ~fetch_err),
		.instr_i(if_instr_rdata),
		.instr_o(instr_decompressed),
		.is_compressed_o(instr_is_compressed),
		.illegal_instr_o(illegal_c_insn)
	);
	// Trace: design.sv:41614:3
	generate
		if (DummyInstructions) begin : gen_dummy_instr
			// Trace: design.sv:41616:5
			wire insert_dummy_instr;
			// Trace: design.sv:41617:5
			wire [31:0] dummy_instr_data;
			// Trace: design.sv:41619:5
			ibex_dummy_instr #(
				.RndCnstLfsrSeed(RndCnstLfsrSeed),
				.RndCnstLfsrPerm(RndCnstLfsrPerm)
			) dummy_instr_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.dummy_instr_en_i(dummy_instr_en_i),
				.dummy_instr_mask_i(dummy_instr_mask_i),
				.dummy_instr_seed_en_i(dummy_instr_seed_en_i),
				.dummy_instr_seed_i(dummy_instr_seed_i),
				.fetch_valid_i(fetch_valid),
				.id_in_ready_i(id_in_ready_i),
				.insert_dummy_instr_o(insert_dummy_instr),
				.dummy_instr_data_o(dummy_instr_data)
			);
			// Trace: design.sv:41636:5
			assign instr_out = (insert_dummy_instr ? dummy_instr_data : instr_decompressed);
			// Trace: design.sv:41637:5
			assign instr_is_compressed_out = (insert_dummy_instr ? 1'b0 : instr_is_compressed);
			// Trace: design.sv:41638:5
			assign illegal_c_instr_out = (insert_dummy_instr ? 1'b0 : illegal_c_insn);
			// Trace: design.sv:41639:5
			assign instr_err_out = (insert_dummy_instr ? 1'b0 : if_instr_err);
			// Trace: design.sv:41644:5
			assign stall_dummy_instr = insert_dummy_instr;
			// Trace: design.sv:41647:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:41648:7
				if (!rst_ni)
					// Trace: design.sv:41649:9
					dummy_instr_id_o <= 1'b0;
				else if (if_id_pipe_reg_we)
					// Trace: design.sv:41651:9
					dummy_instr_id_o <= insert_dummy_instr;
		end
		else begin : gen_no_dummy_instr
			// Trace: design.sv:41656:5
			wire unused_dummy_en;
			// Trace: design.sv:41657:5
			wire [2:0] unused_dummy_mask;
			// Trace: design.sv:41658:5
			wire unused_dummy_seed_en;
			// Trace: design.sv:41659:5
			wire [31:0] unused_dummy_seed;
			// Trace: design.sv:41661:5
			assign unused_dummy_en = dummy_instr_en_i;
			// Trace: design.sv:41662:5
			assign unused_dummy_mask = dummy_instr_mask_i;
			// Trace: design.sv:41663:5
			assign unused_dummy_seed_en = dummy_instr_seed_en_i;
			// Trace: design.sv:41664:5
			assign unused_dummy_seed = dummy_instr_seed_i;
			// Trace: design.sv:41665:5
			assign instr_out = instr_decompressed;
			// Trace: design.sv:41666:5
			assign instr_is_compressed_out = instr_is_compressed;
			// Trace: design.sv:41667:5
			assign illegal_c_instr_out = illegal_c_insn;
			// Trace: design.sv:41668:5
			assign instr_err_out = if_instr_err;
			// Trace: design.sv:41669:5
			assign stall_dummy_instr = 1'b0;
			// Trace: design.sv:41670:5
			wire [1:1] sv2v_tmp_C8A0C;
			assign sv2v_tmp_C8A0C = 1'b0;
			always @(*) dummy_instr_id_o = sv2v_tmp_C8A0C;
		end
	endgenerate
	// Trace: design.sv:41676:3
	assign instr_valid_id_d = ((if_instr_valid & id_in_ready_i) & ~pc_set_i) | (instr_valid_id_q & ~instr_valid_clear_i);
	// Trace: design.sv:41678:3
	assign instr_new_id_d = if_instr_valid & id_in_ready_i;
	// Trace: design.sv:41680:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:41681:5
		if (!rst_ni) begin
			// Trace: design.sv:41682:7
			instr_valid_id_q <= 1'b0;
			// Trace: design.sv:41683:7
			instr_new_id_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:41685:7
			instr_valid_id_q <= instr_valid_id_d;
			// Trace: design.sv:41686:7
			instr_new_id_q <= instr_new_id_d;
		end
	// Trace: design.sv:41690:3
	assign instr_valid_id_o = instr_valid_id_q;
	// Trace: design.sv:41692:3
	assign instr_new_id_o = instr_new_id_q;
	// Trace: design.sv:41695:3
	assign if_id_pipe_reg_we = instr_new_id_d;
	// Trace: design.sv:41697:3
	generate
		if (ResetAll) begin : g_instr_rdata_ra
			// Trace: design.sv:41698:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:41699:7
				if (!rst_ni) begin
					// Trace: design.sv:41700:9
					instr_rdata_id_o <= 1'sb0;
					// Trace: design.sv:41701:9
					instr_rdata_alu_id_o <= 1'sb0;
					// Trace: design.sv:41702:9
					instr_fetch_err_o <= 1'sb0;
					// Trace: design.sv:41703:9
					instr_fetch_err_plus2_o <= 1'sb0;
					// Trace: design.sv:41704:9
					instr_rdata_c_id_o <= 1'sb0;
					// Trace: design.sv:41705:9
					instr_is_compressed_id_o <= 1'sb0;
					// Trace: design.sv:41706:9
					illegal_c_insn_id_o <= 1'sb0;
					// Trace: design.sv:41707:9
					pc_id_o <= 1'sb0;
				end
				else if (if_id_pipe_reg_we) begin
					// Trace: design.sv:41709:9
					instr_rdata_id_o <= instr_out;
					// Trace: design.sv:41711:9
					instr_rdata_alu_id_o <= instr_out;
					// Trace: design.sv:41712:9
					instr_fetch_err_o <= instr_err_out;
					// Trace: design.sv:41713:9
					instr_fetch_err_plus2_o <= if_instr_err_plus2;
					// Trace: design.sv:41714:9
					instr_rdata_c_id_o <= if_instr_rdata[15:0];
					// Trace: design.sv:41715:9
					instr_is_compressed_id_o <= instr_is_compressed_out;
					// Trace: design.sv:41716:9
					illegal_c_insn_id_o <= illegal_c_instr_out;
					// Trace: design.sv:41717:9
					pc_id_o <= pc_if_o;
				end
		end
		else begin : g_instr_rdata_nr
			// Trace: design.sv:41721:5
			always @(posedge clk_i)
				// Trace: design.sv:41722:7
				if (if_id_pipe_reg_we) begin
					// Trace: design.sv:41723:9
					instr_rdata_id_o <= instr_out;
					// Trace: design.sv:41725:9
					instr_rdata_alu_id_o <= instr_out;
					// Trace: design.sv:41726:9
					instr_fetch_err_o <= instr_err_out;
					// Trace: design.sv:41727:9
					instr_fetch_err_plus2_o <= if_instr_err_plus2;
					// Trace: design.sv:41728:9
					instr_rdata_c_id_o <= if_instr_rdata[15:0];
					// Trace: design.sv:41729:9
					instr_is_compressed_id_o <= instr_is_compressed_out;
					// Trace: design.sv:41730:9
					illegal_c_insn_id_o <= illegal_c_instr_out;
					// Trace: design.sv:41731:9
					pc_id_o <= pc_if_o;
				end
		end
	endgenerate
	// Trace: design.sv:41737:3
	generate
		if (PCIncrCheck) begin : g_secure_pc
			// Trace: design.sv:41739:5
			wire [31:0] prev_instr_addr_incr;
			wire [31:0] prev_instr_addr_incr_buf;
			// Trace: design.sv:41740:5
			reg prev_instr_seq_q;
			wire prev_instr_seq_d;
			// Trace: design.sv:41744:5
			assign prev_instr_seq_d = (((prev_instr_seq_q | instr_new_id_d) & ~branch_req) & ~if_instr_err) & ~stall_dummy_instr;
			// Trace: design.sv:41747:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:41748:7
				if (!rst_ni)
					// Trace: design.sv:41749:9
					prev_instr_seq_q <= 1'b0;
				else
					// Trace: design.sv:41751:9
					prev_instr_seq_q <= prev_instr_seq_d;
			// Trace: design.sv:41755:5
			assign prev_instr_addr_incr = pc_id_o + (instr_is_compressed_id_o ? 32'd2 : 32'd4);
			// Trace: design.sv:41758:5
			prim_buf #(.Width(32)) u_prev_instr_addr_incr_buf(
				.in_i(prev_instr_addr_incr),
				.out_o(prev_instr_addr_incr_buf)
			);
			// Trace: design.sv:41764:5
			assign pc_mismatch_alert_o = prev_instr_seq_q & (pc_if_o != prev_instr_addr_incr_buf);
		end
		else begin : g_no_secure_pc
			// Trace: design.sv:41767:5
			assign pc_mismatch_alert_o = 1'b0;
		end
	endgenerate
	// Trace: design.sv:41770:3
	generate
		if (BranchPredictor) begin : g_branch_predictor
			// Trace: design.sv:41771:5
			reg [31:0] instr_skid_data_q;
			// Trace: design.sv:41772:5
			reg [31:0] instr_skid_addr_q;
			// Trace: design.sv:41773:5
			reg instr_skid_bp_taken_q;
			// Trace: design.sv:41774:5
			reg instr_skid_valid_q;
			wire instr_skid_valid_d;
			// Trace: design.sv:41775:5
			wire instr_skid_en;
			// Trace: design.sv:41776:5
			reg instr_bp_taken_q;
			wire instr_bp_taken_d;
			// Trace: design.sv:41778:5
			wire predict_branch_taken_raw;
			if (ResetAll) begin : g_bp_taken_ra
				// Trace: design.sv:41782:7
				always @(posedge clk_i or negedge rst_ni)
					// Trace: design.sv:41783:9
					if (!rst_ni)
						// Trace: design.sv:41784:11
						instr_bp_taken_q <= 1'sb0;
					else if (if_id_pipe_reg_we)
						// Trace: design.sv:41786:11
						instr_bp_taken_q <= instr_bp_taken_d;
			end
			else begin : g_bp_taken_nr
				// Trace: design.sv:41790:7
				always @(posedge clk_i)
					// Trace: design.sv:41791:9
					if (if_id_pipe_reg_we)
						// Trace: design.sv:41792:11
						instr_bp_taken_q <= instr_bp_taken_d;
			end
			// Trace: design.sv:41805:5
			assign instr_skid_en = ((predict_branch_taken & ~pc_set_i) & ~id_in_ready_i) & ~instr_skid_valid_q;
			// Trace: design.sv:41807:5
			assign instr_skid_valid_d = ((instr_skid_valid_q & ~id_in_ready_i) & ~stall_dummy_instr) | instr_skid_en;
			// Trace: design.sv:41810:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:41811:7
				if (!rst_ni)
					// Trace: design.sv:41812:9
					instr_skid_valid_q <= 1'b0;
				else
					// Trace: design.sv:41814:9
					instr_skid_valid_q <= instr_skid_valid_d;
			if (ResetAll) begin : g_instr_skid_ra
				// Trace: design.sv:41819:7
				always @(posedge clk_i or negedge rst_ni)
					// Trace: design.sv:41820:9
					if (!rst_ni) begin
						// Trace: design.sv:41821:11
						instr_skid_bp_taken_q <= 1'sb0;
						// Trace: design.sv:41822:11
						instr_skid_data_q <= 1'sb0;
						// Trace: design.sv:41823:11
						instr_skid_addr_q <= 1'sb0;
					end
					else if (instr_skid_en) begin
						// Trace: design.sv:41825:11
						instr_skid_bp_taken_q <= predict_branch_taken;
						// Trace: design.sv:41826:11
						instr_skid_data_q <= fetch_rdata;
						// Trace: design.sv:41827:11
						instr_skid_addr_q <= fetch_addr;
					end
			end
			else begin : g_instr_skid_nr
				// Trace: design.sv:41831:7
				always @(posedge clk_i)
					// Trace: design.sv:41832:9
					if (instr_skid_en) begin
						// Trace: design.sv:41833:11
						instr_skid_bp_taken_q <= predict_branch_taken;
						// Trace: design.sv:41834:11
						instr_skid_data_q <= fetch_rdata;
						// Trace: design.sv:41835:11
						instr_skid_addr_q <= fetch_addr;
					end
			end
			// Trace: design.sv:41840:5
			ibex_branch_predict branch_predict_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.fetch_rdata_i(fetch_rdata),
				.fetch_pc_i(fetch_addr),
				.fetch_valid_i(fetch_valid),
				.predict_branch_taken_o(predict_branch_taken_raw),
				.predict_branch_pc_o(predict_branch_pc)
			);
			// Trace: design.sv:41855:5
			assign predict_branch_taken = (predict_branch_taken_raw & ~instr_skid_valid_q) & ~fetch_err;
			// Trace: design.sv:41857:5
			assign if_instr_valid = fetch_valid | (instr_skid_valid_q & ~nt_branch_mispredict_i);
			// Trace: design.sv:41858:5
			assign if_instr_rdata = (instr_skid_valid_q ? instr_skid_data_q : fetch_rdata);
			// Trace: design.sv:41859:5
			assign if_instr_addr = (instr_skid_valid_q ? instr_skid_addr_q : fetch_addr);
			// Trace: design.sv:41863:5
			assign if_instr_bus_err = ~instr_skid_valid_q & fetch_err;
			// Trace: design.sv:41864:5
			assign instr_bp_taken_d = (instr_skid_valid_q ? instr_skid_bp_taken_q : predict_branch_taken);
			// Trace: design.sv:41866:5
			assign fetch_ready = (id_in_ready_i & ~stall_dummy_instr) & ~instr_skid_valid_q;
			// Trace: design.sv:41868:5
			assign instr_bp_taken_o = instr_bp_taken_q;
		end
		else begin : g_no_branch_predictor
			// Trace: design.sv:41873:5
			assign instr_bp_taken_o = 1'b0;
			// Trace: design.sv:41874:5
			assign predict_branch_taken = 1'b0;
			// Trace: design.sv:41875:5
			assign predict_branch_pc = 32'b00000000000000000000000000000000;
			// Trace: design.sv:41877:5
			assign if_instr_valid = fetch_valid;
			// Trace: design.sv:41878:5
			assign if_instr_rdata = fetch_rdata;
			// Trace: design.sv:41879:5
			assign if_instr_addr = fetch_addr;
			// Trace: design.sv:41880:5
			assign if_instr_bus_err = fetch_err;
			// Trace: design.sv:41881:5
			assign fetch_ready = id_in_ready_i & ~stall_dummy_instr;
		end
	endgenerate
	// Trace: design.sv:41891:3
	initial _sv2v_0 = 0;
endmodule
module ibex_load_store_unit (
	clk_i,
	rst_ni,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_err_i,
	data_pmp_err_i,
	data_addr_o,
	data_we_o,
	data_be_o,
	data_wdata_o,
	data_rdata_i,
	lsu_we_i,
	lsu_type_i,
	lsu_wdata_i,
	lsu_sign_ext_i,
	lsu_rdata_o,
	lsu_rdata_valid_o,
	lsu_req_i,
	adder_result_ex_i,
	addr_incr_req_o,
	addr_last_o,
	lsu_req_done_o,
	lsu_resp_valid_o,
	load_err_o,
	store_err_o,
	busy_o,
	perf_load_o,
	perf_store_o
);
	reg _sv2v_0;
	// Trace: design.sv:42022:3
	input wire clk_i;
	// Trace: design.sv:42023:3
	input wire rst_ni;
	// Trace: design.sv:42026:3
	output reg data_req_o;
	// Trace: design.sv:42027:3
	input wire data_gnt_i;
	// Trace: design.sv:42028:3
	input wire data_rvalid_i;
	// Trace: design.sv:42029:3
	input wire data_err_i;
	// Trace: design.sv:42030:3
	input wire data_pmp_err_i;
	// Trace: design.sv:42032:3
	output wire [31:0] data_addr_o;
	// Trace: design.sv:42033:3
	output wire data_we_o;
	// Trace: design.sv:42034:3
	output wire [3:0] data_be_o;
	// Trace: design.sv:42035:3
	output wire [31:0] data_wdata_o;
	// Trace: design.sv:42036:3
	input wire [31:0] data_rdata_i;
	// Trace: design.sv:42039:3
	input wire lsu_we_i;
	// Trace: design.sv:42040:3
	input wire [1:0] lsu_type_i;
	// Trace: design.sv:42041:3
	input wire [31:0] lsu_wdata_i;
	// Trace: design.sv:42042:3
	input wire lsu_sign_ext_i;
	// Trace: design.sv:42044:3
	output wire [31:0] lsu_rdata_o;
	// Trace: design.sv:42045:3
	output wire lsu_rdata_valid_o;
	// Trace: design.sv:42046:3
	input wire lsu_req_i;
	// Trace: design.sv:42048:3
	input wire [31:0] adder_result_ex_i;
	// Trace: design.sv:42050:3
	output reg addr_incr_req_o;
	// Trace: design.sv:42052:3
	output wire [31:0] addr_last_o;
	// Trace: design.sv:42056:3
	output wire lsu_req_done_o;
	// Trace: design.sv:42060:3
	output wire lsu_resp_valid_o;
	// Trace: design.sv:42063:3
	output wire load_err_o;
	// Trace: design.sv:42064:3
	output wire store_err_o;
	// Trace: design.sv:42066:3
	output wire busy_o;
	// Trace: design.sv:42068:3
	output reg perf_load_o;
	// Trace: design.sv:42069:3
	output reg perf_store_o;
	// Trace: design.sv:42072:3
	wire [31:0] data_addr;
	// Trace: design.sv:42073:3
	wire [31:0] data_addr_w_aligned;
	// Trace: design.sv:42074:3
	reg [31:0] addr_last_q;
	wire [31:0] addr_last_d;
	// Trace: design.sv:42076:3
	reg addr_update;
	// Trace: design.sv:42077:3
	reg ctrl_update;
	// Trace: design.sv:42078:3
	reg rdata_update;
	// Trace: design.sv:42079:3
	reg [31:8] rdata_q;
	// Trace: design.sv:42080:3
	reg [1:0] rdata_offset_q;
	// Trace: design.sv:42081:3
	reg [1:0] data_type_q;
	// Trace: design.sv:42082:3
	reg data_sign_ext_q;
	// Trace: design.sv:42083:3
	reg data_we_q;
	// Trace: design.sv:42085:3
	wire [1:0] data_offset;
	// Trace: design.sv:42087:3
	reg [3:0] data_be;
	// Trace: design.sv:42088:3
	reg [31:0] data_wdata;
	// Trace: design.sv:42090:3
	reg [31:0] data_rdata_ext;
	// Trace: design.sv:42092:3
	reg [31:0] rdata_w_ext;
	// Trace: design.sv:42093:3
	reg [31:0] rdata_h_ext;
	// Trace: design.sv:42094:3
	reg [31:0] rdata_b_ext;
	// Trace: design.sv:42096:3
	wire split_misaligned_access;
	// Trace: design.sv:42097:3
	reg handle_misaligned_q;
	reg handle_misaligned_d;
	// Trace: design.sv:42099:3
	reg pmp_err_q;
	reg pmp_err_d;
	// Trace: design.sv:42100:3
	reg lsu_err_q;
	reg lsu_err_d;
	// Trace: design.sv:42101:3
	wire data_or_pmp_err;
	// Trace: design.sv:42103:3
	// removed localparam type ls_fsm_e
	// Trace: design.sv:42108:3
	reg [2:0] ls_fsm_cs;
	reg [2:0] ls_fsm_ns;
	// Trace: design.sv:42110:3
	assign data_addr = adder_result_ex_i;
	// Trace: design.sv:42111:3
	assign data_offset = data_addr[1:0];
	// Trace: design.sv:42117:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42118:5
		(* full_case, parallel_case *)
		case (lsu_type_i)
			2'b00:
				// Trace: design.sv:42120:9
				if (!handle_misaligned_q)
					// Trace: design.sv:42121:11
					(* full_case, parallel_case *)
					case (data_offset)
						2'b00:
							// Trace: design.sv:42122:22
							data_be = 4'b1111;
						2'b01:
							// Trace: design.sv:42123:22
							data_be = 4'b1110;
						2'b10:
							// Trace: design.sv:42124:22
							data_be = 4'b1100;
						2'b11:
							// Trace: design.sv:42125:22
							data_be = 4'b1000;
						default:
							// Trace: design.sv:42126:22
							data_be = 4'b1111;
					endcase
				else
					// Trace: design.sv:42129:11
					(* full_case, parallel_case *)
					case (data_offset)
						2'b00:
							// Trace: design.sv:42130:22
							data_be = 4'b0000;
						2'b01:
							// Trace: design.sv:42131:22
							data_be = 4'b0001;
						2'b10:
							// Trace: design.sv:42132:22
							data_be = 4'b0011;
						2'b11:
							// Trace: design.sv:42133:22
							data_be = 4'b0111;
						default:
							// Trace: design.sv:42134:22
							data_be = 4'b1111;
					endcase
			2'b01:
				// Trace: design.sv:42140:9
				if (!handle_misaligned_q)
					// Trace: design.sv:42141:11
					(* full_case, parallel_case *)
					case (data_offset)
						2'b00:
							// Trace: design.sv:42142:22
							data_be = 4'b0011;
						2'b01:
							// Trace: design.sv:42143:22
							data_be = 4'b0110;
						2'b10:
							// Trace: design.sv:42144:22
							data_be = 4'b1100;
						2'b11:
							// Trace: design.sv:42145:22
							data_be = 4'b1000;
						default:
							// Trace: design.sv:42146:22
							data_be = 4'b1111;
					endcase
				else
					// Trace: design.sv:42149:11
					data_be = 4'b0001;
			2'b10, 2'b11:
				// Trace: design.sv:42155:9
				(* full_case, parallel_case *)
				case (data_offset)
					2'b00:
						// Trace: design.sv:42156:20
						data_be = 4'b0001;
					2'b01:
						// Trace: design.sv:42157:20
						data_be = 4'b0010;
					2'b10:
						// Trace: design.sv:42158:20
						data_be = 4'b0100;
					2'b11:
						// Trace: design.sv:42159:20
						data_be = 4'b1000;
					default:
						// Trace: design.sv:42160:20
						data_be = 4'b1111;
				endcase
			default:
				// Trace: design.sv:42164:20
				data_be = 4'b1111;
		endcase
	end
	// Trace: design.sv:42174:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42175:5
		(* full_case, parallel_case *)
		case (data_offset)
			2'b00:
				// Trace: design.sv:42176:16
				data_wdata = lsu_wdata_i[31:0];
			2'b01:
				// Trace: design.sv:42177:16
				data_wdata = {lsu_wdata_i[23:0], lsu_wdata_i[31:24]};
			2'b10:
				// Trace: design.sv:42178:16
				data_wdata = {lsu_wdata_i[15:0], lsu_wdata_i[31:16]};
			2'b11:
				// Trace: design.sv:42179:16
				data_wdata = {lsu_wdata_i[7:0], lsu_wdata_i[31:8]};
			default:
				// Trace: design.sv:42180:16
				data_wdata = lsu_wdata_i[31:0];
		endcase
	end
	// Trace: design.sv:42189:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:42190:5
		if (!rst_ni)
			// Trace: design.sv:42191:7
			rdata_q <= 1'sb0;
		else if (rdata_update)
			// Trace: design.sv:42193:7
			rdata_q <= data_rdata_i[31:8];
	// Trace: design.sv:42198:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:42199:5
		if (!rst_ni) begin
			// Trace: design.sv:42200:7
			rdata_offset_q <= 2'h0;
			// Trace: design.sv:42201:7
			data_type_q <= 2'h0;
			// Trace: design.sv:42202:7
			data_sign_ext_q <= 1'b0;
			// Trace: design.sv:42203:7
			data_we_q <= 1'b0;
		end
		else if (ctrl_update) begin
			// Trace: design.sv:42205:7
			rdata_offset_q <= data_offset;
			// Trace: design.sv:42206:7
			data_type_q <= lsu_type_i;
			// Trace: design.sv:42207:7
			data_sign_ext_q <= lsu_sign_ext_i;
			// Trace: design.sv:42208:7
			data_we_q <= lsu_we_i;
		end
	// Trace: design.sv:42216:3
	assign addr_last_d = (addr_incr_req_o ? data_addr_w_aligned : data_addr);
	// Trace: design.sv:42218:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:42219:5
		if (!rst_ni)
			// Trace: design.sv:42220:7
			addr_last_q <= 1'sb0;
		else if (addr_update)
			// Trace: design.sv:42222:7
			addr_last_q <= addr_last_d;
	// Trace: design.sv:42227:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42228:5
		(* full_case, parallel_case *)
		case (rdata_offset_q)
			2'b00:
				// Trace: design.sv:42229:16
				rdata_w_ext = data_rdata_i[31:0];
			2'b01:
				// Trace: design.sv:42230:16
				rdata_w_ext = {data_rdata_i[7:0], rdata_q[31:8]};
			2'b10:
				// Trace: design.sv:42231:16
				rdata_w_ext = {data_rdata_i[15:0], rdata_q[31:16]};
			2'b11:
				// Trace: design.sv:42232:16
				rdata_w_ext = {data_rdata_i[23:0], rdata_q[31:24]};
			default:
				// Trace: design.sv:42233:16
				rdata_w_ext = data_rdata_i[31:0];
		endcase
	end
	// Trace: design.sv:42242:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42243:5
		(* full_case, parallel_case *)
		case (rdata_offset_q)
			2'b00:
				// Trace: design.sv:42245:9
				if (!data_sign_ext_q)
					// Trace: design.sv:42246:11
					rdata_h_ext = {16'h0000, data_rdata_i[15:0]};
				else
					// Trace: design.sv:42248:11
					rdata_h_ext = {{16 {data_rdata_i[15]}}, data_rdata_i[15:0]};
			2'b01:
				// Trace: design.sv:42253:9
				if (!data_sign_ext_q)
					// Trace: design.sv:42254:11
					rdata_h_ext = {16'h0000, data_rdata_i[23:8]};
				else
					// Trace: design.sv:42256:11
					rdata_h_ext = {{16 {data_rdata_i[23]}}, data_rdata_i[23:8]};
			2'b10:
				// Trace: design.sv:42261:9
				if (!data_sign_ext_q)
					// Trace: design.sv:42262:11
					rdata_h_ext = {16'h0000, data_rdata_i[31:16]};
				else
					// Trace: design.sv:42264:11
					rdata_h_ext = {{16 {data_rdata_i[31]}}, data_rdata_i[31:16]};
			2'b11:
				// Trace: design.sv:42269:9
				if (!data_sign_ext_q)
					// Trace: design.sv:42270:11
					rdata_h_ext = {16'h0000, data_rdata_i[7:0], rdata_q[31:24]};
				else
					// Trace: design.sv:42272:11
					rdata_h_ext = {{16 {data_rdata_i[7]}}, data_rdata_i[7:0], rdata_q[31:24]};
			default:
				// Trace: design.sv:42276:16
				rdata_h_ext = {16'h0000, data_rdata_i[15:0]};
		endcase
	end
	// Trace: design.sv:42281:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42282:5
		(* full_case, parallel_case *)
		case (rdata_offset_q)
			2'b00:
				// Trace: design.sv:42284:9
				if (!data_sign_ext_q)
					// Trace: design.sv:42285:11
					rdata_b_ext = {24'h000000, data_rdata_i[7:0]};
				else
					// Trace: design.sv:42287:11
					rdata_b_ext = {{24 {data_rdata_i[7]}}, data_rdata_i[7:0]};
			2'b01:
				// Trace: design.sv:42292:9
				if (!data_sign_ext_q)
					// Trace: design.sv:42293:11
					rdata_b_ext = {24'h000000, data_rdata_i[15:8]};
				else
					// Trace: design.sv:42295:11
					rdata_b_ext = {{24 {data_rdata_i[15]}}, data_rdata_i[15:8]};
			2'b10:
				// Trace: design.sv:42300:9
				if (!data_sign_ext_q)
					// Trace: design.sv:42301:11
					rdata_b_ext = {24'h000000, data_rdata_i[23:16]};
				else
					// Trace: design.sv:42303:11
					rdata_b_ext = {{24 {data_rdata_i[23]}}, data_rdata_i[23:16]};
			2'b11:
				// Trace: design.sv:42308:9
				if (!data_sign_ext_q)
					// Trace: design.sv:42309:11
					rdata_b_ext = {24'h000000, data_rdata_i[31:24]};
				else
					// Trace: design.sv:42311:11
					rdata_b_ext = {{24 {data_rdata_i[31]}}, data_rdata_i[31:24]};
			default:
				// Trace: design.sv:42315:16
				rdata_b_ext = {24'h000000, data_rdata_i[7:0]};
		endcase
	end
	// Trace: design.sv:42320:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42321:5
		(* full_case, parallel_case *)
		case (data_type_q)
			2'b00:
				// Trace: design.sv:42322:20
				data_rdata_ext = rdata_w_ext;
			2'b01:
				// Trace: design.sv:42323:20
				data_rdata_ext = rdata_h_ext;
			2'b10, 2'b11:
				// Trace: design.sv:42324:20
				data_rdata_ext = rdata_b_ext;
			default:
				// Trace: design.sv:42325:20
				data_rdata_ext = rdata_w_ext;
		endcase
	end
	// Trace: design.sv:42334:3
	assign split_misaligned_access = ((lsu_type_i == 2'b00) && (data_offset != 2'b00)) || ((lsu_type_i == 2'b01) && (data_offset == 2'b11));
	// Trace: design.sv:42339:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42340:5
		ls_fsm_ns = ls_fsm_cs;
		// Trace: design.sv:42342:5
		data_req_o = 1'b0;
		// Trace: design.sv:42343:5
		addr_incr_req_o = 1'b0;
		// Trace: design.sv:42344:5
		handle_misaligned_d = handle_misaligned_q;
		// Trace: design.sv:42345:5
		pmp_err_d = pmp_err_q;
		// Trace: design.sv:42346:5
		lsu_err_d = lsu_err_q;
		// Trace: design.sv:42348:5
		addr_update = 1'b0;
		// Trace: design.sv:42349:5
		ctrl_update = 1'b0;
		// Trace: design.sv:42350:5
		rdata_update = 1'b0;
		// Trace: design.sv:42352:5
		perf_load_o = 1'b0;
		// Trace: design.sv:42353:5
		perf_store_o = 1'b0;
		// Trace: design.sv:42355:5
		(* full_case, parallel_case *)
		case (ls_fsm_cs)
			3'd0: begin
				// Trace: design.sv:42358:9
				pmp_err_d = 1'b0;
				// Trace: design.sv:42359:9
				if (lsu_req_i) begin
					// Trace: design.sv:42360:11
					data_req_o = 1'b1;
					// Trace: design.sv:42361:11
					pmp_err_d = data_pmp_err_i;
					// Trace: design.sv:42362:11
					lsu_err_d = 1'b0;
					// Trace: design.sv:42363:11
					perf_load_o = ~lsu_we_i;
					// Trace: design.sv:42364:11
					perf_store_o = lsu_we_i;
					// Trace: design.sv:42366:11
					if (data_gnt_i) begin
						// Trace: design.sv:42367:13
						ctrl_update = 1'b1;
						// Trace: design.sv:42368:13
						addr_update = 1'b1;
						// Trace: design.sv:42369:13
						handle_misaligned_d = split_misaligned_access;
						// Trace: design.sv:42370:13
						ls_fsm_ns = (split_misaligned_access ? 3'd2 : 3'd0);
					end
					else
						// Trace: design.sv:42372:13
						ls_fsm_ns = (split_misaligned_access ? 3'd1 : 3'd3);
				end
			end
			3'd1: begin
				// Trace: design.sv:42378:9
				data_req_o = 1'b1;
				// Trace: design.sv:42383:9
				if (data_gnt_i || pmp_err_q) begin
					// Trace: design.sv:42384:11
					addr_update = 1'b1;
					// Trace: design.sv:42385:11
					ctrl_update = 1'b1;
					// Trace: design.sv:42386:11
					handle_misaligned_d = 1'b1;
					// Trace: design.sv:42387:11
					ls_fsm_ns = 3'd2;
				end
			end
			3'd2: begin
				// Trace: design.sv:42393:9
				data_req_o = 1'b1;
				// Trace: design.sv:42395:9
				addr_incr_req_o = 1'b1;
				// Trace: design.sv:42398:9
				if (data_rvalid_i || pmp_err_q) begin
					// Trace: design.sv:42400:11
					pmp_err_d = data_pmp_err_i;
					// Trace: design.sv:42402:11
					lsu_err_d = data_err_i | pmp_err_q;
					// Trace: design.sv:42404:11
					rdata_update = ~data_we_q;
					// Trace: design.sv:42406:11
					ls_fsm_ns = (data_gnt_i ? 3'd0 : 3'd3);
					// Trace: design.sv:42408:11
					addr_update = data_gnt_i & ~(data_err_i | pmp_err_q);
					// Trace: design.sv:42410:11
					handle_misaligned_d = ~data_gnt_i;
				end
				else
					// Trace: design.sv:42413:11
					if (data_gnt_i) begin
						// Trace: design.sv:42415:13
						ls_fsm_ns = 3'd4;
						// Trace: design.sv:42416:13
						handle_misaligned_d = 1'b0;
					end
			end
			3'd3: begin
				// Trace: design.sv:42423:9
				addr_incr_req_o = handle_misaligned_q;
				// Trace: design.sv:42424:9
				data_req_o = 1'b1;
				// Trace: design.sv:42425:9
				if (data_gnt_i || pmp_err_q) begin
					// Trace: design.sv:42426:11
					ctrl_update = 1'b1;
					// Trace: design.sv:42428:11
					addr_update = ~lsu_err_q;
					// Trace: design.sv:42429:11
					ls_fsm_ns = 3'd0;
					// Trace: design.sv:42430:11
					handle_misaligned_d = 1'b0;
				end
			end
			3'd4: begin
				// Trace: design.sv:42437:9
				addr_incr_req_o = 1'b1;
				// Trace: design.sv:42439:9
				if (data_rvalid_i) begin
					// Trace: design.sv:42441:11
					pmp_err_d = data_pmp_err_i;
					// Trace: design.sv:42443:11
					lsu_err_d = data_err_i;
					// Trace: design.sv:42445:11
					addr_update = ~data_err_i;
					// Trace: design.sv:42447:11
					rdata_update = ~data_we_q;
					// Trace: design.sv:42449:11
					ls_fsm_ns = 3'd0;
				end
			end
			default:
				// Trace: design.sv:42454:9
				ls_fsm_ns = 3'd0;
		endcase
	end
	// Trace: design.sv:42459:3
	assign lsu_req_done_o = (lsu_req_i | (ls_fsm_cs != 3'd0)) & (ls_fsm_ns == 3'd0);
	// Trace: design.sv:42462:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:42463:5
		if (!rst_ni) begin
			// Trace: design.sv:42464:7
			ls_fsm_cs <= 3'd0;
			// Trace: design.sv:42465:7
			handle_misaligned_q <= 1'sb0;
			// Trace: design.sv:42466:7
			pmp_err_q <= 1'sb0;
			// Trace: design.sv:42467:7
			lsu_err_q <= 1'sb0;
		end
		else begin
			// Trace: design.sv:42469:7
			ls_fsm_cs <= ls_fsm_ns;
			// Trace: design.sv:42470:7
			handle_misaligned_q <= handle_misaligned_d;
			// Trace: design.sv:42471:7
			pmp_err_q <= pmp_err_d;
			// Trace: design.sv:42472:7
			lsu_err_q <= lsu_err_d;
		end
	// Trace: design.sv:42480:3
	assign data_or_pmp_err = (lsu_err_q | data_err_i) | pmp_err_q;
	// Trace: design.sv:42481:3
	assign lsu_resp_valid_o = (data_rvalid_i | pmp_err_q) & (ls_fsm_cs == 3'd0);
	// Trace: design.sv:42482:3
	assign lsu_rdata_valid_o = (((ls_fsm_cs == 3'd0) & data_rvalid_i) & ~data_or_pmp_err) & ~data_we_q;
	// Trace: design.sv:42485:3
	assign lsu_rdata_o = data_rdata_ext;
	// Trace: design.sv:42488:3
	assign data_addr_w_aligned = {data_addr[31:2], 2'b00};
	// Trace: design.sv:42491:3
	assign data_addr_o = data_addr_w_aligned;
	// Trace: design.sv:42492:3
	assign data_wdata_o = data_wdata;
	// Trace: design.sv:42493:3
	assign data_we_o = lsu_we_i;
	// Trace: design.sv:42494:3
	assign data_be_o = data_be;
	// Trace: design.sv:42497:3
	assign addr_last_o = addr_last_q;
	// Trace: design.sv:42500:3
	assign load_err_o = (data_or_pmp_err & ~data_we_q) & lsu_resp_valid_o;
	// Trace: design.sv:42501:3
	assign store_err_o = (data_or_pmp_err & data_we_q) & lsu_resp_valid_o;
	// Trace: design.sv:42503:3
	assign busy_o = ls_fsm_cs != 3'd0;
	initial _sv2v_0 = 0;
endmodule
module ibex_multdiv_fast (
	clk_i,
	rst_ni,
	mult_en_i,
	div_en_i,
	mult_sel_i,
	div_sel_i,
	operator_i,
	signed_mode_i,
	op_a_i,
	op_b_i,
	alu_adder_ext_i,
	alu_adder_i,
	equal_to_zero_i,
	data_ind_timing_i,
	alu_operand_a_o,
	alu_operand_b_o,
	imd_val_q_i,
	imd_val_d_o,
	imd_val_we_o,
	multdiv_ready_id_i,
	multdiv_result_o,
	valid_o
);
	reg _sv2v_0;
	// Trace: design.sv:42549:13
	// removed localparam type ibex_pkg_rv32m_e
	parameter integer RV32M = 32'sd2;
	// Trace: design.sv:42551:3
	input wire clk_i;
	// Trace: design.sv:42552:3
	input wire rst_ni;
	// Trace: design.sv:42553:3
	input wire mult_en_i;
	// Trace: design.sv:42554:3
	input wire div_en_i;
	// Trace: design.sv:42555:3
	input wire mult_sel_i;
	// Trace: design.sv:42556:3
	input wire div_sel_i;
	// Trace: design.sv:42557:3
	// removed localparam type ibex_pkg_md_op_e
	input wire [1:0] operator_i;
	// Trace: design.sv:42558:3
	input wire [1:0] signed_mode_i;
	// Trace: design.sv:42559:3
	input wire [31:0] op_a_i;
	// Trace: design.sv:42560:3
	input wire [31:0] op_b_i;
	// Trace: design.sv:42561:3
	input wire [33:0] alu_adder_ext_i;
	// Trace: design.sv:42562:3
	input wire [31:0] alu_adder_i;
	// Trace: design.sv:42563:3
	input wire equal_to_zero_i;
	// Trace: design.sv:42564:3
	input wire data_ind_timing_i;
	// Trace: design.sv:42566:3
	output reg [32:0] alu_operand_a_o;
	// Trace: design.sv:42567:3
	output reg [32:0] alu_operand_b_o;
	// Trace: design.sv:42569:3
	input wire [67:0] imd_val_q_i;
	// Trace: design.sv:42570:3
	output wire [67:0] imd_val_d_o;
	// Trace: design.sv:42571:3
	output wire [1:0] imd_val_we_o;
	// Trace: design.sv:42573:3
	input wire multdiv_ready_id_i;
	// Trace: design.sv:42575:3
	output wire [31:0] multdiv_result_o;
	// Trace: design.sv:42576:3
	output wire valid_o;
	// Trace: design.sv:42579:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:42582:3
	wire signed [34:0] mac_res_signed;
	// Trace: design.sv:42583:3
	wire [34:0] mac_res_ext;
	// Trace: design.sv:42584:3
	reg [33:0] accum;
	// Trace: design.sv:42585:3
	reg sign_a;
	reg sign_b;
	// Trace: design.sv:42586:3
	reg mult_valid;
	// Trace: design.sv:42587:3
	wire signed_mult;
	// Trace: design.sv:42590:3
	reg [33:0] mac_res_d;
	reg [33:0] op_remainder_d;
	// Trace: design.sv:42592:3
	wire [33:0] mac_res;
	// Trace: design.sv:42595:3
	wire div_sign_a;
	wire div_sign_b;
	// Trace: design.sv:42596:3
	reg is_greater_equal;
	// Trace: design.sv:42597:3
	wire div_change_sign;
	wire rem_change_sign;
	// Trace: design.sv:42598:3
	wire [31:0] one_shift;
	// Trace: design.sv:42599:3
	wire [31:0] op_denominator_q;
	// Trace: design.sv:42600:3
	reg [31:0] op_numerator_q;
	// Trace: design.sv:42601:3
	reg [31:0] op_quotient_q;
	// Trace: design.sv:42602:3
	reg [31:0] op_denominator_d;
	// Trace: design.sv:42603:3
	reg [31:0] op_numerator_d;
	// Trace: design.sv:42604:3
	reg [31:0] op_quotient_d;
	// Trace: design.sv:42605:3
	wire [31:0] next_remainder;
	// Trace: design.sv:42606:3
	wire [32:0] next_quotient;
	// Trace: design.sv:42607:3
	wire [31:0] res_adder_h;
	// Trace: design.sv:42608:3
	reg div_valid;
	// Trace: design.sv:42609:3
	reg [4:0] div_counter_q;
	reg [4:0] div_counter_d;
	// Trace: design.sv:42610:3
	wire multdiv_en;
	// Trace: design.sv:42611:3
	reg mult_hold;
	// Trace: design.sv:42612:3
	reg div_hold;
	// Trace: design.sv:42613:3
	reg div_by_zero_d;
	reg div_by_zero_q;
	// Trace: design.sv:42615:3
	wire mult_en_internal;
	// Trace: design.sv:42616:3
	wire div_en_internal;
	// Trace: design.sv:42618:3
	// removed localparam type md_fsm_e
	// Trace: design.sv:42621:3
	reg [2:0] md_state_q;
	reg [2:0] md_state_d;
	// Trace: design.sv:42623:3
	wire unused_mult_sel_i;
	// Trace: design.sv:42624:3
	assign unused_mult_sel_i = mult_sel_i;
	// Trace: design.sv:42626:3
	assign mult_en_internal = mult_en_i & ~mult_hold;
	// Trace: design.sv:42627:3
	assign div_en_internal = div_en_i & ~div_hold;
	// Trace: design.sv:42629:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:42630:5
		if (!rst_ni) begin
			// Trace: design.sv:42631:7
			div_counter_q <= 1'sb0;
			// Trace: design.sv:42632:7
			md_state_q <= 3'd0;
			// Trace: design.sv:42633:7
			op_numerator_q <= 1'sb0;
			// Trace: design.sv:42634:7
			op_quotient_q <= 1'sb0;
			// Trace: design.sv:42635:7
			div_by_zero_q <= 1'sb0;
		end
		else if (div_en_internal) begin
			// Trace: design.sv:42637:7
			div_counter_q <= div_counter_d;
			// Trace: design.sv:42638:7
			op_numerator_q <= op_numerator_d;
			// Trace: design.sv:42639:7
			op_quotient_q <= op_quotient_d;
			// Trace: design.sv:42640:7
			md_state_q <= md_state_d;
			// Trace: design.sv:42641:7
			div_by_zero_q <= div_by_zero_d;
		end
	// Trace: design.sv:42649:3
	assign multdiv_en = mult_en_internal | div_en_internal;
	// Trace: design.sv:42652:3
	assign imd_val_d_o[34+:34] = (div_sel_i ? op_remainder_d : mac_res_d);
	// Trace: design.sv:42653:3
	assign imd_val_we_o[0] = multdiv_en;
	// Trace: design.sv:42655:3
	assign imd_val_d_o[0+:34] = {2'b00, op_denominator_d};
	// Trace: design.sv:42656:3
	assign imd_val_we_o[1] = div_en_internal;
	// Trace: design.sv:42657:3
	assign op_denominator_q = imd_val_q_i[31-:32];
	// Trace: design.sv:42658:3
	wire [1:0] unused_imd_val;
	// Trace: design.sv:42659:3
	assign unused_imd_val = imd_val_q_i[33-:2];
	// Trace: design.sv:42660:3
	wire unused_mac_res_ext;
	// Trace: design.sv:42661:3
	assign unused_mac_res_ext = mac_res_ext[34];
	// Trace: design.sv:42663:3
	assign signed_mult = signed_mode_i != 2'b00;
	// Trace: design.sv:42664:3
	assign multdiv_result_o = (div_sel_i ? imd_val_q_i[65-:32] : mac_res_d[31:0]);
	// Trace: design.sv:42668:3
	generate
		if (RV32M == 32'sd3) begin : gen_mult_single_cycle
			// Trace: design.sv:42670:5
			// removed localparam type mult_fsm_e
			// Trace: design.sv:42673:5
			reg mult_state_q;
			reg mult_state_d;
			// Trace: design.sv:42675:5
			wire signed [33:0] mult1_res;
			wire signed [33:0] mult2_res;
			wire signed [33:0] mult3_res;
			// Trace: design.sv:42676:5
			wire [33:0] mult1_res_uns;
			// Trace: design.sv:42677:5
			wire [33:32] unused_mult1_res_uns;
			// Trace: design.sv:42678:5
			wire [15:0] mult1_op_a;
			wire [15:0] mult1_op_b;
			// Trace: design.sv:42679:5
			wire [15:0] mult2_op_a;
			wire [15:0] mult2_op_b;
			// Trace: design.sv:42680:5
			reg [15:0] mult3_op_a;
			reg [15:0] mult3_op_b;
			// Trace: design.sv:42681:5
			wire mult1_sign_a;
			wire mult1_sign_b;
			// Trace: design.sv:42682:5
			wire mult2_sign_a;
			wire mult2_sign_b;
			// Trace: design.sv:42683:5
			reg mult3_sign_a;
			reg mult3_sign_b;
			// Trace: design.sv:42684:5
			reg [33:0] summand1;
			reg [33:0] summand2;
			reg [33:0] summand3;
			// Trace: design.sv:42686:5
			assign mult1_res = $signed({mult1_sign_a, mult1_op_a}) * $signed({mult1_sign_b, mult1_op_b});
			// Trace: design.sv:42687:5
			assign mult2_res = $signed({mult2_sign_a, mult2_op_a}) * $signed({mult2_sign_b, mult2_op_b});
			// Trace: design.sv:42688:5
			assign mult3_res = $signed({mult3_sign_a, mult3_op_a}) * $signed({mult3_sign_b, mult3_op_b});
			// Trace: design.sv:42690:5
			assign mac_res_signed = ($signed(summand1) + $signed(summand2)) + $signed(summand3);
			// Trace: design.sv:42692:5
			assign mult1_res_uns = $unsigned(mult1_res);
			// Trace: design.sv:42693:5
			assign mac_res_ext = $unsigned(mac_res_signed);
			// Trace: design.sv:42694:5
			assign mac_res = mac_res_ext[33:0];
			// Trace: design.sv:42696:5
			wire [1:1] sv2v_tmp_5ADA8;
			assign sv2v_tmp_5ADA8 = signed_mode_i[0] & op_a_i[31];
			always @(*) sign_a = sv2v_tmp_5ADA8;
			// Trace: design.sv:42697:5
			wire [1:1] sv2v_tmp_C5449;
			assign sv2v_tmp_C5449 = signed_mode_i[1] & op_b_i[31];
			always @(*) sign_b = sv2v_tmp_C5449;
			// Trace: design.sv:42701:5
			assign mult1_sign_a = 1'b0;
			// Trace: design.sv:42702:5
			assign mult1_sign_b = 1'b0;
			// Trace: design.sv:42703:5
			assign mult1_op_a = op_a_i[15:0];
			// Trace: design.sv:42704:5
			assign mult1_op_b = op_b_i[15:0];
			// Trace: design.sv:42707:5
			assign mult2_sign_a = 1'b0;
			// Trace: design.sv:42708:5
			assign mult2_sign_b = sign_b;
			// Trace: design.sv:42709:5
			assign mult2_op_a = op_a_i[15:0];
			// Trace: design.sv:42710:5
			assign mult2_op_b = op_b_i[31:16];
			// Trace: design.sv:42713:5
			wire [18:1] sv2v_tmp_6FF3F;
			assign sv2v_tmp_6FF3F = imd_val_q_i[67-:18];
			always @(*) accum[17:0] = sv2v_tmp_6FF3F;
			// Trace: design.sv:42714:5
			wire [16:1] sv2v_tmp_A7770;
			assign sv2v_tmp_A7770 = {16 {signed_mult & imd_val_q_i[67]}};
			always @(*) accum[33:18] = sv2v_tmp_A7770;
			// Trace: design.sv:42716:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:42720:7
				mult3_sign_a = sign_a;
				// Trace: design.sv:42721:7
				mult3_sign_b = 1'b0;
				// Trace: design.sv:42722:7
				mult3_op_a = op_a_i[31:16];
				// Trace: design.sv:42723:7
				mult3_op_b = op_b_i[15:0];
				// Trace: design.sv:42725:7
				summand1 = {18'h00000, mult1_res_uns[31:16]};
				// Trace: design.sv:42726:7
				summand2 = $unsigned(mult2_res);
				// Trace: design.sv:42727:7
				summand3 = $unsigned(mult3_res);
				// Trace: design.sv:42730:7
				mac_res_d = {2'b00, mac_res[15:0], mult1_res_uns[15:0]};
				// Trace: design.sv:42731:7
				mult_valid = mult_en_i;
				// Trace: design.sv:42732:7
				mult_state_d = 1'd0;
				// Trace: design.sv:42734:7
				mult_hold = 1'b0;
				// Trace: design.sv:42736:7
				(* full_case, parallel_case *)
				case (mult_state_q)
					1'd0:
						// Trace: design.sv:42739:11
						if (operator_i != 2'd0) begin
							// Trace: design.sv:42740:13
							mac_res_d = mac_res;
							// Trace: design.sv:42741:13
							mult_valid = 1'b0;
							// Trace: design.sv:42742:13
							mult_state_d = 1'd1;
						end
						else
							// Trace: design.sv:42744:13
							mult_hold = ~multdiv_ready_id_i;
					1'd1: begin
						// Trace: design.sv:42750:11
						mult3_sign_a = sign_a;
						// Trace: design.sv:42751:11
						mult3_sign_b = sign_b;
						// Trace: design.sv:42752:11
						mult3_op_a = op_a_i[31:16];
						// Trace: design.sv:42753:11
						mult3_op_b = op_b_i[31:16];
						// Trace: design.sv:42754:11
						mac_res_d = mac_res;
						// Trace: design.sv:42756:11
						summand1 = 1'sb0;
						// Trace: design.sv:42757:11
						summand2 = accum;
						// Trace: design.sv:42758:11
						summand3 = $unsigned(mult3_res);
						// Trace: design.sv:42760:11
						mult_state_d = 1'd0;
						// Trace: design.sv:42761:11
						mult_valid = 1'b1;
						// Trace: design.sv:42763:11
						mult_hold = ~multdiv_ready_id_i;
					end
					default:
						// Trace: design.sv:42767:11
						mult_state_d = 1'd0;
				endcase
			end
			// Trace: design.sv:42773:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:42774:7
				if (!rst_ni)
					// Trace: design.sv:42775:9
					mult_state_q <= 1'd0;
				else
					// Trace: design.sv:42777:9
					if (mult_en_internal)
						// Trace: design.sv:42778:11
						mult_state_q <= mult_state_d;
			// Trace: design.sv:42783:5
			assign unused_mult1_res_uns = mult1_res_uns[33:32];
		end
		else begin : gen_mult_fast
			// Trace: design.sv:42791:5
			reg [15:0] mult_op_a;
			// Trace: design.sv:42792:5
			reg [15:0] mult_op_b;
			// Trace: design.sv:42794:5
			// removed localparam type mult_fsm_e
			// Trace: design.sv:42797:5
			reg [1:0] mult_state_q;
			reg [1:0] mult_state_d;
			// Trace: design.sv:42803:5
			assign mac_res_signed = ($signed({sign_a, mult_op_a}) * $signed({sign_b, mult_op_b})) + $signed(accum);
			// Trace: design.sv:42805:5
			assign mac_res_ext = $unsigned(mac_res_signed);
			// Trace: design.sv:42806:5
			assign mac_res = mac_res_ext[33:0];
			// Trace: design.sv:42808:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:42809:7
				mult_op_a = op_a_i[15:0];
				// Trace: design.sv:42810:7
				mult_op_b = op_b_i[15:0];
				// Trace: design.sv:42811:7
				sign_a = 1'b0;
				// Trace: design.sv:42812:7
				sign_b = 1'b0;
				// Trace: design.sv:42813:7
				accum = imd_val_q_i[34+:34];
				// Trace: design.sv:42814:7
				mac_res_d = mac_res;
				// Trace: design.sv:42815:7
				mult_state_d = mult_state_q;
				// Trace: design.sv:42816:7
				mult_valid = 1'b0;
				// Trace: design.sv:42817:7
				mult_hold = 1'b0;
				// Trace: design.sv:42819:7
				(* full_case, parallel_case *)
				case (mult_state_q)
					2'd0: begin
						// Trace: design.sv:42823:11
						mult_op_a = op_a_i[15:0];
						// Trace: design.sv:42824:11
						mult_op_b = op_b_i[15:0];
						// Trace: design.sv:42825:11
						sign_a = 1'b0;
						// Trace: design.sv:42826:11
						sign_b = 1'b0;
						// Trace: design.sv:42827:11
						accum = 1'sb0;
						// Trace: design.sv:42828:11
						mac_res_d = mac_res;
						// Trace: design.sv:42829:11
						mult_state_d = 2'd1;
					end
					2'd1: begin
						// Trace: design.sv:42834:11
						mult_op_a = op_a_i[15:0];
						// Trace: design.sv:42835:11
						mult_op_b = op_b_i[31:16];
						// Trace: design.sv:42836:11
						sign_a = 1'b0;
						// Trace: design.sv:42837:11
						sign_b = signed_mode_i[1] & op_b_i[31];
						// Trace: design.sv:42839:11
						accum = {18'b000000000000000000, imd_val_q_i[65-:16]};
						// Trace: design.sv:42840:11
						if (operator_i == 2'd0)
							// Trace: design.sv:42841:13
							mac_res_d = {2'b00, mac_res[15:0], imd_val_q_i[49-:16]};
						else
							// Trace: design.sv:42844:13
							mac_res_d = mac_res;
						// Trace: design.sv:42846:11
						mult_state_d = 2'd2;
					end
					2'd2: begin
						// Trace: design.sv:42851:11
						mult_op_a = op_a_i[31:16];
						// Trace: design.sv:42852:11
						mult_op_b = op_b_i[15:0];
						// Trace: design.sv:42853:11
						sign_a = signed_mode_i[0] & op_a_i[31];
						// Trace: design.sv:42854:11
						sign_b = 1'b0;
						// Trace: design.sv:42855:11
						if (operator_i == 2'd0) begin
							// Trace: design.sv:42856:13
							accum = {18'b000000000000000000, imd_val_q_i[65-:16]};
							// Trace: design.sv:42857:13
							mac_res_d = {2'b00, mac_res[15:0], imd_val_q_i[49-:16]};
							// Trace: design.sv:42858:13
							mult_valid = 1'b1;
							// Trace: design.sv:42861:13
							mult_state_d = 2'd0;
							// Trace: design.sv:42862:13
							mult_hold = ~multdiv_ready_id_i;
						end
						else begin
							// Trace: design.sv:42864:13
							accum = imd_val_q_i[34+:34];
							// Trace: design.sv:42865:13
							mac_res_d = mac_res;
							// Trace: design.sv:42866:13
							mult_state_d = 2'd3;
						end
					end
					2'd3: begin
						// Trace: design.sv:42873:11
						mult_op_a = op_a_i[31:16];
						// Trace: design.sv:42874:11
						mult_op_b = op_b_i[31:16];
						// Trace: design.sv:42875:11
						sign_a = signed_mode_i[0] & op_a_i[31];
						// Trace: design.sv:42876:11
						sign_b = signed_mode_i[1] & op_b_i[31];
						// Trace: design.sv:42877:11
						accum[17:0] = imd_val_q_i[67-:18];
						// Trace: design.sv:42878:11
						accum[33:18] = {16 {signed_mult & imd_val_q_i[67]}};
						// Trace: design.sv:42880:11
						mac_res_d = mac_res;
						// Trace: design.sv:42881:11
						mult_valid = 1'b1;
						// Trace: design.sv:42884:11
						mult_state_d = 2'd0;
						// Trace: design.sv:42885:11
						mult_hold = ~multdiv_ready_id_i;
					end
					default:
						// Trace: design.sv:42888:11
						mult_state_d = 2'd0;
				endcase
			end
			// Trace: design.sv:42893:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:42894:7
				if (!rst_ni)
					// Trace: design.sv:42895:9
					mult_state_q <= 2'd0;
				else
					// Trace: design.sv:42897:9
					if (mult_en_internal)
						// Trace: design.sv:42898:11
						mult_state_q <= mult_state_d;
		end
	endgenerate
	// Trace: design.sv:42909:3
	assign res_adder_h = alu_adder_ext_i[32:1];
	// Trace: design.sv:42910:3
	wire [1:0] unused_alu_adder_ext;
	// Trace: design.sv:42911:3
	assign unused_alu_adder_ext = {alu_adder_ext_i[33], alu_adder_ext_i[0]};
	// Trace: design.sv:42913:3
	assign next_remainder = (is_greater_equal ? res_adder_h[31:0] : imd_val_q_i[65-:32]);
	// Trace: design.sv:42914:3
	assign next_quotient = (is_greater_equal ? {1'b0, op_quotient_q} | {1'b0, one_shift} : {1'b0, op_quotient_q});
	// Trace: design.sv:42917:3
	assign one_shift = 32'b00000000000000000000000000000001 << div_counter_q;
	// Trace: design.sv:42922:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42923:5
		if ((imd_val_q_i[65] ^ op_denominator_q[31]) == 1'b0)
			// Trace: design.sv:42924:7
			is_greater_equal = res_adder_h[31] == 1'b0;
		else
			// Trace: design.sv:42926:7
			is_greater_equal = imd_val_q_i[65];
	end
	// Trace: design.sv:42930:3
	assign div_sign_a = op_a_i[31] & signed_mode_i[0];
	// Trace: design.sv:42931:3
	assign div_sign_b = op_b_i[31] & signed_mode_i[1];
	// Trace: design.sv:42932:3
	assign div_change_sign = (div_sign_a ^ div_sign_b) & ~div_by_zero_q;
	// Trace: design.sv:42933:3
	assign rem_change_sign = div_sign_a;
	// Trace: design.sv:42936:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:42937:5
		div_counter_d = div_counter_q - 5'h01;
		// Trace: design.sv:42938:5
		op_remainder_d = imd_val_q_i[34+:34];
		// Trace: design.sv:42939:5
		op_quotient_d = op_quotient_q;
		// Trace: design.sv:42940:5
		md_state_d = md_state_q;
		// Trace: design.sv:42941:5
		op_numerator_d = op_numerator_q;
		// Trace: design.sv:42942:5
		op_denominator_d = op_denominator_q;
		// Trace: design.sv:42943:5
		alu_operand_a_o = 33'h000000001;
		// Trace: design.sv:42944:5
		alu_operand_b_o = {~op_b_i, 1'b1};
		// Trace: design.sv:42945:5
		div_valid = 1'b0;
		// Trace: design.sv:42946:5
		div_hold = 1'b0;
		// Trace: design.sv:42947:5
		div_by_zero_d = div_by_zero_q;
		// Trace: design.sv:42949:5
		(* full_case, parallel_case *)
		case (md_state_q)
			3'd0: begin
				// Trace: design.sv:42951:9
				if (operator_i == 2'd2) begin
					// Trace: design.sv:42956:11
					op_remainder_d = 1'sb1;
					// Trace: design.sv:42958:11
					md_state_d = (!data_ind_timing_i && equal_to_zero_i ? 3'd6 : 3'd1);
					// Trace: design.sv:42961:11
					div_by_zero_d = equal_to_zero_i;
				end
				else begin
					// Trace: design.sv:42967:11
					op_remainder_d = {2'b00, op_a_i};
					// Trace: design.sv:42969:11
					md_state_d = (!data_ind_timing_i && equal_to_zero_i ? 3'd6 : 3'd1);
				end
				// Trace: design.sv:42972:9
				alu_operand_a_o = 33'h000000001;
				// Trace: design.sv:42973:9
				alu_operand_b_o = {~op_b_i, 1'b1};
				// Trace: design.sv:42974:9
				div_counter_d = 5'd31;
			end
			3'd1: begin
				// Trace: design.sv:42979:9
				op_quotient_d = 1'sb0;
				// Trace: design.sv:42981:9
				op_numerator_d = (div_sign_a ? alu_adder_i : op_a_i);
				// Trace: design.sv:42982:9
				md_state_d = 3'd2;
				// Trace: design.sv:42983:9
				div_counter_d = 5'd31;
				// Trace: design.sv:42985:9
				alu_operand_a_o = 33'h000000001;
				// Trace: design.sv:42986:9
				alu_operand_b_o = {~op_a_i, 1'b1};
			end
			3'd2: begin
				// Trace: design.sv:42991:9
				op_remainder_d = {33'h000000000, op_numerator_q[31]};
				// Trace: design.sv:42993:9
				op_denominator_d = (div_sign_b ? alu_adder_i : op_b_i);
				// Trace: design.sv:42994:9
				md_state_d = 3'd3;
				// Trace: design.sv:42995:9
				div_counter_d = 5'd31;
				// Trace: design.sv:42997:9
				alu_operand_a_o = 33'h000000001;
				// Trace: design.sv:42998:9
				alu_operand_b_o = {~op_b_i, 1'b1};
			end
			3'd3: begin
				// Trace: design.sv:43002:9
				op_remainder_d = {1'b0, next_remainder[31:0], op_numerator_q[div_counter_d]};
				// Trace: design.sv:43003:9
				op_quotient_d = next_quotient[31:0];
				// Trace: design.sv:43004:9
				md_state_d = (div_counter_q == 5'd1 ? 3'd4 : 3'd3);
				// Trace: design.sv:43006:9
				alu_operand_a_o = {imd_val_q_i[65-:32], 1'b1};
				// Trace: design.sv:43007:9
				alu_operand_b_o = {~op_denominator_q[31:0], 1'b1};
			end
			3'd4: begin
				// Trace: design.sv:43011:9
				if (operator_i == 2'd2)
					// Trace: design.sv:43014:11
					op_remainder_d = {1'b0, next_quotient};
				else
					// Trace: design.sv:43017:11
					op_remainder_d = {2'b00, next_remainder[31:0]};
				// Trace: design.sv:43020:9
				alu_operand_a_o = {imd_val_q_i[65-:32], 1'b1};
				// Trace: design.sv:43021:9
				alu_operand_b_o = {~op_denominator_q[31:0], 1'b1};
				// Trace: design.sv:43023:9
				md_state_d = 3'd5;
			end
			3'd5: begin
				// Trace: design.sv:43027:9
				md_state_d = 3'd6;
				// Trace: design.sv:43028:9
				if (operator_i == 2'd2)
					// Trace: design.sv:43029:11
					op_remainder_d = (div_change_sign ? {2'h0, alu_adder_i} : imd_val_q_i[34+:34]);
				else
					// Trace: design.sv:43031:11
					op_remainder_d = (rem_change_sign ? {2'h0, alu_adder_i} : imd_val_q_i[34+:34]);
				// Trace: design.sv:43034:9
				alu_operand_a_o = 33'h000000001;
				// Trace: design.sv:43035:9
				alu_operand_b_o = {~imd_val_q_i[65-:32], 1'b1};
			end
			3'd6: begin
				// Trace: design.sv:43041:9
				md_state_d = 3'd0;
				// Trace: design.sv:43042:9
				div_hold = ~multdiv_ready_id_i;
				// Trace: design.sv:43043:9
				div_valid = 1'b1;
			end
			default:
				// Trace: design.sv:43047:9
				md_state_d = 3'd0;
		endcase
	end
	// Trace: design.sv:43052:3
	assign valid_o = mult_valid | div_valid;
	initial _sv2v_0 = 0;
endmodule
module ibex_multdiv_slow (
	clk_i,
	rst_ni,
	mult_en_i,
	div_en_i,
	mult_sel_i,
	div_sel_i,
	operator_i,
	signed_mode_i,
	op_a_i,
	op_b_i,
	alu_adder_ext_i,
	alu_adder_i,
	equal_to_zero_i,
	data_ind_timing_i,
	alu_operand_a_o,
	alu_operand_b_o,
	imd_val_q_i,
	imd_val_d_o,
	imd_val_we_o,
	multdiv_ready_id_i,
	multdiv_result_o,
	valid_o
);
	reg _sv2v_0;
	// Trace: design.sv:43080:3
	input wire clk_i;
	// Trace: design.sv:43081:3
	input wire rst_ni;
	// Trace: design.sv:43082:3
	input wire mult_en_i;
	// Trace: design.sv:43083:3
	input wire div_en_i;
	// Trace: design.sv:43084:3
	input wire mult_sel_i;
	// Trace: design.sv:43085:3
	input wire div_sel_i;
	// Trace: design.sv:43086:3
	// removed localparam type ibex_pkg_md_op_e
	input wire [1:0] operator_i;
	// Trace: design.sv:43087:3
	input wire [1:0] signed_mode_i;
	// Trace: design.sv:43088:3
	input wire [31:0] op_a_i;
	// Trace: design.sv:43089:3
	input wire [31:0] op_b_i;
	// Trace: design.sv:43090:3
	input wire [33:0] alu_adder_ext_i;
	// Trace: design.sv:43091:3
	input wire [31:0] alu_adder_i;
	// Trace: design.sv:43092:3
	input wire equal_to_zero_i;
	// Trace: design.sv:43093:3
	input wire data_ind_timing_i;
	// Trace: design.sv:43095:3
	output reg [32:0] alu_operand_a_o;
	// Trace: design.sv:43096:3
	output reg [32:0] alu_operand_b_o;
	// Trace: design.sv:43098:3
	input wire [67:0] imd_val_q_i;
	// Trace: design.sv:43099:3
	output wire [67:0] imd_val_d_o;
	// Trace: design.sv:43100:3
	output wire [1:0] imd_val_we_o;
	// Trace: design.sv:43102:3
	input wire multdiv_ready_id_i;
	// Trace: design.sv:43104:3
	output wire [31:0] multdiv_result_o;
	// Trace: design.sv:43106:3
	output wire valid_o;
	// Trace: design.sv:43109:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:43111:3
	// removed localparam type md_fsm_e
	// Trace: design.sv:43114:3
	reg [2:0] md_state_q;
	reg [2:0] md_state_d;
	// Trace: design.sv:43116:3
	wire [32:0] accum_window_q;
	reg [32:0] accum_window_d;
	// Trace: design.sv:43117:3
	wire unused_imd_val0;
	// Trace: design.sv:43118:3
	wire [1:0] unused_imd_val1;
	// Trace: design.sv:43120:3
	wire [32:0] res_adder_l;
	// Trace: design.sv:43121:3
	wire [32:0] res_adder_h;
	// Trace: design.sv:43123:3
	reg [4:0] multdiv_count_q;
	reg [4:0] multdiv_count_d;
	// Trace: design.sv:43124:3
	reg [32:0] op_b_shift_q;
	reg [32:0] op_b_shift_d;
	// Trace: design.sv:43125:3
	reg [32:0] op_a_shift_q;
	reg [32:0] op_a_shift_d;
	// Trace: design.sv:43126:3
	wire [32:0] op_a_ext;
	wire [32:0] op_b_ext;
	// Trace: design.sv:43127:3
	wire [32:0] one_shift;
	// Trace: design.sv:43128:3
	wire [32:0] op_a_bw_pp;
	wire [32:0] op_a_bw_last_pp;
	// Trace: design.sv:43129:3
	wire [31:0] b_0;
	// Trace: design.sv:43130:3
	wire sign_a;
	wire sign_b;
	// Trace: design.sv:43131:3
	wire [32:0] next_quotient;
	// Trace: design.sv:43132:3
	wire [31:0] next_remainder;
	// Trace: design.sv:43133:3
	wire [31:0] op_numerator_q;
	reg [31:0] op_numerator_d;
	// Trace: design.sv:43134:3
	wire is_greater_equal;
	// Trace: design.sv:43135:3
	wire div_change_sign;
	wire rem_change_sign;
	// Trace: design.sv:43136:3
	reg div_by_zero_d;
	reg div_by_zero_q;
	// Trace: design.sv:43137:3
	reg multdiv_hold;
	// Trace: design.sv:43138:3
	wire multdiv_en;
	// Trace: design.sv:43141:3
	assign res_adder_l = alu_adder_ext_i[32:0];
	// Trace: design.sv:43143:3
	assign res_adder_h = alu_adder_ext_i[33:1];
	// Trace: design.sv:43150:3
	assign imd_val_d_o[34+:34] = {1'b0, accum_window_d};
	// Trace: design.sv:43151:3
	assign imd_val_we_o[0] = ~multdiv_hold;
	// Trace: design.sv:43152:3
	assign accum_window_q = imd_val_q_i[66-:33];
	// Trace: design.sv:43153:3
	assign unused_imd_val0 = imd_val_q_i[67];
	// Trace: design.sv:43155:3
	assign imd_val_d_o[0+:34] = {2'b00, op_numerator_d};
	// Trace: design.sv:43156:3
	assign imd_val_we_o[1] = multdiv_en;
	// Trace: design.sv:43157:3
	assign op_numerator_q = imd_val_q_i[31-:32];
	// Trace: design.sv:43158:3
	assign unused_imd_val1 = imd_val_q_i[33-:2];
	// Trace: design.sv:43160:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:43161:5
		alu_operand_a_o = accum_window_q;
		// Trace: design.sv:43163:5
		(* full_case, parallel_case *)
		case (operator_i)
			2'd0:
				// Trace: design.sv:43166:9
				alu_operand_b_o = op_a_bw_pp;
			2'd1:
				// Trace: design.sv:43170:9
				alu_operand_b_o = (md_state_q == 3'd4 ? op_a_bw_last_pp : op_a_bw_pp);
			2'd2, 2'd3:
				// Trace: design.sv:43175:9
				(* full_case, parallel_case *)
				case (md_state_q)
					3'd0: begin
						// Trace: design.sv:43178:13
						alu_operand_a_o = 33'h000000001;
						// Trace: design.sv:43179:13
						alu_operand_b_o = {~op_b_i, 1'b1};
					end
					3'd1: begin
						// Trace: design.sv:43183:13
						alu_operand_a_o = 33'h000000001;
						// Trace: design.sv:43184:13
						alu_operand_b_o = {~op_a_i, 1'b1};
					end
					3'd2: begin
						// Trace: design.sv:43188:13
						alu_operand_a_o = 33'h000000001;
						// Trace: design.sv:43189:13
						alu_operand_b_o = {~op_b_i, 1'b1};
					end
					3'd5: begin
						// Trace: design.sv:43193:13
						alu_operand_a_o = 33'h000000001;
						// Trace: design.sv:43194:13
						alu_operand_b_o = {~accum_window_q[31:0], 1'b1};
					end
					default: begin
						// Trace: design.sv:43198:13
						alu_operand_a_o = {accum_window_q[31:0], 1'b1};
						// Trace: design.sv:43199:13
						alu_operand_b_o = {~op_b_shift_q[31:0], 1'b1};
					end
				endcase
			default: begin
				// Trace: design.sv:43204:9
				alu_operand_a_o = accum_window_q;
				// Trace: design.sv:43205:9
				alu_operand_b_o = {~op_b_shift_q[31:0], 1'b1};
			end
		endcase
	end
	// Trace: design.sv:43211:3
	assign b_0 = {32 {op_b_shift_q[0]}};
	// Trace: design.sv:43212:3
	assign op_a_bw_pp = {~(op_a_shift_q[32] & op_b_shift_q[0]), op_a_shift_q[31:0] & b_0};
	// Trace: design.sv:43213:3
	assign op_a_bw_last_pp = {op_a_shift_q[32] & op_b_shift_q[0], ~(op_a_shift_q[31:0] & b_0)};
	// Trace: design.sv:43216:3
	assign sign_a = op_a_i[31] & signed_mode_i[0];
	// Trace: design.sv:43217:3
	assign sign_b = op_b_i[31] & signed_mode_i[1];
	// Trace: design.sv:43219:3
	assign op_a_ext = {sign_a, op_a_i};
	// Trace: design.sv:43220:3
	assign op_b_ext = {sign_b, op_b_i};
	// Trace: design.sv:43227:3
	assign is_greater_equal = (accum_window_q[31] == op_b_shift_q[31] ? ~res_adder_h[31] : accum_window_q[31]);
	// Trace: design.sv:43230:3
	assign one_shift = 33'b000000000000000000000000000000001 << multdiv_count_q;
	// Trace: design.sv:43232:3
	assign next_remainder = (is_greater_equal ? res_adder_h[31:0] : accum_window_q[31:0]);
	// Trace: design.sv:43233:3
	assign next_quotient = (is_greater_equal ? op_a_shift_q | one_shift : op_a_shift_q);
	// Trace: design.sv:43235:3
	assign div_change_sign = (sign_a ^ sign_b) & ~div_by_zero_q;
	// Trace: design.sv:43236:3
	assign rem_change_sign = sign_a;
	// Trace: design.sv:43238:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:43239:5
		multdiv_count_d = multdiv_count_q;
		// Trace: design.sv:43240:5
		accum_window_d = accum_window_q;
		// Trace: design.sv:43241:5
		op_b_shift_d = op_b_shift_q;
		// Trace: design.sv:43242:5
		op_a_shift_d = op_a_shift_q;
		// Trace: design.sv:43243:5
		op_numerator_d = op_numerator_q;
		// Trace: design.sv:43244:5
		md_state_d = md_state_q;
		// Trace: design.sv:43245:5
		multdiv_hold = 1'b0;
		// Trace: design.sv:43246:5
		div_by_zero_d = div_by_zero_q;
		// Trace: design.sv:43247:5
		if (mult_sel_i || div_sel_i)
			// Trace: design.sv:43248:7
			(* full_case, parallel_case *)
			case (md_state_q)
				3'd0: begin
					// Trace: design.sv:43250:11
					(* full_case, parallel_case *)
					case (operator_i)
						2'd0: begin
							// Trace: design.sv:43252:15
							op_a_shift_d = op_a_ext << 1;
							// Trace: design.sv:43253:15
							accum_window_d = {~(op_a_ext[32] & op_b_i[0]), op_a_ext[31:0] & {32 {op_b_i[0]}}};
							// Trace: design.sv:43255:15
							op_b_shift_d = op_b_ext >> 1;
							// Trace: design.sv:43258:15
							md_state_d = (!data_ind_timing_i && ((op_b_ext >> 1) == 0) ? 3'd4 : 3'd3);
						end
						2'd1: begin
							// Trace: design.sv:43261:15
							op_a_shift_d = op_a_ext;
							// Trace: design.sv:43262:15
							accum_window_d = {1'b1, ~(op_a_ext[32] & op_b_i[0]), op_a_ext[31:1] & {31 {op_b_i[0]}}};
							// Trace: design.sv:43264:15
							op_b_shift_d = op_b_ext >> 1;
							// Trace: design.sv:43265:15
							md_state_d = 3'd3;
						end
						2'd2: begin
							// Trace: design.sv:43272:15
							accum_window_d = {33 {1'b1}};
							// Trace: design.sv:43274:15
							md_state_d = (!data_ind_timing_i && equal_to_zero_i ? 3'd6 : 3'd1);
							// Trace: design.sv:43277:15
							div_by_zero_d = equal_to_zero_i;
						end
						2'd3: begin
							// Trace: design.sv:43284:15
							accum_window_d = op_a_ext;
							// Trace: design.sv:43286:15
							md_state_d = (!data_ind_timing_i && equal_to_zero_i ? 3'd6 : 3'd1);
						end
						default:
							;
					endcase
					// Trace: design.sv:43290:11
					multdiv_count_d = 5'd31;
				end
				3'd1: begin
					// Trace: design.sv:43295:11
					op_a_shift_d = 1'sb0;
					// Trace: design.sv:43297:11
					op_numerator_d = (sign_a ? alu_adder_i : op_a_i);
					// Trace: design.sv:43298:11
					md_state_d = 3'd2;
				end
				3'd2: begin
					// Trace: design.sv:43303:11
					accum_window_d = {32'h00000000, op_numerator_q[31]};
					// Trace: design.sv:43305:11
					op_b_shift_d = (sign_b ? {1'b0, alu_adder_i} : {1'b0, op_b_i});
					// Trace: design.sv:43306:11
					md_state_d = 3'd3;
				end
				3'd3: begin
					// Trace: design.sv:43310:11
					multdiv_count_d = multdiv_count_q - 5'h01;
					// Trace: design.sv:43311:11
					(* full_case, parallel_case *)
					case (operator_i)
						2'd0: begin
							// Trace: design.sv:43313:15
							accum_window_d = res_adder_l;
							// Trace: design.sv:43314:15
							op_a_shift_d = op_a_shift_q << 1;
							// Trace: design.sv:43315:15
							op_b_shift_d = op_b_shift_q >> 1;
							// Trace: design.sv:43319:15
							md_state_d = ((!data_ind_timing_i && (op_b_shift_d == 0)) || (multdiv_count_q == 5'd1) ? 3'd4 : 3'd3);
						end
						2'd1: begin
							// Trace: design.sv:43323:15
							accum_window_d = res_adder_h;
							// Trace: design.sv:43324:15
							op_a_shift_d = op_a_shift_q;
							// Trace: design.sv:43325:15
							op_b_shift_d = op_b_shift_q >> 1;
							// Trace: design.sv:43326:15
							md_state_d = (multdiv_count_q == 5'd1 ? 3'd4 : 3'd3);
						end
						2'd2, 2'd3: begin
							// Trace: design.sv:43330:15
							accum_window_d = {next_remainder[31:0], op_numerator_q[multdiv_count_d]};
							// Trace: design.sv:43331:15
							op_a_shift_d = next_quotient;
							// Trace: design.sv:43332:15
							md_state_d = (multdiv_count_q == 5'd1 ? 3'd4 : 3'd3);
						end
						default:
							;
					endcase
				end
				3'd4:
					// Trace: design.sv:43339:11
					(* full_case, parallel_case *)
					case (operator_i)
						2'd0: begin
							// Trace: design.sv:43341:15
							accum_window_d = res_adder_l;
							// Trace: design.sv:43344:15
							md_state_d = 3'd0;
							// Trace: design.sv:43345:15
							multdiv_hold = ~multdiv_ready_id_i;
						end
						2'd1: begin
							// Trace: design.sv:43348:15
							accum_window_d = res_adder_l;
							// Trace: design.sv:43349:15
							md_state_d = 3'd0;
							// Trace: design.sv:43352:15
							md_state_d = 3'd0;
							// Trace: design.sv:43353:15
							multdiv_hold = ~multdiv_ready_id_i;
						end
						2'd2: begin
							// Trace: design.sv:43358:15
							accum_window_d = next_quotient;
							// Trace: design.sv:43359:15
							md_state_d = 3'd5;
						end
						2'd3: begin
							// Trace: design.sv:43363:15
							accum_window_d = {1'b0, next_remainder[31:0]};
							// Trace: design.sv:43364:15
							md_state_d = 3'd5;
						end
						default:
							;
					endcase
				3'd5: begin
					// Trace: design.sv:43371:11
					md_state_d = 3'd6;
					// Trace: design.sv:43372:11
					(* full_case, parallel_case *)
					case (operator_i)
						2'd2:
							// Trace: design.sv:43374:15
							accum_window_d = (div_change_sign ? {1'b0, alu_adder_i} : accum_window_q);
						2'd3:
							// Trace: design.sv:43376:15
							accum_window_d = (rem_change_sign ? {1'b0, alu_adder_i} : accum_window_q);
						default:
							;
					endcase
				end
				3'd6: begin
					// Trace: design.sv:43383:11
					md_state_d = 3'd0;
					// Trace: design.sv:43384:11
					multdiv_hold = ~multdiv_ready_id_i;
				end
				default:
					// Trace: design.sv:43388:11
					md_state_d = 3'd0;
			endcase
	end
	// Trace: design.sv:43398:3
	assign multdiv_en = (mult_en_i | div_en_i) & ~multdiv_hold;
	// Trace: design.sv:43400:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:43401:5
		if (!rst_ni) begin
			// Trace: design.sv:43402:7
			multdiv_count_q <= 5'h00;
			// Trace: design.sv:43403:7
			op_b_shift_q <= 33'h000000000;
			// Trace: design.sv:43404:7
			op_a_shift_q <= 33'h000000000;
			// Trace: design.sv:43405:7
			md_state_q <= 3'd0;
			// Trace: design.sv:43406:7
			div_by_zero_q <= 1'b0;
		end
		else if (multdiv_en) begin
			// Trace: design.sv:43408:7
			multdiv_count_q <= multdiv_count_d;
			// Trace: design.sv:43409:7
			op_b_shift_q <= op_b_shift_d;
			// Trace: design.sv:43410:7
			op_a_shift_q <= op_a_shift_d;
			// Trace: design.sv:43411:7
			md_state_q <= md_state_d;
			// Trace: design.sv:43412:7
			div_by_zero_q <= div_by_zero_d;
		end
	// Trace: design.sv:43420:3
	assign valid_o = (md_state_q == 3'd6) | ((md_state_q == 3'd4) & ((operator_i == 2'd0) | (operator_i == 2'd1)));
	// Trace: design.sv:43425:3
	assign multdiv_result_o = (div_en_i ? accum_window_q[31:0] : res_adder_l[31:0]);
	initial _sv2v_0 = 0;
endmodule
module ibex_prefetch_buffer (
	clk_i,
	rst_ni,
	req_i,
	branch_i,
	branch_mispredict_i,
	mispredict_addr_i,
	addr_i,
	ready_i,
	valid_o,
	rdata_o,
	addr_o,
	err_o,
	err_plus2_o,
	instr_req_o,
	instr_gnt_i,
	instr_addr_o,
	instr_rdata_i,
	instr_err_i,
	instr_rvalid_i,
	busy_o
);
	// Trace: design.sv:43455:13
	parameter [0:0] ResetAll = 1'b0;
	// Trace: design.sv:43457:3
	input wire clk_i;
	// Trace: design.sv:43458:3
	input wire rst_ni;
	// Trace: design.sv:43460:3
	input wire req_i;
	// Trace: design.sv:43462:3
	input wire branch_i;
	// Trace: design.sv:43463:3
	input wire branch_mispredict_i;
	// Trace: design.sv:43464:3
	input wire [31:0] mispredict_addr_i;
	// Trace: design.sv:43465:3
	input wire [31:0] addr_i;
	// Trace: design.sv:43468:3
	input wire ready_i;
	// Trace: design.sv:43469:3
	output wire valid_o;
	// Trace: design.sv:43470:3
	output wire [31:0] rdata_o;
	// Trace: design.sv:43471:3
	output wire [31:0] addr_o;
	// Trace: design.sv:43472:3
	output wire err_o;
	// Trace: design.sv:43473:3
	output wire err_plus2_o;
	// Trace: design.sv:43476:3
	output wire instr_req_o;
	// Trace: design.sv:43477:3
	input wire instr_gnt_i;
	// Trace: design.sv:43478:3
	output wire [31:0] instr_addr_o;
	// Trace: design.sv:43479:3
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:43480:3
	input wire instr_err_i;
	// Trace: design.sv:43481:3
	input wire instr_rvalid_i;
	// Trace: design.sv:43484:3
	output wire busy_o;
	// Trace: design.sv:43487:3
	localparam [31:0] NUM_REQS = 2;
	// Trace: design.sv:43489:3
	wire valid_new_req;
	wire valid_req;
	// Trace: design.sv:43490:3
	wire valid_req_d;
	reg valid_req_q;
	// Trace: design.sv:43491:3
	wire discard_req_d;
	reg discard_req_q;
	// Trace: design.sv:43492:3
	wire [1:0] rdata_outstanding_n;
	wire [1:0] rdata_outstanding_s;
	reg [1:0] rdata_outstanding_q;
	// Trace: design.sv:43493:3
	wire [1:0] branch_discard_n;
	wire [1:0] branch_discard_s;
	reg [1:0] branch_discard_q;
	// Trace: design.sv:43494:3
	wire [1:0] rdata_outstanding_rev;
	// Trace: design.sv:43496:3
	wire [31:0] stored_addr_d;
	reg [31:0] stored_addr_q;
	// Trace: design.sv:43497:3
	wire stored_addr_en;
	// Trace: design.sv:43498:3
	wire [31:0] fetch_addr_d;
	reg [31:0] fetch_addr_q;
	// Trace: design.sv:43499:3
	wire fetch_addr_en;
	// Trace: design.sv:43500:3
	wire [31:0] instr_addr;
	wire [31:0] instr_addr_w_aligned;
	// Trace: design.sv:43502:3
	wire fifo_valid;
	// Trace: design.sv:43503:3
	wire [31:0] fifo_addr;
	// Trace: design.sv:43504:3
	wire fifo_ready;
	// Trace: design.sv:43505:3
	wire fifo_clear;
	// Trace: design.sv:43506:3
	wire [1:0] fifo_busy;
	// Trace: design.sv:43508:3
	wire valid_raw;
	// Trace: design.sv:43510:3
	wire branch_or_mispredict;
	// Trace: design.sv:43516:3
	assign busy_o = |rdata_outstanding_q | instr_req_o;
	// Trace: design.sv:43518:3
	assign branch_or_mispredict = branch_i | branch_mispredict_i;
	// Trace: design.sv:43527:3
	assign fifo_clear = branch_or_mispredict;
	// Trace: design.sv:43530:3
	genvar _gv_i_67;
	generate
		for (_gv_i_67 = 0; _gv_i_67 < NUM_REQS; _gv_i_67 = _gv_i_67 + 1) begin : gen_rd_rev
			localparam i = _gv_i_67;
			// Trace: design.sv:43531:5
			assign rdata_outstanding_rev[i] = rdata_outstanding_q[1 - i];
		end
	endgenerate
	// Trace: design.sv:43537:3
	assign fifo_ready = ~&(fifo_busy | rdata_outstanding_rev);
	// Trace: design.sv:43539:3
	ibex_fetch_fifo #(
		.NUM_REQS(NUM_REQS),
		.ResetAll(ResetAll)
	) fifo_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clear_i(fifo_clear),
		.busy_o(fifo_busy),
		.in_valid_i(fifo_valid),
		.in_addr_i(fifo_addr),
		.in_rdata_i(instr_rdata_i),
		.in_err_i(instr_err_i),
		.out_valid_o(valid_raw),
		.out_ready_i(ready_i),
		.out_rdata_o(rdata_o),
		.out_addr_o(addr_o),
		.out_err_o(err_o),
		.out_err_plus2_o(err_plus2_o)
	);
	// Trace: design.sv:43567:3
	assign valid_new_req = (req_i & (fifo_ready | branch_or_mispredict)) & ~rdata_outstanding_q[1];
	// Trace: design.sv:43570:3
	assign valid_req = valid_req_q | valid_new_req;
	// Trace: design.sv:43573:3
	assign valid_req_d = valid_req & ~instr_gnt_i;
	// Trace: design.sv:43576:3
	assign discard_req_d = valid_req_q & (branch_or_mispredict | discard_req_q);
	// Trace: design.sv:43595:3
	assign stored_addr_en = (valid_new_req & ~valid_req_q) & ~instr_gnt_i;
	// Trace: design.sv:43598:3
	assign stored_addr_d = instr_addr;
	// Trace: design.sv:43601:3
	generate
		if (ResetAll) begin : g_stored_addr_ra
			// Trace: design.sv:43602:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:43603:7
				if (!rst_ni)
					// Trace: design.sv:43604:9
					stored_addr_q <= 1'sb0;
				else if (stored_addr_en)
					// Trace: design.sv:43606:9
					stored_addr_q <= stored_addr_d;
		end
		else begin : g_stored_addr_nr
			// Trace: design.sv:43610:5
			always @(posedge clk_i)
				// Trace: design.sv:43611:7
				if (stored_addr_en)
					// Trace: design.sv:43612:9
					stored_addr_q <= stored_addr_d;
		end
	endgenerate
	// Trace: design.sv:43619:3
	assign fetch_addr_en = branch_or_mispredict | (valid_new_req & ~valid_req_q);
	// Trace: design.sv:43621:3
	assign fetch_addr_d = (branch_i ? addr_i : (branch_mispredict_i ? {mispredict_addr_i[31:2], 2'b00} : {fetch_addr_q[31:2], 2'b00})) + {{29 {1'b0}}, valid_new_req & ~valid_req_q, 2'b00};
	// Trace: design.sv:43627:3
	generate
		if (ResetAll) begin : g_fetch_addr_ra
			// Trace: design.sv:43628:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:43629:7
				if (!rst_ni)
					// Trace: design.sv:43630:9
					fetch_addr_q <= 1'sb0;
				else if (fetch_addr_en)
					// Trace: design.sv:43632:9
					fetch_addr_q <= fetch_addr_d;
		end
		else begin : g_fetch_addr_nr
			// Trace: design.sv:43636:5
			always @(posedge clk_i)
				// Trace: design.sv:43637:7
				if (fetch_addr_en)
					// Trace: design.sv:43638:9
					fetch_addr_q <= fetch_addr_d;
		end
	endgenerate
	// Trace: design.sv:43644:3
	assign instr_addr = (valid_req_q ? stored_addr_q : (branch_i ? addr_i : (branch_mispredict_i ? mispredict_addr_i : fetch_addr_q)));
	// Trace: design.sv:43649:3
	assign instr_addr_w_aligned = {instr_addr[31:2], 2'b00};
	// Trace: design.sv:43655:3
	genvar _gv_i_68;
	generate
		for (_gv_i_68 = 0; _gv_i_68 < NUM_REQS; _gv_i_68 = _gv_i_68 + 1) begin : g_outstanding_reqs
			localparam i = _gv_i_68;
			if (i == 0) begin : g_req0
				// Trace: design.sv:43660:7
				assign rdata_outstanding_n[i] = (valid_req & instr_gnt_i) | rdata_outstanding_q[i];
				// Trace: design.sv:43664:7
				assign branch_discard_n[i] = (((valid_req & instr_gnt_i) & discard_req_d) | (branch_or_mispredict & rdata_outstanding_q[i])) | branch_discard_q[i];
			end
			else begin : g_reqtop
				// Trace: design.sv:43672:7
				assign rdata_outstanding_n[i] = ((valid_req & instr_gnt_i) & rdata_outstanding_q[i - 1]) | rdata_outstanding_q[i];
				// Trace: design.sv:43675:7
				assign branch_discard_n[i] = ((((valid_req & instr_gnt_i) & discard_req_d) & rdata_outstanding_q[i - 1]) | (branch_or_mispredict & rdata_outstanding_q[i])) | branch_discard_q[i];
			end
		end
	endgenerate
	// Trace: design.sv:43683:3
	assign rdata_outstanding_s = (instr_rvalid_i ? {1'b0, rdata_outstanding_n[1:1]} : rdata_outstanding_n);
	// Trace: design.sv:43685:3
	assign branch_discard_s = (instr_rvalid_i ? {1'b0, branch_discard_n[1:1]} : branch_discard_n);
	// Trace: design.sv:43689:3
	assign fifo_valid = instr_rvalid_i & ~branch_discard_q[0];
	// Trace: design.sv:43691:3
	assign fifo_addr = (branch_i ? addr_i : mispredict_addr_i);
	// Trace: design.sv:43697:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:43698:5
		if (!rst_ni) begin
			// Trace: design.sv:43699:7
			valid_req_q <= 1'b0;
			// Trace: design.sv:43700:7
			discard_req_q <= 1'b0;
			// Trace: design.sv:43701:7
			rdata_outstanding_q <= 'b0;
			// Trace: design.sv:43702:7
			branch_discard_q <= 'b0;
		end
		else begin
			// Trace: design.sv:43704:7
			valid_req_q <= valid_req_d;
			// Trace: design.sv:43705:7
			discard_req_q <= discard_req_d;
			// Trace: design.sv:43706:7
			rdata_outstanding_q <= rdata_outstanding_s;
			// Trace: design.sv:43707:7
			branch_discard_q <= branch_discard_s;
		end
	// Trace: design.sv:43715:3
	assign instr_req_o = valid_req;
	// Trace: design.sv:43716:3
	assign instr_addr_o = instr_addr_w_aligned;
	// Trace: design.sv:43718:3
	assign valid_o = valid_raw & ~branch_mispredict_i;
endmodule
module ibex_pmp (
	clk_i,
	rst_ni,
	csr_pmp_cfg_i,
	csr_pmp_addr_i,
	csr_pmp_mseccfg_i,
	priv_mode_i,
	pmp_req_addr_i,
	pmp_req_type_i,
	pmp_req_err_o
);
	reg _sv2v_0;
	// Trace: design.sv:43728:13
	parameter [31:0] PMPGranularity = 0;
	// Trace: design.sv:43730:13
	parameter [31:0] PMPNumChan = 2;
	// Trace: design.sv:43732:13
	parameter [31:0] PMPNumRegions = 4;
	// Trace: design.sv:43735:3
	input wire clk_i;
	// Trace: design.sv:43736:3
	input wire rst_ni;
	// Trace: design.sv:43739:3
	// removed localparam type ibex_pkg_pmp_cfg_mode_e
	// removed localparam type ibex_pkg_pmp_cfg_t
	input wire [(PMPNumRegions * 6) - 1:0] csr_pmp_cfg_i;
	// Trace: design.sv:43740:3
	input wire [(PMPNumRegions * 34) - 1:0] csr_pmp_addr_i;
	// Trace: design.sv:43741:3
	// removed localparam type ibex_pkg_pmp_mseccfg_t
	input wire [2:0] csr_pmp_mseccfg_i;
	// Trace: design.sv:43743:3
	// removed localparam type ibex_pkg_priv_lvl_e
	input wire [(PMPNumChan * 2) - 1:0] priv_mode_i;
	// Trace: design.sv:43745:3
	input wire [(PMPNumChan * 34) - 1:0] pmp_req_addr_i;
	// Trace: design.sv:43746:3
	// removed localparam type ibex_pkg_pmp_req_e
	input wire [(PMPNumChan * 2) - 1:0] pmp_req_type_i;
	// Trace: design.sv:43747:3
	output wire [0:PMPNumChan - 1] pmp_req_err_o;
	// Trace: design.sv:43751:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:43754:3
	wire [33:0] region_start_addr [0:PMPNumRegions - 1];
	// Trace: design.sv:43755:3
	wire [33:PMPGranularity + 2] region_addr_mask [0:PMPNumRegions - 1];
	// Trace: design.sv:43756:3
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_match_gt;
	// Trace: design.sv:43757:3
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_match_lt;
	// Trace: design.sv:43758:3
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_match_eq;
	// Trace: design.sv:43759:3
	reg [(PMPNumChan * PMPNumRegions) - 1:0] region_match_all;
	// Trace: design.sv:43760:3
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_basic_perm_check;
	// Trace: design.sv:43761:3
	reg [(PMPNumChan * PMPNumRegions) - 1:0] region_mml_perm_check;
	// Trace: design.sv:43762:3
	reg [PMPNumChan - 1:0] access_fault;
	// Trace: design.sv:43769:3
	genvar _gv_r_3;
	generate
		for (_gv_r_3 = 0; _gv_r_3 < PMPNumRegions; _gv_r_3 = _gv_r_3 + 1) begin : g_addr_exp
			localparam r = _gv_r_3;
			if (r == 0) begin : g_entry0
				// Trace: design.sv:43772:7
				assign region_start_addr[r] = (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] == 2'b01 ? 34'h000000000 : csr_pmp_addr_i[((PMPNumRegions - 1) - r) * 34+:34]);
			end
			else begin : g_oth
				// Trace: design.sv:43775:7
				assign region_start_addr[r] = (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] == 2'b01 ? csr_pmp_addr_i[((PMPNumRegions - 1) - (r - 1)) * 34+:34] : csr_pmp_addr_i[((PMPNumRegions - 1) - r) * 34+:34]);
			end
			genvar _gv_b_1;
			for (_gv_b_1 = PMPGranularity + 2; _gv_b_1 < 34; _gv_b_1 = _gv_b_1 + 1) begin : g_bitmask
				localparam b = _gv_b_1;
				if (b == 2) begin : g_bit0
					// Trace: design.sv:43782:9
					assign region_addr_mask[r][b] = csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] != 2'b11;
				end
				else begin : g_others
					if (PMPGranularity == 0) begin : g_region_addr_mask_zero_granularity
						// Trace: design.sv:43790:11
						assign region_addr_mask[r][b] = (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] != 2'b11) | ~&csr_pmp_addr_i[(((PMPNumRegions - 1) - r) * 34) + ((b - 1) >= 2 ? b - 1 : ((b - 1) + ((b - 1) >= 2 ? b - 2 : 4 - b)) - 1)-:((b - 1) >= 2 ? b - 2 : 4 - b)];
					end
					else begin : g_region_addr_mask_other_granularity
						// Trace: design.sv:43793:11
						assign region_addr_mask[r][b] = (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] != 2'b11) | ~&csr_pmp_addr_i[(((PMPNumRegions - 1) - r) * 34) + ((b - 1) >= (PMPGranularity + 1) ? b - 1 : ((b - 1) + ((b - 1) >= (PMPGranularity + 1) ? ((b - 1) - (PMPGranularity + 1)) + 1 : ((PMPGranularity + 1) - (b - 1)) + 1)) - 1)-:((b - 1) >= (PMPGranularity + 1) ? ((b - 1) - (PMPGranularity + 1)) + 1 : ((PMPGranularity + 1) - (b - 1)) + 1)];
					end
				end
			end
		end
	endgenerate
	// Trace: design.sv:43800:3
	genvar _gv_c_1;
	generate
		for (_gv_c_1 = 0; _gv_c_1 < PMPNumChan; _gv_c_1 = _gv_c_1 + 1) begin : g_access_check
			localparam c = _gv_c_1;
			genvar _gv_r_4;
			for (_gv_r_4 = 0; _gv_r_4 < PMPNumRegions; _gv_r_4 = _gv_r_4 + 1) begin : g_regions
				localparam r = _gv_r_4;
				// Trace: design.sv:43803:7
				assign region_match_eq[(c * PMPNumRegions) + r] = (pmp_req_addr_i[(((PMPNumChan - 1) - c) * 34) + (33 >= (PMPGranularity + 2) ? 33 : (33 + (33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)) - 1)-:(33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)] & region_addr_mask[r]) == (region_start_addr[r][33:PMPGranularity + 2] & region_addr_mask[r]);
				// Trace: design.sv:43807:7
				assign region_match_gt[(c * PMPNumRegions) + r] = pmp_req_addr_i[(((PMPNumChan - 1) - c) * 34) + (33 >= (PMPGranularity + 2) ? 33 : (33 + (33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)) - 1)-:(33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)] > region_start_addr[r][33:PMPGranularity + 2];
				// Trace: design.sv:43809:7
				assign region_match_lt[(c * PMPNumRegions) + r] = pmp_req_addr_i[(((PMPNumChan - 1) - c) * 34) + (33 >= (PMPGranularity + 2) ? 33 : (33 + (33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)) - 1)-:(33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)] < csr_pmp_addr_i[(((PMPNumRegions - 1) - r) * 34) + (33 >= (PMPGranularity + 2) ? 33 : (33 + (33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)) - 1)-:(33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)];
				// Trace: design.sv:43812:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:43813:9
					region_match_all[(c * PMPNumRegions) + r] = 1'b0;
					// Trace: design.sv:43814:9
					(* full_case, parallel_case *)
					case (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2])
						2'b00:
							// Trace: design.sv:43815:27
							region_match_all[(c * PMPNumRegions) + r] = 1'b0;
						2'b10:
							// Trace: design.sv:43816:27
							region_match_all[(c * PMPNumRegions) + r] = region_match_eq[(c * PMPNumRegions) + r];
						2'b11:
							// Trace: design.sv:43817:27
							region_match_all[(c * PMPNumRegions) + r] = region_match_eq[(c * PMPNumRegions) + r];
						2'b01:
							// Trace: design.sv:43819:13
							region_match_all[(c * PMPNumRegions) + r] = (region_match_eq[(c * PMPNumRegions) + r] | region_match_gt[(c * PMPNumRegions) + r]) & region_match_lt[(c * PMPNumRegions) + r];
						default:
							// Trace: design.sv:43822:27
							region_match_all[(c * PMPNumRegions) + r] = 1'b0;
					endcase
				end
				// Trace: design.sv:43827:7
				assign region_basic_perm_check[(c * PMPNumRegions) + r] = (((pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b00) & csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 2]) | ((pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b01) & csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 1])) | ((pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b10) & csr_pmp_cfg_i[((PMPNumRegions - 1) - r) * 6]);
				// Trace: design.sv:43834:7
				always @(*) begin
					if (_sv2v_0)
						;
					// Trace: design.sv:43835:9
					region_mml_perm_check[(c * PMPNumRegions) + r] = 1'b0;
					// Trace: design.sv:43837:9
					if (!csr_pmp_cfg_i[((PMPNumRegions - 1) - r) * 6] && csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 1])
						// Trace: design.sv:43839:11
						(* full_case, parallel_case *)
						case ({csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 5], csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 2]})
							2'b00:
								// Trace: design.sv:43841:20
								region_mml_perm_check[(c * PMPNumRegions) + r] = (pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b10) | ((pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b01) & (priv_mode_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b11));
							2'b01:
								// Trace: design.sv:43845:20
								region_mml_perm_check[(c * PMPNumRegions) + r] = (pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b10) | (pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b01);
							2'b10:
								// Trace: design.sv:43848:20
								region_mml_perm_check[(c * PMPNumRegions) + r] = pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b00;
							2'b11:
								// Trace: design.sv:43850:20
								region_mml_perm_check[(c * PMPNumRegions) + r] = (pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b00) | ((pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b10) & (priv_mode_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b11));
							default:
								;
						endcase
					else
						// Trace: design.sv:43856:11
						if (((csr_pmp_cfg_i[((PMPNumRegions - 1) - r) * 6] & csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 1]) & csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 2]) & csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 5])
							// Trace: design.sv:43859:13
							region_mml_perm_check[(c * PMPNumRegions) + r] = pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b10;
						else
							// Trace: design.sv:43863:13
							region_mml_perm_check[(c * PMPNumRegions) + r] = (priv_mode_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b11 ? csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 5] & region_basic_perm_check[(c * PMPNumRegions) + r] : ~csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 5] & region_basic_perm_check[(c * PMPNumRegions) + r]);
				end
			end
			// Trace: design.sv:43872:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:43875:7
				access_fault[c] = csr_pmp_mseccfg_i[1] | (priv_mode_i[((PMPNumChan - 1) - c) * 2+:2] != 2'b11);
				// Trace: design.sv:43879:7
				begin : sv2v_autoblock_1
					// Trace: design.sv:43879:12
					reg signed [31:0] r;
					// Trace: design.sv:43879:12
					for (r = PMPNumRegions - 1; r >= 0; r = r - 1)
						begin
							// Trace: design.sv:43880:9
							if (region_match_all[(c * PMPNumRegions) + r]) begin
								begin
									// Trace: design.sv:43881:11
									if (csr_pmp_mseccfg_i[0])
										// Trace: design.sv:43883:13
										access_fault[c] = ~region_mml_perm_check[(c * PMPNumRegions) + r];
									else
										// Trace: design.sv:43886:13
										access_fault[c] = (priv_mode_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b11 ? csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 5] & ~region_basic_perm_check[(c * PMPNumRegions) + r] : ~region_basic_perm_check[(c * PMPNumRegions) + r]);
								end
							end
						end
				end
			end
			// Trace: design.sv:43897:5
			assign pmp_req_err_o[c] = access_fault[c];
		end
	endgenerate
	// Trace: design.sv:43902:3
	wire unused_csr_pmp_mseccfg_rlb;
	// Trace: design.sv:43903:3
	assign unused_csr_pmp_mseccfg_rlb = csr_pmp_mseccfg_i[2];
	initial _sv2v_0 = 0;
endmodule
module ibex_wb_stage (
	clk_i,
	rst_ni,
	en_wb_i,
	instr_type_wb_i,
	pc_id_i,
	instr_is_compressed_id_i,
	instr_perf_count_id_i,
	ready_wb_o,
	rf_write_wb_o,
	outstanding_load_wb_o,
	outstanding_store_wb_o,
	pc_wb_o,
	perf_instr_ret_wb_o,
	perf_instr_ret_compressed_wb_o,
	perf_instr_ret_wb_spec_o,
	perf_instr_ret_compressed_wb_spec_o,
	rf_waddr_id_i,
	rf_wdata_id_i,
	rf_we_id_i,
	rf_wdata_lsu_i,
	rf_we_lsu_i,
	rf_wdata_fwd_wb_o,
	rf_waddr_wb_o,
	rf_wdata_wb_o,
	rf_we_wb_o,
	lsu_resp_valid_i,
	lsu_resp_err_i,
	instr_done_wb_o
);
	// Trace: design.sv:43922:13
	parameter [0:0] ResetAll = 1'b0;
	// Trace: design.sv:43923:13
	parameter [0:0] WritebackStage = 1'b0;
	// Trace: design.sv:43925:3
	input wire clk_i;
	// Trace: design.sv:43926:3
	input wire rst_ni;
	// Trace: design.sv:43928:3
	input wire en_wb_i;
	// Trace: design.sv:43929:3
	// removed localparam type ibex_pkg_wb_instr_type_e
	input wire [1:0] instr_type_wb_i;
	// Trace: design.sv:43930:3
	input wire [31:0] pc_id_i;
	// Trace: design.sv:43931:3
	input wire instr_is_compressed_id_i;
	// Trace: design.sv:43932:3
	input wire instr_perf_count_id_i;
	// Trace: design.sv:43934:3
	output wire ready_wb_o;
	// Trace: design.sv:43935:3
	output wire rf_write_wb_o;
	// Trace: design.sv:43936:3
	output wire outstanding_load_wb_o;
	// Trace: design.sv:43937:3
	output wire outstanding_store_wb_o;
	// Trace: design.sv:43938:3
	output wire [31:0] pc_wb_o;
	// Trace: design.sv:43939:3
	output wire perf_instr_ret_wb_o;
	// Trace: design.sv:43940:3
	output wire perf_instr_ret_compressed_wb_o;
	// Trace: design.sv:43941:3
	output wire perf_instr_ret_wb_spec_o;
	// Trace: design.sv:43942:3
	output wire perf_instr_ret_compressed_wb_spec_o;
	// Trace: design.sv:43944:3
	input wire [4:0] rf_waddr_id_i;
	// Trace: design.sv:43945:3
	input wire [31:0] rf_wdata_id_i;
	// Trace: design.sv:43946:3
	input wire rf_we_id_i;
	// Trace: design.sv:43948:3
	input wire [31:0] rf_wdata_lsu_i;
	// Trace: design.sv:43949:3
	input wire rf_we_lsu_i;
	// Trace: design.sv:43951:3
	output wire [31:0] rf_wdata_fwd_wb_o;
	// Trace: design.sv:43953:3
	output wire [4:0] rf_waddr_wb_o;
	// Trace: design.sv:43954:3
	output wire [31:0] rf_wdata_wb_o;
	// Trace: design.sv:43955:3
	output wire rf_we_wb_o;
	// Trace: design.sv:43957:3
	input wire lsu_resp_valid_i;
	// Trace: design.sv:43958:3
	input wire lsu_resp_err_i;
	// Trace: design.sv:43960:3
	output wire instr_done_wb_o;
	// Trace: design.sv:43963:3
	// removed import ibex_pkg::*;
	// Trace: design.sv:43967:3
	wire [31:0] rf_wdata_wb_mux [0:1];
	// Trace: design.sv:43968:3
	wire [1:0] rf_wdata_wb_mux_we;
	// Trace: design.sv:43970:3
	generate
		if (WritebackStage) begin : g_writeback_stage
			// Trace: design.sv:43971:5
			reg [31:0] rf_wdata_wb_q;
			// Trace: design.sv:43972:5
			reg rf_we_wb_q;
			// Trace: design.sv:43973:5
			reg [4:0] rf_waddr_wb_q;
			// Trace: design.sv:43975:5
			wire wb_done;
			// Trace: design.sv:43977:5
			reg wb_valid_q;
			// Trace: design.sv:43978:5
			reg [31:0] wb_pc_q;
			// Trace: design.sv:43979:5
			reg wb_compressed_q;
			// Trace: design.sv:43980:5
			reg wb_count_q;
			// Trace: design.sv:43981:5
			reg [1:0] wb_instr_type_q;
			// Trace: design.sv:43983:5
			wire wb_valid_d;
			// Trace: design.sv:43987:5
			assign wb_valid_d = (en_wb_i & ready_wb_o) | (wb_valid_q & ~wb_done);
			// Trace: design.sv:43992:5
			assign wb_done = (wb_instr_type_q == 2'd2) | lsu_resp_valid_i;
			// Trace: design.sv:43994:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:43995:7
				if (!rst_ni)
					// Trace: design.sv:43996:9
					wb_valid_q <= 1'b0;
				else
					// Trace: design.sv:43998:9
					wb_valid_q <= wb_valid_d;
			if (ResetAll) begin : g_wb_regs_ra
				// Trace: design.sv:44003:7
				always @(posedge clk_i or negedge rst_ni)
					// Trace: design.sv:44004:9
					if (!rst_ni) begin
						// Trace: design.sv:44005:11
						rf_we_wb_q <= 1'sb0;
						// Trace: design.sv:44006:11
						rf_waddr_wb_q <= 1'sb0;
						// Trace: design.sv:44007:11
						rf_wdata_wb_q <= 1'sb0;
						// Trace: design.sv:44008:11
						wb_instr_type_q <= 2'd0;
						// Trace: design.sv:44009:11
						wb_pc_q <= 1'sb0;
						// Trace: design.sv:44010:11
						wb_compressed_q <= 1'sb0;
						// Trace: design.sv:44011:11
						wb_count_q <= 1'sb0;
					end
					else if (en_wb_i) begin
						// Trace: design.sv:44013:11
						rf_we_wb_q <= rf_we_id_i;
						// Trace: design.sv:44014:11
						rf_waddr_wb_q <= rf_waddr_id_i;
						// Trace: design.sv:44015:11
						rf_wdata_wb_q <= rf_wdata_id_i;
						// Trace: design.sv:44016:11
						wb_instr_type_q <= instr_type_wb_i;
						// Trace: design.sv:44017:11
						wb_pc_q <= pc_id_i;
						// Trace: design.sv:44018:11
						wb_compressed_q <= instr_is_compressed_id_i;
						// Trace: design.sv:44019:11
						wb_count_q <= instr_perf_count_id_i;
					end
			end
			else begin : g_wb_regs_nr
				// Trace: design.sv:44023:7
				always @(posedge clk_i)
					// Trace: design.sv:44024:9
					if (en_wb_i) begin
						// Trace: design.sv:44025:11
						rf_we_wb_q <= rf_we_id_i;
						// Trace: design.sv:44026:11
						rf_waddr_wb_q <= rf_waddr_id_i;
						// Trace: design.sv:44027:11
						rf_wdata_wb_q <= rf_wdata_id_i;
						// Trace: design.sv:44028:11
						wb_instr_type_q <= instr_type_wb_i;
						// Trace: design.sv:44029:11
						wb_pc_q <= pc_id_i;
						// Trace: design.sv:44030:11
						wb_compressed_q <= instr_is_compressed_id_i;
						// Trace: design.sv:44031:11
						wb_count_q <= instr_perf_count_id_i;
					end
			end
			// Trace: design.sv:44036:5
			assign rf_waddr_wb_o = rf_waddr_wb_q;
			// Trace: design.sv:44037:5
			assign rf_wdata_wb_mux[0] = rf_wdata_wb_q;
			// Trace: design.sv:44038:5
			assign rf_wdata_wb_mux_we[0] = rf_we_wb_q & wb_valid_q;
			// Trace: design.sv:44040:5
			assign ready_wb_o = ~wb_valid_q | wb_done;
			// Trace: design.sv:44044:5
			assign rf_write_wb_o = wb_valid_q & (rf_we_wb_q | (wb_instr_type_q == 2'd0));
			// Trace: design.sv:44046:5
			assign outstanding_load_wb_o = wb_valid_q & (wb_instr_type_q == 2'd0);
			// Trace: design.sv:44047:5
			assign outstanding_store_wb_o = wb_valid_q & (wb_instr_type_q == 2'd1);
			// Trace: design.sv:44049:5
			assign pc_wb_o = wb_pc_q;
			// Trace: design.sv:44051:5
			assign instr_done_wb_o = wb_valid_q & wb_done;
			// Trace: design.sv:44057:5
			assign perf_instr_ret_wb_spec_o = wb_count_q;
			// Trace: design.sv:44058:5
			assign perf_instr_ret_compressed_wb_spec_o = perf_instr_ret_wb_spec_o & wb_compressed_q;
			// Trace: design.sv:44059:5
			assign perf_instr_ret_wb_o = (instr_done_wb_o & wb_count_q) & ~(lsu_resp_valid_i & lsu_resp_err_i);
			// Trace: design.sv:44061:5
			assign perf_instr_ret_compressed_wb_o = perf_instr_ret_wb_o & wb_compressed_q;
			// Trace: design.sv:44066:5
			assign rf_wdata_fwd_wb_o = rf_wdata_wb_q;
		end
		else begin : g_bypass_wb
			// Trace: design.sv:44069:5
			assign rf_waddr_wb_o = rf_waddr_id_i;
			// Trace: design.sv:44070:5
			assign rf_wdata_wb_mux[0] = rf_wdata_id_i;
			// Trace: design.sv:44071:5
			assign rf_wdata_wb_mux_we[0] = rf_we_id_i;
			// Trace: design.sv:44076:5
			assign perf_instr_ret_wb_spec_o = 1'b0;
			// Trace: design.sv:44077:5
			assign perf_instr_ret_compressed_wb_spec_o = 1'b0;
			// Trace: design.sv:44078:5
			assign perf_instr_ret_wb_o = (instr_perf_count_id_i & en_wb_i) & ~(lsu_resp_valid_i & lsu_resp_err_i);
			// Trace: design.sv:44080:5
			assign perf_instr_ret_compressed_wb_o = perf_instr_ret_wb_o & instr_is_compressed_id_i;
			// Trace: design.sv:44083:5
			assign ready_wb_o = 1'b1;
			// Trace: design.sv:44088:5
			wire unused_clk;
			// Trace: design.sv:44089:5
			wire unused_rst;
			// Trace: design.sv:44090:5
			wire [1:0] unused_instr_type_wb;
			// Trace: design.sv:44091:5
			wire [31:0] unused_pc_id;
			// Trace: design.sv:44093:5
			assign unused_clk = clk_i;
			// Trace: design.sv:44094:5
			assign unused_rst = rst_ni;
			// Trace: design.sv:44095:5
			assign unused_instr_type_wb = instr_type_wb_i;
			// Trace: design.sv:44096:5
			assign unused_pc_id = pc_id_i;
			// Trace: design.sv:44098:5
			assign outstanding_load_wb_o = 1'b0;
			// Trace: design.sv:44099:5
			assign outstanding_store_wb_o = 1'b0;
			// Trace: design.sv:44100:5
			assign pc_wb_o = 1'sb0;
			// Trace: design.sv:44101:5
			assign rf_write_wb_o = 1'b0;
			// Trace: design.sv:44102:5
			assign rf_wdata_fwd_wb_o = 32'b00000000000000000000000000000000;
			// Trace: design.sv:44103:5
			assign instr_done_wb_o = 1'b0;
		end
	endgenerate
	// Trace: design.sv:44106:3
	assign rf_wdata_wb_mux[1] = rf_wdata_lsu_i;
	// Trace: design.sv:44107:3
	assign rf_wdata_wb_mux_we[1] = rf_we_lsu_i;
	// Trace: design.sv:44111:3
	assign rf_wdata_wb_o = ({32 {rf_wdata_wb_mux_we[0]}} & rf_wdata_wb_mux[0]) | ({32 {rf_wdata_wb_mux_we[1]}} & rf_wdata_wb_mux[1]);
	// Trace: design.sv:44113:3
	assign rf_we_wb_o = |rf_wdata_wb_mux_we;
endmodule
module ibex_dummy_instr (
	clk_i,
	rst_ni,
	dummy_instr_en_i,
	dummy_instr_mask_i,
	dummy_instr_seed_en_i,
	dummy_instr_seed_i,
	fetch_valid_i,
	id_in_ready_i,
	insert_dummy_instr_o,
	dummy_instr_data_o
);
	reg _sv2v_0;
	// removed import ibex_pkg::*;
	// Trace: design.sv:44131:15
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	// removed localparam type ibex_pkg_lfsr_seed_t
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	// Trace: design.sv:44132:15
	// removed localparam type ibex_pkg_lfsr_perm_t
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	// Trace: design.sv:44135:3
	input wire clk_i;
	// Trace: design.sv:44136:3
	input wire rst_ni;
	// Trace: design.sv:44139:3
	input wire dummy_instr_en_i;
	// Trace: design.sv:44140:3
	input wire [2:0] dummy_instr_mask_i;
	// Trace: design.sv:44141:3
	input wire dummy_instr_seed_en_i;
	// Trace: design.sv:44142:3
	input wire [31:0] dummy_instr_seed_i;
	// Trace: design.sv:44145:3
	input wire fetch_valid_i;
	// Trace: design.sv:44146:3
	input wire id_in_ready_i;
	// Trace: design.sv:44147:3
	output wire insert_dummy_instr_o;
	// Trace: design.sv:44148:3
	output wire [31:0] dummy_instr_data_o;
	// Trace: design.sv:44151:3
	localparam [31:0] TIMEOUT_CNT_W = 5;
	// Trace: design.sv:44152:3
	localparam [31:0] OP_W = 5;
	// Trace: design.sv:44154:3
	// removed localparam type dummy_instr_e
	// Trace: design.sv:44161:3
	// removed localparam type lfsr_data_t
	// Trace: design.sv:44167:3
	localparam [31:0] LFSR_OUT_W = 17;
	// Trace: design.sv:44169:3
	wire [16:0] lfsr_data;
	// Trace: design.sv:44170:3
	wire [4:0] dummy_cnt_incr;
	wire [4:0] dummy_cnt_threshold;
	// Trace: design.sv:44171:3
	wire [4:0] dummy_cnt_d;
	reg [4:0] dummy_cnt_q;
	// Trace: design.sv:44172:3
	wire dummy_cnt_en;
	// Trace: design.sv:44173:3
	wire lfsr_en;
	// Trace: design.sv:44174:3
	wire [16:0] lfsr_state;
	// Trace: design.sv:44175:3
	wire insert_dummy_instr;
	// Trace: design.sv:44176:3
	reg [6:0] dummy_set;
	// Trace: design.sv:44177:3
	reg [2:0] dummy_opcode;
	// Trace: design.sv:44178:3
	wire [31:0] dummy_instr;
	// Trace: design.sv:44179:3
	reg [31:0] dummy_instr_seed_q;
	wire [31:0] dummy_instr_seed_d;
	// Trace: design.sv:44182:3
	assign lfsr_en = insert_dummy_instr & id_in_ready_i;
	// Trace: design.sv:44184:3
	assign dummy_instr_seed_d = dummy_instr_seed_q ^ dummy_instr_seed_i;
	// Trace: design.sv:44186:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:44187:5
		if (!rst_ni)
			// Trace: design.sv:44188:7
			dummy_instr_seed_q <= 1'sb0;
		else if (dummy_instr_seed_en_i)
			// Trace: design.sv:44190:7
			dummy_instr_seed_q <= dummy_instr_seed_d;
	// Trace: design.sv:44194:3
	prim_lfsr #(
		.LfsrDw(ibex_pkg_LfsrWidth),
		.StateOutDw(LFSR_OUT_W),
		.DefaultSeed(RndCnstLfsrSeed),
		.StatePermEn(1'b1),
		.StatePerm(RndCnstLfsrPerm)
	) lfsr_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.seed_en_i(dummy_instr_seed_en_i),
		.seed_i(dummy_instr_seed_d),
		.lfsr_en_i(lfsr_en),
		.entropy_i(1'sb0),
		.state_o(lfsr_state)
	);
	// Trace: design.sv:44211:3
	function automatic [16:0] sv2v_cast_92F3A;
		input reg [16:0] inp;
		sv2v_cast_92F3A = inp;
	endfunction
	assign lfsr_data = sv2v_cast_92F3A(lfsr_state);
	// Trace: design.sv:44215:3
	assign dummy_cnt_threshold = lfsr_data[4-:TIMEOUT_CNT_W] & {dummy_instr_mask_i, {2 {1'b1}}};
	// Trace: design.sv:44216:3
	assign dummy_cnt_incr = dummy_cnt_q + {{4 {1'b0}}, 1'b1};
	// Trace: design.sv:44218:3
	assign dummy_cnt_d = (insert_dummy_instr ? {5 {1'sb0}} : dummy_cnt_incr);
	// Trace: design.sv:44221:3
	assign dummy_cnt_en = (dummy_instr_en_i & id_in_ready_i) & (fetch_valid_i | insert_dummy_instr);
	// Trace: design.sv:44224:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:44225:5
		if (!rst_ni)
			// Trace: design.sv:44226:7
			dummy_cnt_q <= 1'sb0;
		else if (dummy_cnt_en)
			// Trace: design.sv:44228:7
			dummy_cnt_q <= dummy_cnt_d;
	// Trace: design.sv:44233:3
	assign insert_dummy_instr = dummy_instr_en_i & (dummy_cnt_q == dummy_cnt_threshold);
	// Trace: design.sv:44236:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:44237:5
		(* full_case, parallel_case *)
		case (lfsr_data[16-:2])
			2'b00: begin
				// Trace: design.sv:44239:9
				dummy_set = 7'b0000000;
				// Trace: design.sv:44240:9
				dummy_opcode = 3'b000;
			end
			2'b01: begin
				// Trace: design.sv:44243:9
				dummy_set = 7'b0000001;
				// Trace: design.sv:44244:9
				dummy_opcode = 3'b000;
			end
			2'b10: begin
				// Trace: design.sv:44247:9
				dummy_set = 7'b0000001;
				// Trace: design.sv:44248:9
				dummy_opcode = 3'b100;
			end
			2'b11: begin
				// Trace: design.sv:44251:9
				dummy_set = 7'b0000000;
				// Trace: design.sv:44252:9
				dummy_opcode = 3'b111;
			end
			default: begin
				// Trace: design.sv:44255:9
				dummy_set = 7'b0000000;
				// Trace: design.sv:44256:9
				dummy_opcode = 3'b000;
			end
		endcase
	end
	// Trace: design.sv:44262:3
	assign dummy_instr = {dummy_set, lfsr_data[14-:5], lfsr_data[9-:5], dummy_opcode, 12'h033};
	// Trace: design.sv:44265:3
	assign insert_dummy_instr_o = insert_dummy_instr;
	// Trace: design.sv:44266:3
	assign dummy_instr_data_o = dummy_instr;
	initial _sv2v_0 = 0;
endmodule
module ibex_core (
	clk_i,
	rst_ni,
	hart_id_i,
	boot_addr_i,
	instr_req_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_addr_o,
	instr_rdata_i,
	instr_err_i,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_we_o,
	data_be_o,
	data_addr_o,
	data_wdata_o,
	data_rdata_i,
	data_err_i,
	dummy_instr_id_o,
	rf_raddr_a_o,
	rf_raddr_b_o,
	rf_waddr_wb_o,
	rf_we_wb_o,
	rf_wdata_wb_ecc_o,
	rf_rdata_a_ecc_i,
	rf_rdata_b_ecc_i,
	ic_tag_req_o,
	ic_tag_write_o,
	ic_tag_addr_o,
	ic_tag_wdata_o,
	ic_tag_rdata_i,
	ic_data_req_o,
	ic_data_write_o,
	ic_data_addr_o,
	ic_data_wdata_o,
	ic_data_rdata_i,
	ic_scr_key_valid_i,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	irq_fast_i,
	irq_nm_i,
	irq_pending_o,
	debug_req_i,
	crash_dump_o,
	double_fault_seen_o,
	fetch_enable_i,
	alert_minor_o,
	alert_major_o,
	icache_inval_o,
	core_sleep_o
);
	// removed import ibex_pkg::*;
	// Trace: design.sv:44284:13
	parameter [0:0] PMPEnable = 1'b0;
	// Trace: design.sv:44285:13
	parameter [31:0] PMPGranularity = 0;
	// Trace: design.sv:44286:13
	parameter [31:0] PMPNumRegions = 4;
	// Trace: design.sv:44287:13
	parameter [31:0] MHPMCounterNum = 0;
	// Trace: design.sv:44288:13
	parameter [31:0] MHPMCounterWidth = 40;
	// Trace: design.sv:44289:13
	parameter [0:0] RV32E = 1'b0;
	// Trace: design.sv:44290:13
	// removed localparam type ibex_pkg_rv32m_e
	parameter integer RV32M = 32'sd2;
	// Trace: design.sv:44291:13
	// removed localparam type ibex_pkg_rv32b_e
	parameter integer RV32B = 32'sd0;
	// Trace: design.sv:44292:13
	parameter [0:0] BranchTargetALU = 1'b0;
	// Trace: design.sv:44293:13
	parameter [0:0] WritebackStage = 1'b0;
	// Trace: design.sv:44294:13
	parameter [0:0] ICache = 1'b0;
	// Trace: design.sv:44295:13
	parameter [0:0] ICacheECC = 1'b0;
	// Trace: design.sv:44296:13
	localparam [31:0] ibex_pkg_BUS_SIZE = 32;
	parameter [31:0] BusSizeECC = ibex_pkg_BUS_SIZE;
	// Trace: design.sv:44297:13
	localparam [31:0] ibex_pkg_ADDR_W = 32;
	localparam [31:0] ibex_pkg_IC_LINE_SIZE = 64;
	localparam [31:0] ibex_pkg_IC_LINE_BYTES = 8;
	localparam [31:0] ibex_pkg_IC_NUM_WAYS = 2;
	localparam [31:0] ibex_pkg_IC_SIZE_BYTES = 4096;
	localparam [31:0] ibex_pkg_IC_NUM_LINES = (ibex_pkg_IC_SIZE_BYTES / ibex_pkg_IC_NUM_WAYS) / ibex_pkg_IC_LINE_BYTES;
	localparam [31:0] ibex_pkg_IC_INDEX_W = $clog2(ibex_pkg_IC_NUM_LINES);
	localparam [31:0] ibex_pkg_IC_LINE_W = 3;
	localparam [31:0] ibex_pkg_IC_TAG_SIZE = ((ibex_pkg_ADDR_W - ibex_pkg_IC_INDEX_W) - ibex_pkg_IC_LINE_W) + 1;
	parameter [31:0] TagSizeECC = ibex_pkg_IC_TAG_SIZE;
	// Trace: design.sv:44298:13
	parameter [31:0] LineSizeECC = ibex_pkg_IC_LINE_SIZE;
	// Trace: design.sv:44299:13
	parameter [0:0] BranchPredictor = 1'b0;
	// Trace: design.sv:44300:13
	parameter [0:0] DbgTriggerEn = 1'b0;
	// Trace: design.sv:44301:13
	parameter [31:0] DbgHwBreakNum = 1;
	// Trace: design.sv:44302:13
	parameter [0:0] ResetAll = 1'b0;
	// Trace: design.sv:44303:13
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	// removed localparam type ibex_pkg_lfsr_seed_t
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	// Trace: design.sv:44304:13
	// removed localparam type ibex_pkg_lfsr_perm_t
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	// Trace: design.sv:44305:13
	parameter [0:0] SecureIbex = 1'b0;
	// Trace: design.sv:44306:13
	parameter [0:0] DummyInstructions = 1'b0;
	// Trace: design.sv:44307:13
	parameter [0:0] RegFileECC = 1'b0;
	// Trace: design.sv:44308:13
	parameter [31:0] RegFileDataWidth = 32;
	// Trace: design.sv:44309:13
	parameter [31:0] DmHaltAddr = 32'h1a110800;
	// Trace: design.sv:44310:13
	parameter [31:0] DmExceptionAddr = 32'h1a110808;
	// Trace: design.sv:44313:3
	input wire clk_i;
	// Trace: design.sv:44314:3
	input wire rst_ni;
	// Trace: design.sv:44316:3
	input wire [31:0] hart_id_i;
	// Trace: design.sv:44317:3
	input wire [31:0] boot_addr_i;
	// Trace: design.sv:44320:3
	output wire instr_req_o;
	// Trace: design.sv:44321:3
	input wire instr_gnt_i;
	// Trace: design.sv:44322:3
	input wire instr_rvalid_i;
	// Trace: design.sv:44323:3
	output wire [31:0] instr_addr_o;
	// Trace: design.sv:44324:3
	input wire [31:0] instr_rdata_i;
	// Trace: design.sv:44325:3
	input wire instr_err_i;
	// Trace: design.sv:44328:3
	output wire data_req_o;
	// Trace: design.sv:44329:3
	input wire data_gnt_i;
	// Trace: design.sv:44330:3
	input wire data_rvalid_i;
	// Trace: design.sv:44331:3
	output wire data_we_o;
	// Trace: design.sv:44332:3
	output wire [3:0] data_be_o;
	// Trace: design.sv:44333:3
	output wire [31:0] data_addr_o;
	// Trace: design.sv:44334:3
	output wire [31:0] data_wdata_o;
	// Trace: design.sv:44335:3
	input wire [31:0] data_rdata_i;
	// Trace: design.sv:44336:3
	input wire data_err_i;
	// Trace: design.sv:44339:3
	output wire dummy_instr_id_o;
	// Trace: design.sv:44340:3
	output wire [4:0] rf_raddr_a_o;
	// Trace: design.sv:44341:3
	output wire [4:0] rf_raddr_b_o;
	// Trace: design.sv:44342:3
	output wire [4:0] rf_waddr_wb_o;
	// Trace: design.sv:44343:3
	output wire rf_we_wb_o;
	// Trace: design.sv:44344:3
	output wire [RegFileDataWidth - 1:0] rf_wdata_wb_ecc_o;
	// Trace: design.sv:44345:3
	input wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc_i;
	// Trace: design.sv:44346:3
	input wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc_i;
	// Trace: design.sv:44349:3
	output wire [1:0] ic_tag_req_o;
	// Trace: design.sv:44350:3
	output wire ic_tag_write_o;
	// Trace: design.sv:44351:3
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr_o;
	// Trace: design.sv:44352:3
	output wire [TagSizeECC - 1:0] ic_tag_wdata_o;
	// Trace: design.sv:44353:3
	input wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata_i;
	// Trace: design.sv:44354:3
	output wire [1:0] ic_data_req_o;
	// Trace: design.sv:44355:3
	output wire ic_data_write_o;
	// Trace: design.sv:44356:3
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr_o;
	// Trace: design.sv:44357:3
	output wire [LineSizeECC - 1:0] ic_data_wdata_o;
	// Trace: design.sv:44358:3
	input wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata_i;
	// Trace: design.sv:44359:3
	input wire ic_scr_key_valid_i;
	// Trace: design.sv:44362:3
	input wire irq_software_i;
	// Trace: design.sv:44363:3
	input wire irq_timer_i;
	// Trace: design.sv:44364:3
	input wire irq_external_i;
	// Trace: design.sv:44365:3
	input wire [14:0] irq_fast_i;
	// Trace: design.sv:44366:3
	input wire irq_nm_i;
	// Trace: design.sv:44367:3
	output wire irq_pending_o;
	// Trace: design.sv:44370:3
	input wire debug_req_i;
	// Trace: design.sv:44371:3
	// removed localparam type ibex_pkg_crash_dump_t
	output wire [127:0] crash_dump_o;
	// Trace: design.sv:44374:3
	output wire double_fault_seen_o;
	// Trace: design.sv:44411:3
	input wire fetch_enable_i;
	// Trace: design.sv:44412:3
	output wire alert_minor_o;
	// Trace: design.sv:44413:3
	output wire alert_major_o;
	// Trace: design.sv:44414:3
	output wire icache_inval_o;
	// Trace: design.sv:44415:3
	output wire core_sleep_o;
	// Trace: design.sv:44418:3
	localparam [31:0] PMP_NUM_CHAN = 3;
	// Trace: design.sv:44420:3
	localparam [0:0] DataIndTiming = SecureIbex;
	// Trace: design.sv:44421:3
	localparam [0:0] PCIncrCheck = SecureIbex;
	// Trace: design.sv:44422:3
	localparam [0:0] ShadowCSR = 1'b0;
	// Trace: design.sv:44425:3
	wire dummy_instr_id;
	// Trace: design.sv:44426:3
	wire instr_valid_id;
	// Trace: design.sv:44427:3
	wire instr_new_id;
	// Trace: design.sv:44428:3
	wire [31:0] instr_rdata_id;
	// Trace: design.sv:44429:3
	wire [31:0] instr_rdata_alu_id;
	// Trace: design.sv:44431:3
	wire [15:0] instr_rdata_c_id;
	// Trace: design.sv:44432:3
	wire instr_is_compressed_id;
	// Trace: design.sv:44433:3
	wire instr_perf_count_id;
	// Trace: design.sv:44434:3
	wire instr_bp_taken_id;
	// Trace: design.sv:44435:3
	wire instr_fetch_err;
	// Trace: design.sv:44436:3
	wire instr_fetch_err_plus2;
	// Trace: design.sv:44437:3
	wire illegal_c_insn_id;
	// Trace: design.sv:44438:3
	wire [31:0] pc_if;
	// Trace: design.sv:44439:3
	wire [31:0] pc_id;
	// Trace: design.sv:44440:3
	wire [31:0] pc_wb;
	// Trace: design.sv:44441:3
	wire [67:0] imd_val_d_ex;
	// Trace: design.sv:44442:3
	wire [67:0] imd_val_q_ex;
	// Trace: design.sv:44443:3
	wire [1:0] imd_val_we_ex;
	// Trace: design.sv:44445:3
	wire data_ind_timing;
	// Trace: design.sv:44446:3
	wire dummy_instr_en;
	// Trace: design.sv:44447:3
	wire [2:0] dummy_instr_mask;
	// Trace: design.sv:44448:3
	wire dummy_instr_seed_en;
	// Trace: design.sv:44449:3
	wire [31:0] dummy_instr_seed;
	// Trace: design.sv:44450:3
	wire icache_enable;
	// Trace: design.sv:44451:3
	wire icache_inval;
	// Trace: design.sv:44452:3
	wire icache_ecc_error;
	// Trace: design.sv:44453:3
	wire pc_mismatch_alert;
	// Trace: design.sv:44454:3
	wire csr_shadow_err;
	// Trace: design.sv:44456:3
	wire instr_first_cycle_id;
	// Trace: design.sv:44457:3
	wire instr_valid_clear;
	// Trace: design.sv:44458:3
	wire pc_set;
	// Trace: design.sv:44459:3
	wire nt_branch_mispredict;
	// Trace: design.sv:44460:3
	wire [31:0] nt_branch_addr;
	// Trace: design.sv:44461:3
	// removed localparam type ibex_pkg_pc_sel_e
	wire [2:0] pc_mux_id;
	// Trace: design.sv:44462:3
	// removed localparam type ibex_pkg_exc_pc_sel_e
	wire [1:0] exc_pc_mux_id;
	// Trace: design.sv:44463:3
	// removed localparam type ibex_pkg_exc_cause_e
	wire [5:0] exc_cause;
	// Trace: design.sv:44465:3
	wire lsu_load_err;
	// Trace: design.sv:44466:3
	wire lsu_store_err;
	// Trace: design.sv:44469:3
	wire lsu_addr_incr_req;
	// Trace: design.sv:44470:3
	wire [31:0] lsu_addr_last;
	// Trace: design.sv:44473:3
	wire [31:0] branch_target_ex;
	// Trace: design.sv:44474:3
	wire branch_decision;
	// Trace: design.sv:44477:3
	wire ctrl_busy;
	// Trace: design.sv:44478:3
	wire if_busy;
	// Trace: design.sv:44479:3
	wire lsu_busy;
	// Trace: design.sv:44482:3
	wire [4:0] rf_raddr_a;
	// Trace: design.sv:44483:3
	wire [31:0] rf_rdata_a;
	// Trace: design.sv:44484:3
	wire [4:0] rf_raddr_b;
	// Trace: design.sv:44485:3
	wire [31:0] rf_rdata_b;
	// Trace: design.sv:44486:3
	wire rf_ren_a;
	// Trace: design.sv:44487:3
	wire rf_ren_b;
	// Trace: design.sv:44488:3
	wire [4:0] rf_waddr_wb;
	// Trace: design.sv:44489:3
	wire [31:0] rf_wdata_wb;
	// Trace: design.sv:44492:3
	wire [31:0] rf_wdata_fwd_wb;
	// Trace: design.sv:44493:3
	wire [31:0] rf_wdata_lsu;
	// Trace: design.sv:44494:3
	wire rf_we_wb;
	// Trace: design.sv:44495:3
	wire rf_we_lsu;
	// Trace: design.sv:44496:3
	wire rf_ecc_err_comb;
	// Trace: design.sv:44498:3
	wire [4:0] rf_waddr_id;
	// Trace: design.sv:44499:3
	wire [31:0] rf_wdata_id;
	// Trace: design.sv:44500:3
	wire rf_we_id;
	// Trace: design.sv:44501:3
	wire rf_rd_a_wb_match;
	// Trace: design.sv:44502:3
	wire rf_rd_b_wb_match;
	// Trace: design.sv:44505:3
	// removed localparam type ibex_pkg_alu_op_e
	wire [6:0] alu_operator_ex;
	// Trace: design.sv:44506:3
	wire [31:0] alu_operand_a_ex;
	// Trace: design.sv:44507:3
	wire [31:0] alu_operand_b_ex;
	// Trace: design.sv:44509:3
	wire [31:0] bt_a_operand;
	// Trace: design.sv:44510:3
	wire [31:0] bt_b_operand;
	// Trace: design.sv:44512:3
	wire [31:0] alu_adder_result_ex;
	// Trace: design.sv:44513:3
	wire [31:0] result_ex;
	// Trace: design.sv:44516:3
	wire mult_en_ex;
	// Trace: design.sv:44517:3
	wire div_en_ex;
	// Trace: design.sv:44518:3
	wire mult_sel_ex;
	// Trace: design.sv:44519:3
	wire div_sel_ex;
	// Trace: design.sv:44520:3
	// removed localparam type ibex_pkg_md_op_e
	wire [1:0] multdiv_operator_ex;
	// Trace: design.sv:44521:3
	wire [1:0] multdiv_signed_mode_ex;
	// Trace: design.sv:44522:3
	wire [31:0] multdiv_operand_a_ex;
	// Trace: design.sv:44523:3
	wire [31:0] multdiv_operand_b_ex;
	// Trace: design.sv:44524:3
	wire multdiv_ready_id;
	// Trace: design.sv:44527:3
	wire csr_access;
	// Trace: design.sv:44528:3
	// removed localparam type ibex_pkg_csr_op_e
	wire [1:0] csr_op;
	// Trace: design.sv:44529:3
	wire csr_op_en;
	// Trace: design.sv:44530:3
	// removed localparam type ibex_pkg_csr_num_e
	wire [11:0] csr_addr;
	// Trace: design.sv:44531:3
	wire [31:0] csr_rdata;
	// Trace: design.sv:44532:3
	wire [31:0] csr_wdata;
	// Trace: design.sv:44533:3
	wire illegal_csr_insn_id;
	// Trace: design.sv:44538:3
	wire lsu_we;
	// Trace: design.sv:44539:3
	wire [1:0] lsu_type;
	// Trace: design.sv:44540:3
	wire lsu_sign_ext;
	// Trace: design.sv:44541:3
	wire lsu_req;
	// Trace: design.sv:44542:3
	wire [31:0] lsu_wdata;
	// Trace: design.sv:44543:3
	wire lsu_req_done;
	// Trace: design.sv:44546:3
	wire id_in_ready;
	// Trace: design.sv:44547:3
	wire ex_valid;
	// Trace: design.sv:44549:3
	wire lsu_resp_valid;
	// Trace: design.sv:44550:3
	wire lsu_resp_err;
	// Trace: design.sv:44553:3
	wire instr_req_int;
	// Trace: design.sv:44554:3
	wire instr_req_gated;
	// Trace: design.sv:44557:3
	wire en_wb;
	// Trace: design.sv:44558:3
	// removed localparam type ibex_pkg_wb_instr_type_e
	wire [1:0] instr_type_wb;
	// Trace: design.sv:44559:3
	wire ready_wb;
	// Trace: design.sv:44560:3
	wire rf_write_wb;
	// Trace: design.sv:44561:3
	wire outstanding_load_wb;
	// Trace: design.sv:44562:3
	wire outstanding_store_wb;
	// Trace: design.sv:44565:3
	wire nmi_mode;
	// Trace: design.sv:44566:3
	// removed localparam type ibex_pkg_irqs_t
	wire [17:0] irqs;
	// Trace: design.sv:44567:3
	wire csr_mstatus_mie;
	// Trace: design.sv:44568:3
	wire [31:0] csr_mepc;
	wire [31:0] csr_depc;
	// Trace: design.sv:44571:3
	wire [(PMPNumRegions * 34) - 1:0] csr_pmp_addr;
	// Trace: design.sv:44572:3
	// removed localparam type ibex_pkg_pmp_cfg_mode_e
	// removed localparam type ibex_pkg_pmp_cfg_t
	wire [(PMPNumRegions * 6) - 1:0] csr_pmp_cfg;
	// Trace: design.sv:44573:3
	// removed localparam type ibex_pkg_pmp_mseccfg_t
	wire [2:0] csr_pmp_mseccfg;
	// Trace: design.sv:44574:3
	wire [0:2] pmp_req_err;
	// Trace: design.sv:44575:3
	wire data_req_out;
	// Trace: design.sv:44577:3
	wire csr_save_if;
	// Trace: design.sv:44578:3
	wire csr_save_id;
	// Trace: design.sv:44579:3
	wire csr_save_wb;
	// Trace: design.sv:44580:3
	wire csr_restore_mret_id;
	// Trace: design.sv:44581:3
	wire csr_restore_dret_id;
	// Trace: design.sv:44582:3
	wire csr_save_cause;
	// Trace: design.sv:44583:3
	wire csr_mtvec_init;
	// Trace: design.sv:44584:3
	wire [31:0] csr_mtvec;
	// Trace: design.sv:44585:3
	wire [31:0] csr_mtval;
	// Trace: design.sv:44586:3
	wire csr_mstatus_tw;
	// Trace: design.sv:44587:3
	// removed localparam type ibex_pkg_priv_lvl_e
	wire [1:0] priv_mode_id;
	// Trace: design.sv:44588:3
	wire [1:0] priv_mode_lsu;
	// Trace: design.sv:44591:3
	wire debug_mode;
	// Trace: design.sv:44592:3
	// removed localparam type ibex_pkg_dbg_cause_e
	wire [2:0] debug_cause;
	// Trace: design.sv:44593:3
	wire debug_csr_save;
	// Trace: design.sv:44594:3
	wire debug_single_step;
	// Trace: design.sv:44595:3
	wire debug_ebreakm;
	// Trace: design.sv:44596:3
	wire debug_ebreaku;
	// Trace: design.sv:44597:3
	wire trigger_match;
	// Trace: design.sv:44601:3
	wire instr_id_done;
	// Trace: design.sv:44602:3
	wire instr_done_wb;
	// Trace: design.sv:44604:3
	wire perf_instr_ret_wb;
	// Trace: design.sv:44605:3
	wire perf_instr_ret_compressed_wb;
	// Trace: design.sv:44606:3
	wire perf_instr_ret_wb_spec;
	// Trace: design.sv:44607:3
	wire perf_instr_ret_compressed_wb_spec;
	// Trace: design.sv:44608:3
	wire perf_iside_wait;
	// Trace: design.sv:44609:3
	wire perf_dside_wait;
	// Trace: design.sv:44610:3
	wire perf_mul_wait;
	// Trace: design.sv:44611:3
	wire perf_div_wait;
	// Trace: design.sv:44612:3
	wire perf_jump;
	// Trace: design.sv:44613:3
	wire perf_branch;
	// Trace: design.sv:44614:3
	wire perf_tbranch;
	// Trace: design.sv:44615:3
	wire perf_load;
	// Trace: design.sv:44616:3
	wire perf_store;
	// Trace: design.sv:44619:3
	wire illegal_insn_id;
	wire unused_illegal_insn_id;
	// Trace: design.sv:44630:3
	wire clk;
	// Trace: design.sv:44631:3
	wire fetch_enable;
	// Trace: design.sv:44632:3
	wire wake_from_sleep;
	// Trace: design.sv:44634:3
	cve2_sleep_unit sleep_unit_i(
		.clk_ungated_i(clk_i),
		.rst_n(rst_ni),
		.clk_gated_o(clk),
		.scan_cg_en_i(1'b0),
		.core_sleep_o(core_sleep_o),
		.fetch_enable_i(fetch_enable_i),
		.fetch_enable_o(fetch_enable),
		.if_busy_i(if_busy),
		.ctrl_busy_i(ctrl_busy),
		.lsu_busy_i(lsu_busy),
		.wake_from_sleep_i(wake_from_sleep)
	);
	// Trace: design.sv:44662:3
	localparam [31:0] ibex_pkg_PMP_I = 0;
	localparam [31:0] ibex_pkg_PMP_I2 = 1;
	ibex_if_stage #(
		.DmHaltAddr(DmHaltAddr),
		.DmExceptionAddr(DmExceptionAddr),
		.DummyInstructions(DummyInstructions),
		.ICache(ICache),
		.ICacheECC(ICacheECC),
		.BusSizeECC(BusSizeECC),
		.TagSizeECC(TagSizeECC),
		.LineSizeECC(LineSizeECC),
		.PCIncrCheck(PCIncrCheck),
		.ResetAll(ResetAll),
		.RndCnstLfsrSeed(RndCnstLfsrSeed),
		.RndCnstLfsrPerm(RndCnstLfsrPerm),
		.BranchPredictor(BranchPredictor)
	) if_stage_i(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.boot_addr_i(boot_addr_i),
		.req_i(instr_req_gated),
		.instr_req_o(instr_req_o),
		.instr_addr_o(instr_addr_o),
		.instr_gnt_i(instr_gnt_i),
		.instr_rvalid_i(instr_rvalid_i),
		.instr_rdata_i(instr_rdata_i),
		.instr_err_i(instr_err_i),
		.ic_tag_req_o(ic_tag_req_o),
		.ic_tag_write_o(ic_tag_write_o),
		.ic_tag_addr_o(ic_tag_addr_o),
		.ic_tag_wdata_o(ic_tag_wdata_o),
		.ic_tag_rdata_i(ic_tag_rdata_i),
		.ic_data_req_o(ic_data_req_o),
		.ic_data_write_o(ic_data_write_o),
		.ic_data_addr_o(ic_data_addr_o),
		.ic_data_wdata_o(ic_data_wdata_o),
		.ic_data_rdata_i(ic_data_rdata_i),
		.ic_scr_key_valid_i(ic_scr_key_valid_i),
		.instr_valid_id_o(instr_valid_id),
		.instr_new_id_o(instr_new_id),
		.instr_rdata_id_o(instr_rdata_id),
		.instr_rdata_alu_id_o(instr_rdata_alu_id),
		.instr_rdata_c_id_o(instr_rdata_c_id),
		.instr_is_compressed_id_o(instr_is_compressed_id),
		.instr_bp_taken_o(instr_bp_taken_id),
		.instr_fetch_err_o(instr_fetch_err),
		.instr_fetch_err_plus2_o(instr_fetch_err_plus2),
		.illegal_c_insn_id_o(illegal_c_insn_id),
		.dummy_instr_id_o(dummy_instr_id),
		.pc_if_o(pc_if),
		.pc_id_o(pc_id),
		.pmp_err_if_i(pmp_req_err[ibex_pkg_PMP_I]),
		.pmp_err_if_plus2_i(pmp_req_err[ibex_pkg_PMP_I2]),
		.instr_valid_clear_i(instr_valid_clear),
		.pc_set_i(pc_set),
		.pc_mux_i(pc_mux_id),
		.nt_branch_mispredict_i(nt_branch_mispredict),
		.exc_pc_mux_i(exc_pc_mux_id),
		.exc_cause(exc_cause),
		.dummy_instr_en_i(dummy_instr_en),
		.dummy_instr_mask_i(dummy_instr_mask),
		.dummy_instr_seed_en_i(dummy_instr_seed_en),
		.dummy_instr_seed_i(dummy_instr_seed),
		.icache_enable_i(icache_enable),
		.icache_inval_i(icache_inval),
		.icache_ecc_error_o(icache_ecc_error),
		.branch_target_ex_i(branch_target_ex),
		.nt_branch_addr_i(nt_branch_addr),
		.csr_mepc_i(csr_mepc),
		.csr_depc_i(csr_depc),
		.csr_mtvec_i(csr_mtvec),
		.csr_mtvec_init_o(csr_mtvec_init),
		.id_in_ready_i(id_in_ready),
		.pc_mismatch_alert_o(pc_mismatch_alert),
		.if_busy_o(if_busy)
	);
	// Trace: design.sv:44754:3
	assign perf_iside_wait = id_in_ready & ~instr_valid_id;
	// Trace: design.sv:44757:3
	assign instr_req_gated = instr_req_int & fetch_enable;
	// Trace: design.sv:44763:3
	ibex_id_stage #(
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU),
		.DataIndTiming(DataIndTiming),
		.WritebackStage(WritebackStage),
		.BranchPredictor(BranchPredictor)
	) id_stage_i(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.ctrl_busy_o(ctrl_busy),
		.illegal_insn_o(illegal_insn_id),
		.instr_valid_i(instr_valid_id),
		.instr_rdata_i(instr_rdata_id),
		.instr_rdata_alu_i(instr_rdata_alu_id),
		.instr_rdata_c_i(instr_rdata_c_id),
		.instr_is_compressed_i(instr_is_compressed_id),
		.instr_bp_taken_i(instr_bp_taken_id),
		.branch_decision_i(branch_decision),
		.instr_first_cycle_id_o(instr_first_cycle_id),
		.instr_valid_clear_o(instr_valid_clear),
		.id_in_ready_o(id_in_ready),
		.instr_req_o(instr_req_int),
		.pc_set_o(pc_set),
		.pc_mux_o(pc_mux_id),
		.nt_branch_mispredict_o(nt_branch_mispredict),
		.nt_branch_addr_o(nt_branch_addr),
		.exc_pc_mux_o(exc_pc_mux_id),
		.exc_cause_o(exc_cause),
		.icache_inval_o(icache_inval),
		.instr_fetch_err_i(instr_fetch_err),
		.instr_fetch_err_plus2_i(instr_fetch_err_plus2),
		.illegal_c_insn_i(illegal_c_insn_id),
		.pc_id_i(pc_id),
		.ex_valid_i(ex_valid),
		.lsu_resp_valid_i(lsu_resp_valid),
		.alu_operator_ex_o(alu_operator_ex),
		.alu_operand_a_ex_o(alu_operand_a_ex),
		.alu_operand_b_ex_o(alu_operand_b_ex),
		.imd_val_q_ex_o(imd_val_q_ex),
		.imd_val_d_ex_i(imd_val_d_ex),
		.imd_val_we_ex_i(imd_val_we_ex),
		.bt_a_operand_o(bt_a_operand),
		.bt_b_operand_o(bt_b_operand),
		.mult_en_ex_o(mult_en_ex),
		.div_en_ex_o(div_en_ex),
		.mult_sel_ex_o(mult_sel_ex),
		.div_sel_ex_o(div_sel_ex),
		.multdiv_operator_ex_o(multdiv_operator_ex),
		.multdiv_signed_mode_ex_o(multdiv_signed_mode_ex),
		.multdiv_operand_a_ex_o(multdiv_operand_a_ex),
		.multdiv_operand_b_ex_o(multdiv_operand_b_ex),
		.multdiv_ready_id_o(multdiv_ready_id),
		.csr_access_o(csr_access),
		.csr_op_o(csr_op),
		.csr_op_en_o(csr_op_en),
		.csr_save_if_o(csr_save_if),
		.csr_save_id_o(csr_save_id),
		.csr_save_wb_o(csr_save_wb),
		.csr_restore_mret_id_o(csr_restore_mret_id),
		.csr_restore_dret_id_o(csr_restore_dret_id),
		.csr_save_cause_o(csr_save_cause),
		.csr_mtval_o(csr_mtval),
		.priv_mode_i(priv_mode_id),
		.csr_mstatus_tw_i(csr_mstatus_tw),
		.illegal_csr_insn_i(illegal_csr_insn_id),
		.data_ind_timing_i(data_ind_timing),
		.lsu_req_o(lsu_req),
		.lsu_we_o(lsu_we),
		.lsu_type_o(lsu_type),
		.lsu_sign_ext_o(lsu_sign_ext),
		.lsu_wdata_o(lsu_wdata),
		.lsu_req_done_i(lsu_req_done),
		.lsu_addr_incr_req_i(lsu_addr_incr_req),
		.lsu_addr_last_i(lsu_addr_last),
		.lsu_load_err_i(lsu_load_err),
		.lsu_store_err_i(lsu_store_err),
		.csr_mstatus_mie_i(csr_mstatus_mie),
		.irq_pending_i(irq_pending_o),
		.irqs_i(irqs),
		.irq_nm_i(irq_nm_i),
		.nmi_mode_o(nmi_mode),
		.debug_mode_o(debug_mode),
		.debug_cause_o(debug_cause),
		.debug_csr_save_o(debug_csr_save),
		.debug_req_i(debug_req_i),
		.debug_single_step_i(debug_single_step),
		.debug_ebreakm_i(debug_ebreakm),
		.debug_ebreaku_i(debug_ebreaku),
		.trigger_match_i(trigger_match),
		.wake_from_sleep_o(wake_from_sleep),
		.result_ex_i(result_ex),
		.csr_rdata_i(csr_rdata),
		.rf_raddr_a_o(rf_raddr_a),
		.rf_rdata_a_i(rf_rdata_a),
		.rf_raddr_b_o(rf_raddr_b),
		.rf_rdata_b_i(rf_rdata_b),
		.rf_ren_a_o(rf_ren_a),
		.rf_ren_b_o(rf_ren_b),
		.rf_waddr_id_o(rf_waddr_id),
		.rf_wdata_id_o(rf_wdata_id),
		.rf_we_id_o(rf_we_id),
		.rf_rd_a_wb_match_o(rf_rd_a_wb_match),
		.rf_rd_b_wb_match_o(rf_rd_b_wb_match),
		.rf_waddr_wb_i(rf_waddr_wb),
		.rf_wdata_fwd_wb_i(rf_wdata_fwd_wb),
		.rf_write_wb_i(rf_write_wb),
		.en_wb_o(en_wb),
		.instr_type_wb_o(instr_type_wb),
		.instr_perf_count_id_o(instr_perf_count_id),
		.ready_wb_i(ready_wb),
		.outstanding_load_wb_i(outstanding_load_wb),
		.outstanding_store_wb_i(outstanding_store_wb),
		.perf_jump_o(perf_jump),
		.perf_branch_o(perf_branch),
		.perf_tbranch_o(perf_tbranch),
		.perf_dside_wait_o(perf_dside_wait),
		.perf_mul_wait_o(perf_mul_wait),
		.perf_div_wait_o(perf_div_wait),
		.instr_id_done_o(instr_id_done)
	);
	// Trace: design.sv:44922:3
	assign icache_inval_o = icache_inval;
	// Trace: design.sv:44924:3
	assign unused_illegal_insn_id = illegal_insn_id;
	// Trace: design.sv:44926:3
	ibex_ex_block #(
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU)
	) ex_block_i(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.alu_operator_i(alu_operator_ex),
		.alu_operand_a_i(alu_operand_a_ex),
		.alu_operand_b_i(alu_operand_b_ex),
		.alu_instr_first_cycle_i(instr_first_cycle_id),
		.bt_a_operand_i(bt_a_operand),
		.bt_b_operand_i(bt_b_operand),
		.multdiv_operator_i(multdiv_operator_ex),
		.mult_en_i(mult_en_ex),
		.div_en_i(div_en_ex),
		.mult_sel_i(mult_sel_ex),
		.div_sel_i(div_sel_ex),
		.multdiv_signed_mode_i(multdiv_signed_mode_ex),
		.multdiv_operand_a_i(multdiv_operand_a_ex),
		.multdiv_operand_b_i(multdiv_operand_b_ex),
		.multdiv_ready_id_i(multdiv_ready_id),
		.data_ind_timing_i(data_ind_timing),
		.imd_val_we_o(imd_val_we_ex),
		.imd_val_d_o(imd_val_d_ex),
		.imd_val_q_i(imd_val_q_ex),
		.alu_adder_result_ex_o(alu_adder_result_ex),
		.result_ex_o(result_ex),
		.branch_target_o(branch_target_ex),
		.branch_decision_o(branch_decision),
		.ex_valid_o(ex_valid)
	);
	// Trace: design.sv:44975:3
	localparam [31:0] ibex_pkg_PMP_D = 2;
	assign data_req_o = data_req_out & ~pmp_req_err[ibex_pkg_PMP_D];
	// Trace: design.sv:44976:3
	assign lsu_resp_err = lsu_load_err | lsu_store_err;
	// Trace: design.sv:44978:3
	ibex_load_store_unit load_store_unit_i(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.data_req_o(data_req_out),
		.data_gnt_i(data_gnt_i),
		.data_rvalid_i(data_rvalid_i),
		.data_err_i(data_err_i),
		.data_pmp_err_i(pmp_req_err[ibex_pkg_PMP_D]),
		.data_addr_o(data_addr_o),
		.data_we_o(data_we_o),
		.data_be_o(data_be_o),
		.data_wdata_o(data_wdata_o),
		.data_rdata_i(data_rdata_i),
		.lsu_we_i(lsu_we),
		.lsu_type_i(lsu_type),
		.lsu_wdata_i(lsu_wdata),
		.lsu_sign_ext_i(lsu_sign_ext),
		.lsu_rdata_o(rf_wdata_lsu),
		.lsu_rdata_valid_o(rf_we_lsu),
		.lsu_req_i(lsu_req),
		.lsu_req_done_o(lsu_req_done),
		.adder_result_ex_i(alu_adder_result_ex),
		.addr_incr_req_o(lsu_addr_incr_req),
		.addr_last_o(lsu_addr_last),
		.lsu_resp_valid_o(lsu_resp_valid),
		.load_err_o(lsu_load_err),
		.store_err_o(lsu_store_err),
		.busy_o(lsu_busy),
		.perf_load_o(perf_load),
		.perf_store_o(perf_store)
	);
	// Trace: design.sv:45024:3
	ibex_wb_stage #(
		.ResetAll(ResetAll),
		.WritebackStage(WritebackStage)
	) wb_stage_i(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.en_wb_i(en_wb),
		.instr_type_wb_i(instr_type_wb),
		.pc_id_i(pc_id),
		.instr_is_compressed_id_i(instr_is_compressed_id),
		.instr_perf_count_id_i(instr_perf_count_id),
		.ready_wb_o(ready_wb),
		.rf_write_wb_o(rf_write_wb),
		.outstanding_load_wb_o(outstanding_load_wb),
		.outstanding_store_wb_o(outstanding_store_wb),
		.pc_wb_o(pc_wb),
		.perf_instr_ret_wb_o(perf_instr_ret_wb),
		.perf_instr_ret_compressed_wb_o(perf_instr_ret_compressed_wb),
		.perf_instr_ret_wb_spec_o(perf_instr_ret_wb_spec),
		.perf_instr_ret_compressed_wb_spec_o(perf_instr_ret_compressed_wb_spec),
		.rf_waddr_id_i(rf_waddr_id),
		.rf_wdata_id_i(rf_wdata_id),
		.rf_we_id_i(rf_we_id),
		.rf_wdata_lsu_i(rf_wdata_lsu),
		.rf_we_lsu_i(rf_we_lsu),
		.rf_wdata_fwd_wb_o(rf_wdata_fwd_wb),
		.rf_waddr_wb_o(rf_waddr_wb),
		.rf_wdata_wb_o(rf_wdata_wb),
		.rf_we_wb_o(rf_we_wb),
		.lsu_resp_valid_i(lsu_resp_valid),
		.lsu_resp_err_i(lsu_resp_err),
		.instr_done_wb_o(instr_done_wb)
	);
	// Trace: design.sv:45069:3
	assign dummy_instr_id_o = dummy_instr_id;
	// Trace: design.sv:45070:3
	assign rf_raddr_a_o = rf_raddr_a;
	// Trace: design.sv:45071:3
	assign rf_waddr_wb_o = rf_waddr_wb;
	// Trace: design.sv:45072:3
	assign rf_we_wb_o = rf_we_wb;
	// Trace: design.sv:45073:3
	assign rf_raddr_b_o = rf_raddr_b;
	// Trace: design.sv:45075:3
	generate
		if (RegFileECC) begin : gen_regfile_ecc
			// Trace: design.sv:45078:5
			wire [1:0] rf_ecc_err_a;
			wire [1:0] rf_ecc_err_b;
			// Trace: design.sv:45079:5
			wire rf_ecc_err_a_id;
			wire rf_ecc_err_b_id;
			// Trace: design.sv:45082:5
			prim_secded_inv_39_32_enc regfile_ecc_enc(
				.data_i(rf_wdata_wb),
				.data_o(rf_wdata_wb_ecc_o)
			);
			// Trace: design.sv:45088:5
			prim_secded_inv_39_32_dec regfile_ecc_dec_a(
				.data_i(rf_rdata_a_ecc_i),
				.data_o(),
				.syndrome_o(),
				.err_o(rf_ecc_err_a)
			);
			// Trace: design.sv:45094:5
			prim_secded_inv_39_32_dec regfile_ecc_dec_b(
				.data_i(rf_rdata_b_ecc_i),
				.data_o(),
				.syndrome_o(),
				.err_o(rf_ecc_err_b)
			);
			// Trace: design.sv:45102:5
			assign rf_rdata_a = rf_rdata_a_ecc_i[31:0];
			// Trace: design.sv:45103:5
			assign rf_rdata_b = rf_rdata_b_ecc_i[31:0];
			// Trace: design.sv:45106:5
			assign rf_ecc_err_a_id = (|rf_ecc_err_a & rf_ren_a) & ~rf_rd_a_wb_match;
			// Trace: design.sv:45107:5
			assign rf_ecc_err_b_id = (|rf_ecc_err_b & rf_ren_b) & ~rf_rd_b_wb_match;
			// Trace: design.sv:45110:5
			assign rf_ecc_err_comb = instr_valid_id & (rf_ecc_err_a_id | rf_ecc_err_b_id);
		end
		else begin : gen_no_regfile_ecc
			// Trace: design.sv:45113:5
			wire unused_rf_ren_a;
			wire unused_rf_ren_b;
			// Trace: design.sv:45114:5
			wire unused_rf_rd_a_wb_match;
			wire unused_rf_rd_b_wb_match;
			// Trace: design.sv:45116:5
			assign unused_rf_ren_a = rf_ren_a;
			// Trace: design.sv:45117:5
			assign unused_rf_ren_b = rf_ren_b;
			// Trace: design.sv:45118:5
			assign unused_rf_rd_a_wb_match = rf_rd_a_wb_match;
			// Trace: design.sv:45119:5
			assign unused_rf_rd_b_wb_match = rf_rd_b_wb_match;
			// Trace: design.sv:45120:5
			assign rf_wdata_wb_ecc_o = rf_wdata_wb;
			// Trace: design.sv:45121:5
			assign rf_rdata_a = rf_rdata_a_ecc_i;
			// Trace: design.sv:45122:5
			assign rf_rdata_b = rf_rdata_b_ecc_i;
			// Trace: design.sv:45123:5
			assign rf_ecc_err_comb = 1'b0;
		end
	endgenerate
	// Trace: design.sv:45130:3
	assign crash_dump_o[127-:32] = pc_id;
	// Trace: design.sv:45131:3
	assign crash_dump_o[95-:32] = pc_if;
	// Trace: design.sv:45132:3
	assign crash_dump_o[63-:32] = lsu_addr_last;
	// Trace: design.sv:45133:3
	assign crash_dump_o[31-:32] = csr_mepc;
	// Trace: design.sv:45140:3
	assign alert_minor_o = icache_ecc_error;
	// Trace: design.sv:45143:3
	assign alert_major_o = (rf_ecc_err_comb | pc_mismatch_alert) | csr_shadow_err;
	// Trace: design.sv:45195:3
	assign csr_wdata = alu_operand_a_ex;
	// Trace: design.sv:45196:3
	function automatic [11:0] sv2v_cast_12;
		input reg [11:0] inp;
		sv2v_cast_12 = inp;
	endfunction
	assign csr_addr = sv2v_cast_12((csr_access ? alu_operand_b_ex[11:0] : 12'b000000000000));
	// Trace: design.sv:45198:3
	ibex_cs_registers #(
		.DbgTriggerEn(DbgTriggerEn),
		.DbgHwBreakNum(DbgHwBreakNum),
		.DataIndTiming(DataIndTiming),
		.DummyInstructions(DummyInstructions),
		.ShadowCSR(ShadowCSR),
		.ICache(ICache),
		.MHPMCounterNum(MHPMCounterNum),
		.MHPMCounterWidth(MHPMCounterWidth),
		.PMPEnable(PMPEnable),
		.PMPGranularity(PMPGranularity),
		.PMPNumRegions(PMPNumRegions),
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B)
	) cs_registers_i(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.hart_id_i(hart_id_i),
		.priv_mode_id_o(priv_mode_id),
		.priv_mode_lsu_o(priv_mode_lsu),
		.csr_mtvec_o(csr_mtvec),
		.csr_mtvec_init_i(csr_mtvec_init),
		.boot_addr_i(boot_addr_i),
		.csr_access_i(csr_access),
		.csr_addr_i(csr_addr),
		.csr_wdata_i(csr_wdata),
		.csr_op_i(csr_op),
		.csr_op_en_i(csr_op_en),
		.csr_rdata_o(csr_rdata),
		.irq_software_i(irq_software_i),
		.irq_timer_i(irq_timer_i),
		.irq_external_i(irq_external_i),
		.irq_fast_i(irq_fast_i),
		.nmi_mode_i(nmi_mode),
		.irq_pending_o(irq_pending_o),
		.irqs_o(irqs),
		.csr_mstatus_mie_o(csr_mstatus_mie),
		.csr_mstatus_tw_o(csr_mstatus_tw),
		.csr_mepc_o(csr_mepc),
		.csr_pmp_cfg_o(csr_pmp_cfg),
		.csr_pmp_addr_o(csr_pmp_addr),
		.csr_pmp_mseccfg_o(csr_pmp_mseccfg),
		.csr_depc_o(csr_depc),
		.debug_mode_i(debug_mode),
		.debug_cause_i(debug_cause),
		.debug_csr_save_i(debug_csr_save),
		.debug_single_step_o(debug_single_step),
		.debug_ebreakm_o(debug_ebreakm),
		.debug_ebreaku_o(debug_ebreaku),
		.trigger_match_o(trigger_match),
		.pc_if_i(pc_if),
		.pc_id_i(pc_id),
		.pc_wb_i(pc_wb),
		.data_ind_timing_o(data_ind_timing),
		.dummy_instr_en_o(dummy_instr_en),
		.dummy_instr_mask_o(dummy_instr_mask),
		.dummy_instr_seed_en_o(dummy_instr_seed_en),
		.dummy_instr_seed_o(dummy_instr_seed),
		.icache_enable_o(icache_enable),
		.csr_shadow_err_o(csr_shadow_err),
		.csr_save_if_i(csr_save_if),
		.csr_save_id_i(csr_save_id),
		.csr_save_wb_i(csr_save_wb),
		.csr_restore_mret_i(csr_restore_mret_id),
		.csr_restore_dret_i(csr_restore_dret_id),
		.csr_save_cause_i(csr_save_cause),
		.csr_mcause_i(exc_cause),
		.csr_mtval_i(csr_mtval),
		.illegal_csr_insn_o(illegal_csr_insn_id),
		.double_fault_seen_o(double_fault_seen_o),
		.instr_ret_i(perf_instr_ret_wb),
		.instr_ret_compressed_i(perf_instr_ret_compressed_wb),
		.instr_ret_spec_i(perf_instr_ret_wb_spec),
		.instr_ret_compressed_spec_i(perf_instr_ret_compressed_wb_spec),
		.iside_wait_i(perf_iside_wait),
		.jump_i(perf_jump),
		.branch_i(perf_branch),
		.branch_taken_i(perf_tbranch),
		.mem_load_i(perf_load),
		.mem_store_i(perf_store),
		.dside_wait_i(perf_dside_wait),
		.mul_wait_i(perf_mul_wait),
		.div_wait_i(perf_div_wait)
	);
	// Trace: design.sv:45311:3
	// removed localparam type ibex_pkg_pmp_req_e
	generate
		if (PMPEnable) begin : g_pmp
			// Trace: design.sv:45312:5
			wire [101:0] pmp_req_addr;
			// Trace: design.sv:45313:5
			wire [5:0] pmp_req_type;
			// Trace: design.sv:45314:5
			wire [5:0] pmp_priv_lvl;
			// Trace: design.sv:45316:5
			assign pmp_req_addr[68+:34] = {2'b00, pc_if};
			// Trace: design.sv:45317:5
			assign pmp_req_type[4+:2] = 2'b00;
			// Trace: design.sv:45318:5
			assign pmp_priv_lvl[4+:2] = priv_mode_id;
			// Trace: design.sv:45319:5
			assign pmp_req_addr[34+:34] = {2'b00, pc_if + 32'd2};
			// Trace: design.sv:45320:5
			assign pmp_req_type[2+:2] = 2'b00;
			// Trace: design.sv:45321:5
			assign pmp_priv_lvl[2+:2] = priv_mode_id;
			// Trace: design.sv:45322:5
			assign pmp_req_addr[0+:34] = {2'b00, data_addr_o[31:0]};
			// Trace: design.sv:45323:5
			assign pmp_req_type[0+:2] = (data_we_o ? 2'b01 : 2'b10);
			// Trace: design.sv:45324:5
			assign pmp_priv_lvl[0+:2] = priv_mode_lsu;
			// Trace: design.sv:45326:5
			ibex_pmp #(
				.PMPGranularity(PMPGranularity),
				.PMPNumChan(PMP_NUM_CHAN),
				.PMPNumRegions(PMPNumRegions)
			) pmp_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.csr_pmp_cfg_i(csr_pmp_cfg),
				.csr_pmp_addr_i(csr_pmp_addr),
				.csr_pmp_mseccfg_i(csr_pmp_mseccfg),
				.priv_mode_i(pmp_priv_lvl),
				.pmp_req_addr_i(pmp_req_addr),
				.pmp_req_type_i(pmp_req_type),
				.pmp_req_err_o(pmp_req_err)
			);
		end
		else begin : g_no_pmp
			// Trace: design.sv:45345:5
			wire [1:0] unused_priv_lvl_ls;
			// Trace: design.sv:45346:5
			wire [(PMPNumRegions * 34) - 1:0] unused_csr_pmp_addr;
			// Trace: design.sv:45347:5
			wire [(PMPNumRegions * 6) - 1:0] unused_csr_pmp_cfg;
			// Trace: design.sv:45348:5
			wire [2:0] unused_csr_pmp_mseccfg;
			// Trace: design.sv:45349:5
			assign unused_priv_lvl_ls = priv_mode_lsu;
			// Trace: design.sv:45350:5
			assign unused_csr_pmp_addr = csr_pmp_addr;
			// Trace: design.sv:45351:5
			assign unused_csr_pmp_cfg = csr_pmp_cfg;
			// Trace: design.sv:45352:5
			assign unused_csr_pmp_mseccfg = csr_pmp_mseccfg;
			// Trace: design.sv:45355:5
			assign pmp_req_err[ibex_pkg_PMP_I] = 1'b0;
			// Trace: design.sv:45356:5
			assign pmp_req_err[ibex_pkg_PMP_I2] = 1'b0;
			// Trace: design.sv:45357:5
			assign pmp_req_err[ibex_pkg_PMP_D] = 1'b0;
		end
	endgenerate
	// Trace: design.sv:45867:3
	wire unused_instr_new_id;
	wire unused_instr_id_done;
	wire unused_instr_done_wb;
	// Trace: design.sv:45868:3
	assign unused_instr_id_done = instr_id_done;
	// Trace: design.sv:45869:3
	assign unused_instr_new_id = instr_new_id;
	// Trace: design.sv:45870:3
	assign unused_instr_done_wb = instr_done_wb;
endmodule
module cve2_sleep_unit (
	clk_ungated_i,
	rst_n,
	clk_gated_o,
	scan_cg_en_i,
	core_sleep_o,
	fetch_enable_i,
	fetch_enable_o,
	if_busy_i,
	ctrl_busy_i,
	lsu_busy_i,
	wake_from_sleep_i
);
	// Trace: design.sv:45922:5
	input wire clk_ungated_i;
	// Trace: design.sv:45923:5
	input wire rst_n;
	// Trace: design.sv:45924:5
	output wire clk_gated_o;
	// Trace: design.sv:45925:5
	input wire scan_cg_en_i;
	// Trace: design.sv:45928:5
	output wire core_sleep_o;
	// Trace: design.sv:45931:5
	input wire fetch_enable_i;
	// Trace: design.sv:45932:5
	output wire fetch_enable_o;
	// Trace: design.sv:45935:5
	input wire if_busy_i;
	// Trace: design.sv:45936:5
	input wire ctrl_busy_i;
	// Trace: design.sv:45937:5
	input wire lsu_busy_i;
	// Trace: design.sv:45940:5
	input wire wake_from_sleep_i;
	// Trace: design.sv:45943:3
	reg fetch_enable_q;
	// Trace: design.sv:45944:3
	wire fetch_enable_d;
	// Trace: design.sv:45945:3
	reg core_busy_q;
	// Trace: design.sv:45946:3
	wire core_busy_d;
	// Trace: design.sv:45947:3
	wire clock_en;
	// Trace: design.sv:45954:3
	assign fetch_enable_d = (fetch_enable_i ? 1'b1 : fetch_enable_q);
	// Trace: design.sv:45958:3
	assign core_busy_d = (if_busy_i || ctrl_busy_i) || lsu_busy_i;
	// Trace: design.sv:45961:3
	assign clock_en = fetch_enable_q && (wake_from_sleep_i || core_busy_q);
	// Trace: design.sv:45965:3
	assign core_sleep_o = fetch_enable_q && !clock_en;
	// Trace: design.sv:45968:3
	always @(posedge clk_ungated_i or negedge rst_n)
		// Trace: design.sv:45969:5
		if (rst_n == 1'b0) begin
			// Trace: design.sv:45970:7
			core_busy_q <= 1'b0;
			// Trace: design.sv:45971:7
			fetch_enable_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:45973:7
			core_busy_q <= core_busy_d;
			// Trace: design.sv:45974:7
			fetch_enable_q <= fetch_enable_d;
		end
	// Trace: design.sv:45979:3
	assign fetch_enable_o = fetch_enable_q;
	// Trace: design.sv:45982:3
	cve2_clock_gate core_clock_gate_i(
		.clk_i(clk_ungated_i),
		.en_i(clock_en),
		.scan_cg_en_i(scan_cg_en_i),
		.clk_o(clk_gated_o)
	);
endmodule
module debug_rom (
	clk_i,
	req_i,
	addr_i,
	rdata_o
);
	reg _sv2v_0;
	// Trace: design.sv:46012:3
	input wire clk_i;
	// Trace: design.sv:46013:3
	input wire req_i;
	// Trace: design.sv:46014:3
	input wire [63:0] addr_i;
	// Trace: design.sv:46015:3
	output reg [63:0] rdata_o;
	// Trace: design.sv:46018:3
	localparam [31:0] RomSize = 19;
	// Trace: design.sv:46020:3
	wire [1215:0] mem;
	// Trace: design.sv:46021:3
	assign mem = 1216'h7b2000737b2024737b30257310852423f1402473a85ff06f7b2024737b30257310052223001000737b2024737b3025731005262300c5151300c5551300000517fd5ff06ffa041ce3002474134004440300a40433f140247302041c63001474134004440300a4043310852023f140247300c5151300c55513000005177b3510737b2410730ff0000f04c0006f07c0006f00c0006f;
	// Trace: design.sv:46043:3
	reg [4:0] addr_q;
	// Trace: design.sv:46045:3
	always @(posedge clk_i)
		// Trace: design.sv:46046:5
		if (req_i)
			// Trace: design.sv:46047:7
			addr_q <= addr_i[7:3];
	// Trace: design.sv:46053:3
	function automatic [4:0] sv2v_cast_C6D38;
		input reg [4:0] inp;
		sv2v_cast_C6D38 = inp;
	endfunction
	always @(*) begin : p_outmux
		if (_sv2v_0)
			;
		// Trace: design.sv:46054:5
		rdata_o = 1'sb0;
		// Trace: design.sv:46055:5
		if (addr_q < sv2v_cast_C6D38(RomSize))
			// Trace: design.sv:46056:9
			rdata_o = mem[addr_q * 64+:64];
	end
	initial _sv2v_0 = 0;
endmodule
module debug_rom_one_scratch (
	clk_i,
	req_i,
	addr_i,
	rdata_o
);
	reg _sv2v_0;
	// Trace: design.sv:46078:3
	input wire clk_i;
	// Trace: design.sv:46079:3
	input wire req_i;
	// Trace: design.sv:46080:3
	input wire [63:0] addr_i;
	// Trace: design.sv:46081:3
	output reg [63:0] rdata_o;
	// Trace: design.sv:46084:3
	localparam [31:0] RomSize = 13;
	// Trace: design.sv:46086:3
	wire [831:0] mem;
	// Trace: design.sv:46087:3
	assign mem = 832'h7b2000737b20247310802423f1402473ab1ff06f7b20247310002223001000737b20247310002623fddff06ffc0418e30024741340044403f140247302041263001474134004440310802023f14024737b2410730ff0000f0340006f0500006f00c0006f;
	// Trace: design.sv:46103:3
	reg [3:0] addr_q;
	// Trace: design.sv:46105:3
	always @(posedge clk_i)
		// Trace: design.sv:46106:5
		if (req_i)
			// Trace: design.sv:46107:7
			addr_q <= addr_i[6:3];
	// Trace: design.sv:46113:3
	function automatic [3:0] sv2v_cast_F42D2;
		input reg [3:0] inp;
		sv2v_cast_F42D2 = inp;
	endfunction
	always @(*) begin : p_outmux
		if (_sv2v_0)
			;
		// Trace: design.sv:46114:5
		rdata_o = 1'sb0;
		// Trace: design.sv:46115:5
		if (addr_q < sv2v_cast_F42D2(RomSize))
			// Trace: design.sv:46116:9
			rdata_o = mem[addr_q * 64+:64];
	end
	initial _sv2v_0 = 0;
endmodule
module dm_csrs (
	clk_i,
	rst_ni,
	testmode_i,
	dmi_rst_ni,
	dmi_req_valid_i,
	dmi_req_ready_o,
	dmi_req_i,
	dmi_resp_valid_o,
	dmi_resp_ready_i,
	dmi_resp_o,
	ndmreset_o,
	dmactive_o,
	hartinfo_i,
	halted_i,
	unavailable_i,
	resumeack_i,
	hartsel_o,
	haltreq_o,
	resumereq_o,
	clear_resumeack_o,
	cmd_valid_o,
	cmd_o,
	cmderror_valid_i,
	cmderror_i,
	cmdbusy_i,
	progbuf_o,
	data_o,
	data_i,
	data_valid_i,
	sbaddress_o,
	sbaddress_i,
	sbaddress_write_valid_o,
	sbreadonaddr_o,
	sbautoincrement_o,
	sbaccess_o,
	sbreadondata_o,
	sbdata_o,
	sbdata_read_valid_o,
	sbdata_write_valid_o,
	sbdata_i,
	sbdata_valid_i,
	sbbusy_i,
	sberror_valid_i,
	sberror_i
);
	reg _sv2v_0;
	// Trace: design.sv:46139:13
	parameter [31:0] NrHarts = 1;
	// Trace: design.sv:46140:13
	parameter [31:0] BusWidth = 32;
	// Trace: design.sv:46141:13
	parameter [NrHarts - 1:0] SelectableHarts = {NrHarts {1'b1}};
	// Trace: design.sv:46143:3
	input wire clk_i;
	// Trace: design.sv:46144:3
	input wire rst_ni;
	// Trace: design.sv:46145:3
	input wire testmode_i;
	// Trace: design.sv:46146:3
	input wire dmi_rst_ni;
	// Trace: design.sv:46148:3
	input wire dmi_req_valid_i;
	// Trace: design.sv:46149:3
	output wire dmi_req_ready_o;
	// Trace: design.sv:46150:3
	// removed localparam type dm_dtm_op_e
	// removed localparam type dm_dmi_req_t
	input wire [40:0] dmi_req_i;
	// Trace: design.sv:46152:3
	output wire dmi_resp_valid_o;
	// Trace: design.sv:46153:3
	input wire dmi_resp_ready_i;
	// Trace: design.sv:46154:3
	// removed localparam type dm_dmi_resp_t
	output wire [33:0] dmi_resp_o;
	// Trace: design.sv:46156:3
	output wire ndmreset_o;
	// Trace: design.sv:46157:3
	output wire dmactive_o;
	// Trace: design.sv:46160:3
	// removed localparam type dm_hartinfo_t
	input wire [(NrHarts * 32) - 1:0] hartinfo_i;
	// Trace: design.sv:46161:3
	input wire [NrHarts - 1:0] halted_i;
	// Trace: design.sv:46162:3
	input wire [NrHarts - 1:0] unavailable_i;
	// Trace: design.sv:46163:3
	input wire [NrHarts - 1:0] resumeack_i;
	// Trace: design.sv:46165:3
	output wire [19:0] hartsel_o;
	// Trace: design.sv:46166:3
	output reg [NrHarts - 1:0] haltreq_o;
	// Trace: design.sv:46167:3
	output reg [NrHarts - 1:0] resumereq_o;
	// Trace: design.sv:46168:3
	output reg clear_resumeack_o;
	// Trace: design.sv:46170:3
	output wire cmd_valid_o;
	// Trace: design.sv:46171:3
	// removed localparam type dm_cmd_e
	// removed localparam type dm_command_t
	output wire [31:0] cmd_o;
	// Trace: design.sv:46172:3
	input wire cmderror_valid_i;
	// Trace: design.sv:46173:3
	// removed localparam type dm_cmderr_e
	input wire [2:0] cmderror_i;
	// Trace: design.sv:46174:3
	input wire cmdbusy_i;
	// Trace: design.sv:46176:3
	localparam [4:0] dm_ProgBufSize = 5'h08;
	output wire [255:0] progbuf_o;
	// Trace: design.sv:46177:3
	localparam [3:0] dm_DataCount = 4'h2;
	output wire [63:0] data_o;
	// Trace: design.sv:46179:3
	input wire [63:0] data_i;
	// Trace: design.sv:46180:3
	input wire data_valid_i;
	// Trace: design.sv:46182:3
	output wire [BusWidth - 1:0] sbaddress_o;
	// Trace: design.sv:46183:3
	input wire [BusWidth - 1:0] sbaddress_i;
	// Trace: design.sv:46184:3
	output reg sbaddress_write_valid_o;
	// Trace: design.sv:46186:3
	output wire sbreadonaddr_o;
	// Trace: design.sv:46187:3
	output wire sbautoincrement_o;
	// Trace: design.sv:46188:3
	output wire [2:0] sbaccess_o;
	// Trace: design.sv:46190:3
	output wire sbreadondata_o;
	// Trace: design.sv:46191:3
	output wire [BusWidth - 1:0] sbdata_o;
	// Trace: design.sv:46192:3
	output reg sbdata_read_valid_o;
	// Trace: design.sv:46193:3
	output reg sbdata_write_valid_o;
	// Trace: design.sv:46195:3
	input wire [BusWidth - 1:0] sbdata_i;
	// Trace: design.sv:46196:3
	input wire sbdata_valid_i;
	// Trace: design.sv:46198:3
	input wire sbbusy_i;
	// Trace: design.sv:46199:3
	input wire sberror_valid_i;
	// Trace: design.sv:46200:3
	input wire [2:0] sberror_i;
	// Trace: design.sv:46203:3
	localparam [31:0] HartSelLen = (NrHarts == 1 ? 1 : $clog2(NrHarts));
	// Trace: design.sv:46204:3
	localparam [31:0] NrHartsAligned = 2 ** HartSelLen;
	// Trace: design.sv:46206:3
	wire [1:0] dtm_op;
	// Trace: design.sv:46207:3
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	assign dtm_op = sv2v_cast_2(dmi_req_i[33-:2]);
	// Trace: design.sv:46209:3
	wire resp_queue_full;
	// Trace: design.sv:46210:3
	wire resp_queue_empty;
	// Trace: design.sv:46211:3
	wire resp_queue_push;
	// Trace: design.sv:46212:3
	wire resp_queue_pop;
	// Trace: design.sv:46213:3
	reg [31:0] resp_queue_data;
	// Trace: design.sv:46215:3
	// removed localparam type dm_dm_csr_e
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	localparam [7:0] DataEnd = sv2v_cast_8((8'h04 + {4'h0, dm_DataCount}) - 8'h01);
	// Trace: design.sv:46216:3
	localparam [7:0] ProgBufEnd = sv2v_cast_8((8'h20 + {4'h0, dm_ProgBufSize}) - 8'h01);
	// Trace: design.sv:46218:3
	reg [31:0] haltsum0;
	reg [31:0] haltsum1;
	reg [31:0] haltsum2;
	reg [31:0] haltsum3;
	// Trace: design.sv:46219:3
	reg [((((NrHarts - 1) / 32) + 1) * 32) - 1:0] halted;
	// Trace: design.sv:46220:3
	reg [(((NrHarts - 1) / 32) >= 0 ? ((((NrHarts - 1) / 32) + 1) * 32) - 1 : ((1 - ((NrHarts - 1) / 32)) * 32) + ((((NrHarts - 1) / 32) * 32) - 1)):(((NrHarts - 1) / 32) >= 0 ? 0 : ((NrHarts - 1) / 32) * 32)] halted_reshaped0;
	// Trace: design.sv:46221:3
	reg [(((NrHarts - 1) / 1024) >= 0 ? ((((NrHarts - 1) / 1024) + 1) * 32) - 1 : ((1 - ((NrHarts - 1) / 1024)) * 32) + ((((NrHarts - 1) / 1024) * 32) - 1)):(((NrHarts - 1) / 1024) >= 0 ? 0 : ((NrHarts - 1) / 1024) * 32)] halted_reshaped1;
	// Trace: design.sv:46222:3
	reg [(((NrHarts - 1) / 32768) >= 0 ? ((((NrHarts - 1) / 32768) + 1) * 32) - 1 : ((1 - ((NrHarts - 1) / 32768)) * 32) + ((((NrHarts - 1) / 32768) * 32) - 1)):(((NrHarts - 1) / 32768) >= 0 ? 0 : ((NrHarts - 1) / 32768) * 32)] halted_reshaped2;
	// Trace: design.sv:46223:3
	reg [((((NrHarts - 1) / 1024) + 1) * 32) - 1:0] halted_flat1;
	// Trace: design.sv:46224:3
	reg [((((NrHarts - 1) / 32768) + 1) * 32) - 1:0] halted_flat2;
	// Trace: design.sv:46225:3
	reg [31:0] halted_flat3;
	// Trace: design.sv:46228:3
	reg [14:0] hartsel_idx0;
	// Trace: design.sv:46229:3
	function automatic [14:0] sv2v_cast_15;
		input reg [14:0] inp;
		sv2v_cast_15 = inp;
	endfunction
	always @(*) begin : p_haltsum0
		if (_sv2v_0)
			;
		// Trace: design.sv:46230:5
		halted = 1'sb0;
		// Trace: design.sv:46231:5
		haltsum0 = 1'sb0;
		// Trace: design.sv:46232:5
		hartsel_idx0 = hartsel_o[19:5];
		// Trace: design.sv:46233:5
		halted[NrHarts - 1:0] = halted_i;
		// Trace: design.sv:46234:5
		halted_reshaped0 = halted;
		// Trace: design.sv:46235:5
		if (hartsel_idx0 < sv2v_cast_15(((NrHarts - 1) / 32) + 1))
			// Trace: design.sv:46236:7
			haltsum0 = halted_reshaped0[(((NrHarts - 1) / 32) >= 0 ? hartsel_idx0 : ((NrHarts - 1) / 32) - hartsel_idx0) * 32+:32];
	end
	// Trace: design.sv:46241:3
	reg [9:0] hartsel_idx1;
	// Trace: design.sv:46242:3
	function automatic [9:0] sv2v_cast_10;
		input reg [9:0] inp;
		sv2v_cast_10 = inp;
	endfunction
	always @(*) begin : p_reduction1
		if (_sv2v_0)
			;
		// Trace: design.sv:46243:5
		halted_flat1 = 1'sb0;
		// Trace: design.sv:46244:5
		haltsum1 = 1'sb0;
		// Trace: design.sv:46245:5
		hartsel_idx1 = hartsel_o[19:10];
		// Trace: design.sv:46247:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:46247:10
			reg [31:0] k;
			// Trace: design.sv:46247:10
			for (k = 0; k < (((NrHarts - 1) / 32) + 1); k = k + 1)
				begin
					// Trace: design.sv:46248:7
					halted_flat1[k] = |halted_reshaped0[(((NrHarts - 1) / 32) >= 0 ? k : ((NrHarts - 1) / 32) - k) * 32+:32];
				end
		end
		// Trace: design.sv:46250:5
		halted_reshaped1 = halted_flat1;
		if (hartsel_idx1 < sv2v_cast_10(((NrHarts - 1) / 1024) + 1))
			// Trace: design.sv:46253:7
			haltsum1 = halted_reshaped1[(((NrHarts - 1) / 1024) >= 0 ? hartsel_idx1 : ((NrHarts - 1) / 1024) - hartsel_idx1) * 32+:32];
	end
	// Trace: design.sv:46258:3
	reg [4:0] hartsel_idx2;
	// Trace: design.sv:46259:3
	function automatic [4:0] sv2v_cast_5;
		input reg [4:0] inp;
		sv2v_cast_5 = inp;
	endfunction
	always @(*) begin : p_reduction2
		if (_sv2v_0)
			;
		// Trace: design.sv:46260:5
		halted_flat2 = 1'sb0;
		// Trace: design.sv:46261:5
		haltsum2 = 1'sb0;
		// Trace: design.sv:46262:5
		hartsel_idx2 = hartsel_o[19:15];
		// Trace: design.sv:46264:5
		begin : sv2v_autoblock_2
			// Trace: design.sv:46264:10
			reg [31:0] k;
			// Trace: design.sv:46264:10
			for (k = 0; k < (((NrHarts - 1) / 1024) + 1); k = k + 1)
				begin
					// Trace: design.sv:46265:7
					halted_flat2[k] = |halted_reshaped1[(((NrHarts - 1) / 1024) >= 0 ? k : ((NrHarts - 1) / 1024) - k) * 32+:32];
				end
		end
		// Trace: design.sv:46267:5
		halted_reshaped2 = halted_flat2;
		if (hartsel_idx2 < sv2v_cast_5(((NrHarts - 1) / 32768) + 1))
			// Trace: design.sv:46270:7
			haltsum2 = halted_reshaped2[(((NrHarts - 1) / 32768) >= 0 ? hartsel_idx2 : ((NrHarts - 1) / 32768) - hartsel_idx2) * 32+:32];
	end
	// Trace: design.sv:46275:3
	always @(*) begin : p_reduction3
		if (_sv2v_0)
			;
		// Trace: design.sv:46276:5
		halted_flat3 = 1'sb0;
		// Trace: design.sv:46277:5
		begin : sv2v_autoblock_3
			// Trace: design.sv:46277:10
			reg [31:0] k;
			// Trace: design.sv:46277:10
			for (k = 0; k < ((NrHarts / 32768) + 1); k = k + 1)
				begin
					// Trace: design.sv:46278:7
					halted_flat3[k] = |halted_reshaped2[(((NrHarts - 1) / 32768) >= 0 ? k : ((NrHarts - 1) / 32768) - k) * 32+:32];
				end
		end
		// Trace: design.sv:46280:5
		haltsum3 = halted_flat3;
	end
	// Trace: design.sv:46284:3
	// removed localparam type dm_dmstatus_t
	reg [31:0] dmstatus;
	// Trace: design.sv:46285:3
	// removed localparam type dm_dmcontrol_t
	reg [31:0] dmcontrol_d;
	reg [31:0] dmcontrol_q;
	// Trace: design.sv:46286:3
	// removed localparam type dm_abstractcs_t
	reg [31:0] abstractcs;
	// Trace: design.sv:46287:3
	reg [2:0] cmderr_d;
	reg [2:0] cmderr_q;
	// Trace: design.sv:46288:3
	reg [31:0] command_d;
	reg [31:0] command_q;
	// Trace: design.sv:46289:3
	reg cmd_valid_d;
	reg cmd_valid_q;
	// Trace: design.sv:46290:3
	// removed localparam type dm_abstractauto_t
	reg [31:0] abstractauto_d;
	reg [31:0] abstractauto_q;
	// Trace: design.sv:46291:3
	// removed localparam type dm_sbcs_t
	reg [31:0] sbcs_d;
	reg [31:0] sbcs_q;
	// Trace: design.sv:46292:3
	reg [63:0] sbaddr_d;
	reg [63:0] sbaddr_q;
	// Trace: design.sv:46293:3
	reg [63:0] sbdata_d;
	reg [63:0] sbdata_q;
	// Trace: design.sv:46295:3
	wire [NrHarts - 1:0] havereset_d;
	reg [NrHarts - 1:0] havereset_q;
	// Trace: design.sv:46297:3
	reg [255:0] progbuf_d;
	reg [255:0] progbuf_q;
	// Trace: design.sv:46298:3
	reg [63:0] data_d;
	reg [63:0] data_q;
	// Trace: design.sv:46300:3
	reg [HartSelLen - 1:0] selected_hart;
	// Trace: design.sv:46303:3
	localparam [1:0] dm_DTM_SUCCESS = 2'h0;
	assign dmi_resp_o[1-:2] = dm_DTM_SUCCESS;
	// Trace: design.sv:46304:3
	assign dmi_resp_valid_o = ~resp_queue_empty;
	// Trace: design.sv:46305:3
	assign dmi_req_ready_o = ~resp_queue_full;
	// Trace: design.sv:46306:3
	assign resp_queue_push = dmi_req_valid_i & dmi_req_ready_o;
	// Trace: design.sv:46308:3
	assign sbautoincrement_o = sbcs_q[16];
	// Trace: design.sv:46309:3
	assign sbreadonaddr_o = sbcs_q[20];
	// Trace: design.sv:46310:3
	assign sbreadondata_o = sbcs_q[15];
	// Trace: design.sv:46311:3
	assign sbaccess_o = sbcs_q[19-:3];
	// Trace: design.sv:46312:3
	assign sbdata_o = sbdata_q[BusWidth - 1:0];
	// Trace: design.sv:46313:3
	assign sbaddress_o = sbaddr_q[BusWidth - 1:0];
	// Trace: design.sv:46315:3
	assign hartsel_o = {dmcontrol_q[15-:10], dmcontrol_q[25-:10]};
	// Trace: design.sv:46318:3
	reg [NrHartsAligned - 1:0] havereset_d_aligned;
	wire [NrHartsAligned - 1:0] havereset_q_aligned;
	wire [NrHartsAligned - 1:0] resumeack_aligned;
	wire [NrHartsAligned - 1:0] unavailable_aligned;
	wire [NrHartsAligned - 1:0] halted_aligned;
	// Trace: design.sv:46321:3
	function automatic [NrHartsAligned - 1:0] sv2v_cast_DFF07;
		input reg [NrHartsAligned - 1:0] inp;
		sv2v_cast_DFF07 = inp;
	endfunction
	assign resumeack_aligned = sv2v_cast_DFF07(resumeack_i);
	// Trace: design.sv:46322:3
	assign unavailable_aligned = sv2v_cast_DFF07(unavailable_i);
	// Trace: design.sv:46323:3
	assign halted_aligned = sv2v_cast_DFF07(halted_i);
	// Trace: design.sv:46325:3
	function automatic [NrHarts - 1:0] sv2v_cast_178F2;
		input reg [NrHarts - 1:0] inp;
		sv2v_cast_178F2 = inp;
	endfunction
	assign havereset_d = sv2v_cast_178F2(havereset_d_aligned);
	// Trace: design.sv:46326:3
	assign havereset_q_aligned = sv2v_cast_DFF07(havereset_q);
	// Trace: design.sv:46328:3
	reg [(NrHartsAligned * 32) - 1:0] hartinfo_aligned;
	// Trace: design.sv:46329:3
	always @(*) begin : p_hartinfo_align
		if (_sv2v_0)
			;
		// Trace: design.sv:46330:5
		hartinfo_aligned = 1'sb0;
		// Trace: design.sv:46331:5
		hartinfo_aligned[32 * ((NrHarts - 1) - (NrHarts - 1))+:32 * NrHarts] = hartinfo_i;
	end
	// Trace: design.sv:46335:3
	wire [7:0] dm_csr_addr;
	// Trace: design.sv:46336:3
	reg [31:0] sbcs;
	// Trace: design.sv:46337:3
	reg [31:0] a_abstractcs;
	// Trace: design.sv:46338:3
	wire [3:0] autoexecdata_idx;
	// Trace: design.sv:46341:3
	assign dm_csr_addr = sv2v_cast_8({1'b0, dmi_req_i[40-:7]});
	// Trace: design.sv:46344:3
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	assign autoexecdata_idx = sv2v_cast_4({dm_csr_addr} - 8'h04);
	// Trace: design.sv:46346:3
	localparam [3:0] dm_DbgVersion013 = 4'h2;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	function automatic [$clog2(4'h2) - 1:0] sv2v_cast_68FD0;
		input reg [$clog2(4'h2) - 1:0] inp;
		sv2v_cast_68FD0 = inp;
	endfunction
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [11:0] sv2v_cast_12;
		input reg [11:0] inp;
		sv2v_cast_12 = inp;
	endfunction
	function automatic [15:0] sv2v_cast_16;
		input reg [15:0] inp;
		sv2v_cast_16 = inp;
	endfunction
	function automatic [6:0] sv2v_cast_1B50F;
		input reg [6:0] inp;
		sv2v_cast_1B50F = inp;
	endfunction
	always @(*) begin : csr_read_write
		if (_sv2v_0)
			;
		// Trace: design.sv:46351:5
		dmstatus = 1'sb0;
		// Trace: design.sv:46352:5
		dmstatus[3-:4] = dm_DbgVersion013;
		// Trace: design.sv:46354:5
		dmstatus[7] = 1'b1;
		// Trace: design.sv:46356:5
		dmstatus[5] = 1'b0;
		// Trace: design.sv:46358:5
		dmstatus[19] = havereset_q_aligned[selected_hart];
		// Trace: design.sv:46359:5
		dmstatus[18] = havereset_q_aligned[selected_hart];
		// Trace: design.sv:46361:5
		dmstatus[17] = resumeack_aligned[selected_hart];
		// Trace: design.sv:46362:5
		dmstatus[16] = resumeack_aligned[selected_hart];
		// Trace: design.sv:46364:5
		dmstatus[13] = unavailable_aligned[selected_hart];
		// Trace: design.sv:46365:5
		dmstatus[12] = unavailable_aligned[selected_hart];
		// Trace: design.sv:46369:5
		dmstatus[15] = sv2v_cast_32(hartsel_o) > (NrHarts - 32'sd1);
		// Trace: design.sv:46370:5
		dmstatus[14] = sv2v_cast_32(hartsel_o) > (NrHarts - 32'sd1);
		// Trace: design.sv:46374:5
		dmstatus[9] = halted_aligned[selected_hart] & ~unavailable_aligned[selected_hart];
		// Trace: design.sv:46375:5
		dmstatus[8] = halted_aligned[selected_hart] & ~unavailable_aligned[selected_hart];
		// Trace: design.sv:46377:5
		dmstatus[11] = ~halted_aligned[selected_hart] & ~unavailable_aligned[selected_hart];
		// Trace: design.sv:46378:5
		dmstatus[10] = ~halted_aligned[selected_hart] & ~unavailable_aligned[selected_hart];
		// Trace: design.sv:46381:5
		abstractcs = 1'sb0;
		// Trace: design.sv:46382:5
		abstractcs[3-:4] = dm_DataCount;
		// Trace: design.sv:46383:5
		abstractcs[28-:5] = dm_ProgBufSize;
		// Trace: design.sv:46384:5
		abstractcs[12] = cmdbusy_i;
		// Trace: design.sv:46385:5
		abstractcs[10-:3] = cmderr_q;
		// Trace: design.sv:46388:5
		abstractauto_d = abstractauto_q;
		// Trace: design.sv:46389:5
		abstractauto_d[15-:4] = 1'sb0;
		// Trace: design.sv:46392:5
		havereset_d_aligned = sv2v_cast_DFF07(havereset_q);
		// Trace: design.sv:46393:5
		dmcontrol_d = dmcontrol_q;
		// Trace: design.sv:46394:5
		cmderr_d = cmderr_q;
		// Trace: design.sv:46395:5
		command_d = command_q;
		// Trace: design.sv:46396:5
		progbuf_d = progbuf_q;
		// Trace: design.sv:46397:5
		data_d = data_q;
		// Trace: design.sv:46398:5
		sbcs_d = sbcs_q;
		// Trace: design.sv:46399:5
		sbaddr_d = sv2v_cast_64(sbaddress_i);
		// Trace: design.sv:46400:5
		sbdata_d = sbdata_q;
		// Trace: design.sv:46402:5
		resp_queue_data = 32'h00000000;
		// Trace: design.sv:46403:5
		cmd_valid_d = 1'b0;
		// Trace: design.sv:46404:5
		sbaddress_write_valid_o = 1'b0;
		// Trace: design.sv:46405:5
		sbdata_read_valid_o = 1'b0;
		// Trace: design.sv:46406:5
		sbdata_write_valid_o = 1'b0;
		// Trace: design.sv:46407:5
		clear_resumeack_o = 1'b0;
		// Trace: design.sv:46410:5
		sbcs = 1'sb0;
		// Trace: design.sv:46411:5
		a_abstractcs = 1'sb0;
		// Trace: design.sv:46414:5
		if ((dmi_req_ready_o && dmi_req_valid_i) && (dtm_op == 2'h1)) begin
			begin
				// Trace: design.sv:46415:7
				(* full_case, parallel_case *)
				if ((8'h04 <= dm_csr_addr) && (DataEnd >= dm_csr_addr)) begin
					// Trace: design.sv:46417:11
					resp_queue_data = data_q[sv2v_cast_68FD0(autoexecdata_idx) * 32+:32];
					// Trace: design.sv:46418:11
					if (!cmdbusy_i)
						// Trace: design.sv:46420:13
						cmd_valid_d = abstractauto_q[0 + autoexecdata_idx];
					else if (cmderr_q == 3'd0)
						// Trace: design.sv:46423:13
						cmderr_d = 3'd1;
				end
				else if (dm_csr_addr == 8'h10)
					// Trace: design.sv:46426:27
					resp_queue_data = dmcontrol_q;
				else if (dm_csr_addr == 8'h11)
					// Trace: design.sv:46427:27
					resp_queue_data = dmstatus;
				else if (dm_csr_addr == 8'h12)
					// Trace: design.sv:46428:27
					resp_queue_data = hartinfo_aligned[selected_hart * 32+:32];
				else if (dm_csr_addr == 8'h16)
					// Trace: design.sv:46429:27
					resp_queue_data = abstractcs;
				else if (dm_csr_addr == 8'h18)
					// Trace: design.sv:46430:27
					resp_queue_data = abstractauto_q;
				else if (dm_csr_addr == 8'h17)
					// Trace: design.sv:46432:25
					resp_queue_data = 1'sb0;
				else if ((8'h20 <= dm_csr_addr) && (ProgBufEnd >= dm_csr_addr)) begin
					// Trace: design.sv:46434:11
					resp_queue_data = progbuf_q[dmi_req_i[$clog2(5'h08) + 33:34] * 32+:32];
					// Trace: design.sv:46435:11
					if (!cmdbusy_i)
						// Trace: design.sv:46438:13
						cmd_valid_d = abstractauto_q[0 + {1'b1, dmi_req_i[37:34]}];
					else if (cmderr_q == 3'd0)
						// Trace: design.sv:46442:13
						cmderr_d = 3'd1;
				end
				else if (dm_csr_addr == 8'h40)
					// Trace: design.sv:46445:23
					resp_queue_data = haltsum0;
				else if (dm_csr_addr == 8'h13)
					// Trace: design.sv:46446:23
					resp_queue_data = haltsum1;
				else if (dm_csr_addr == 8'h34)
					// Trace: design.sv:46447:23
					resp_queue_data = haltsum2;
				else if (dm_csr_addr == 8'h35)
					// Trace: design.sv:46448:23
					resp_queue_data = haltsum3;
				else if (dm_csr_addr == 8'h38)
					// Trace: design.sv:46450:11
					resp_queue_data = sbcs_q;
				else if (dm_csr_addr == 8'h39)
					// Trace: design.sv:46453:11
					resp_queue_data = sbaddr_q[31:0];
				else if (dm_csr_addr == 8'h3a)
					// Trace: design.sv:46456:11
					resp_queue_data = sbaddr_q[63:32];
				else if (dm_csr_addr == 8'h3c) begin
					begin
						// Trace: design.sv:46460:11
						if (sbbusy_i || sbcs_q[22])
							// Trace: design.sv:46461:13
							sbcs_d[22] = 1'b1;
						else begin
							// Trace: design.sv:46463:13
							sbdata_read_valid_o = sbcs_q[14-:3] == {3 {1'sb0}};
							// Trace: design.sv:46464:13
							resp_queue_data = sbdata_q[31:0];
						end
					end
				end
				else if (dm_csr_addr == 8'h3d) begin
					begin
						// Trace: design.sv:46469:11
						if (sbbusy_i || sbcs_q[22])
							// Trace: design.sv:46470:13
							sbcs_d[22] = 1'b1;
						else
							// Trace: design.sv:46472:13
							resp_queue_data = sbdata_q[63:32];
					end
				end
			end
		end
		if ((dmi_req_ready_o && dmi_req_valid_i) && (dtm_op == 2'h2)) begin
			begin
				// Trace: design.sv:46481:7
				(* full_case, parallel_case *)
				if ((8'h04 <= dm_csr_addr) && (DataEnd >= dm_csr_addr)) begin
					// Trace: design.sv:46483:11
					// Trace: design.sv:46485:13
					if (!cmdbusy_i) begin
						// Trace: design.sv:46486:15
						data_d[dmi_req_i[$clog2(4'h2) + 33:34] * 32+:32] = dmi_req_i[31-:32];
						// Trace: design.sv:46488:15
						cmd_valid_d = abstractauto_q[0 + autoexecdata_idx];
					end
					else if (cmderr_q == 3'd0)
						// Trace: design.sv:46491:15
						cmderr_d = 3'd1;
				end
				else if (dm_csr_addr == 8'h10) begin
					// Trace: design.sv:46496:11
					dmcontrol_d = dmi_req_i[31-:32];
					// Trace: design.sv:46498:11
					if (dmcontrol_d[28])
						// Trace: design.sv:46499:13
						havereset_d_aligned[selected_hart] = 1'b0;
				end
				else if (dm_csr_addr == 8'h11)
					;
				else if (dm_csr_addr == 8'h12)
					;
				else if (dm_csr_addr == 8'h16) begin
					// Trace: design.sv:46510:11
					a_abstractcs = sv2v_cast_32(dmi_req_i[31-:32]);
					// Trace: design.sv:46512:11
					if (!cmdbusy_i)
						// Trace: design.sv:46513:13
						cmderr_d = sv2v_cast_3(~a_abstractcs[10-:3] & cmderr_q);
					else if (cmderr_q == 3'd0)
						// Trace: design.sv:46515:13
						cmderr_d = 3'd1;
				end
				else if (dm_csr_addr == 8'h17) begin
					begin
						// Trace: design.sv:46520:11
						if (!cmdbusy_i) begin
							// Trace: design.sv:46521:13
							cmd_valid_d = 1'b1;
							// Trace: design.sv:46522:13
							command_d = sv2v_cast_32(dmi_req_i[31-:32]);
						end
						else if (cmderr_q == 3'd0)
							// Trace: design.sv:46526:13
							cmderr_d = 3'd1;
					end
				end
				else if (dm_csr_addr == 8'h18) begin
					begin
						// Trace: design.sv:46531:11
						if (!cmdbusy_i) begin
							// Trace: design.sv:46532:13
							abstractauto_d = 32'h00000000;
							// Trace: design.sv:46533:13
							abstractauto_d[11-:12] = sv2v_cast_12(dmi_req_i[1:0]);
							// Trace: design.sv:46534:13
							abstractauto_d[31-:16] = sv2v_cast_16(dmi_req_i[23:16]);
						end
						else if (cmderr_q == 3'd0)
							// Trace: design.sv:46536:13
							cmderr_d = 3'd1;
					end
				end
				else if ((8'h20 <= dm_csr_addr) && (ProgBufEnd >= dm_csr_addr)) begin
					begin
						// Trace: design.sv:46541:11
						if (!cmdbusy_i) begin
							// Trace: design.sv:46542:13
							progbuf_d[dmi_req_i[$clog2(5'h08) + 33:34] * 32+:32] = dmi_req_i[31-:32];
							// Trace: design.sv:46547:13
							cmd_valid_d = abstractauto_q[0 + {1'b1, dmi_req_i[37:34]}];
						end
						else if (cmderr_q == 3'd0)
							// Trace: design.sv:46550:13
							cmderr_d = 3'd1;
					end
				end
				else if (dm_csr_addr == 8'h38) begin
					begin
						// Trace: design.sv:46555:11
						if (sbbusy_i)
							// Trace: design.sv:46556:13
							sbcs_d[22] = 1'b1;
						else begin
							// Trace: design.sv:46558:13
							sbcs = sv2v_cast_32(dmi_req_i[31-:32]);
							// Trace: design.sv:46559:13
							sbcs_d = sbcs;
							// Trace: design.sv:46561:13
							sbcs_d[22] = sbcs_q[22] & ~sbcs[22];
							// Trace: design.sv:46562:13
							sbcs_d[14-:3] = sbcs_q[14-:3] & {3 {~(sbcs[14-:3] == 3'd1)}};
						end
					end
				end
				else if (dm_csr_addr == 8'h39) begin
					begin
						// Trace: design.sv:46567:11
						if (sbbusy_i || sbcs_q[22])
							// Trace: design.sv:46568:13
							sbcs_d[22] = 1'b1;
						else begin
							// Trace: design.sv:46570:13
							sbaddr_d[31:0] = dmi_req_i[31-:32];
							// Trace: design.sv:46571:13
							sbaddress_write_valid_o = sbcs_q[14-:3] == {3 {1'sb0}};
						end
					end
				end
				else if (dm_csr_addr == 8'h3a) begin
					begin
						// Trace: design.sv:46576:11
						if (sbbusy_i || sbcs_q[22])
							// Trace: design.sv:46577:13
							sbcs_d[22] = 1'b1;
						else
							// Trace: design.sv:46579:13
							sbaddr_d[63:32] = dmi_req_i[31-:32];
					end
				end
				else if (dm_csr_addr == 8'h3c) begin
					begin
						// Trace: design.sv:46584:11
						if (sbbusy_i || sbcs_q[22])
							// Trace: design.sv:46585:12
							sbcs_d[22] = 1'b1;
						else begin
							// Trace: design.sv:46587:13
							sbdata_d[31:0] = dmi_req_i[31-:32];
							// Trace: design.sv:46588:13
							sbdata_write_valid_o = sbcs_q[14-:3] == {3 {1'sb0}};
						end
					end
				end
				else if (dm_csr_addr == 8'h3d) begin
					begin
						// Trace: design.sv:46593:11
						if (sbbusy_i || sbcs_q[22])
							// Trace: design.sv:46594:12
							sbcs_d[22] = 1'b1;
						else
							// Trace: design.sv:46596:13
							sbdata_d[63:32] = dmi_req_i[31-:32];
					end
				end
			end
		end
		if (cmderror_valid_i)
			// Trace: design.sv:46604:7
			cmderr_d = cmderror_i;
		if (data_valid_i)
			// Trace: design.sv:46609:7
			data_d = data_i;
		if (ndmreset_o)
			// Trace: design.sv:46614:7
			havereset_d_aligned[NrHarts - 1:0] = 1'sb1;
		if (sberror_valid_i)
			// Trace: design.sv:46621:7
			sbcs_d[14-:3] = sberror_i;
		if (sbdata_valid_i)
			// Trace: design.sv:46625:7
			sbdata_d = sv2v_cast_64(sbdata_i);
		// Trace: design.sv:46630:5
		dmcontrol_d[26] = 1'b0;
		// Trace: design.sv:46632:5
		dmcontrol_d[29] = 1'b0;
		// Trace: design.sv:46633:5
		dmcontrol_d[3] = 1'b0;
		// Trace: design.sv:46634:5
		dmcontrol_d[2] = 1'b0;
		// Trace: design.sv:46635:5
		dmcontrol_d[27] = 1'sb0;
		// Trace: design.sv:46636:5
		dmcontrol_d[5-:2] = 1'sb0;
		// Trace: design.sv:46638:5
		dmcontrol_d[28] = 1'b0;
		if (!dmcontrol_q[30] && dmcontrol_d[30])
			// Trace: design.sv:46640:7
			clear_resumeack_o = 1'b1;
		if (dmcontrol_q[30] && resumeack_i)
			// Trace: design.sv:46643:7
			dmcontrol_d[30] = 1'b0;
		// Trace: design.sv:46646:5
		sbcs_d[31-:3] = 3'd1;
		// Trace: design.sv:46647:5
		sbcs_d[21] = sbbusy_i;
		// Trace: design.sv:46648:5
		sbcs_d[11-:7] = sv2v_cast_1B50F(BusWidth);
		// Trace: design.sv:46649:5
		sbcs_d[4] = BusWidth >= 32'd128;
		// Trace: design.sv:46650:5
		sbcs_d[3] = BusWidth >= 32'd64;
		// Trace: design.sv:46651:5
		sbcs_d[2] = BusWidth >= 32'd32;
		// Trace: design.sv:46652:5
		sbcs_d[1] = BusWidth >= 32'd16;
		// Trace: design.sv:46653:5
		sbcs_d[0] = BusWidth >= 32'd8;
	end
	// Trace: design.sv:46657:3
	function automatic [HartSelLen - 1:0] sv2v_cast_FFD0D;
		input reg [HartSelLen - 1:0] inp;
		sv2v_cast_FFD0D = inp;
	endfunction
	always @(*) begin : p_outmux
		if (_sv2v_0)
			;
		// Trace: design.sv:46658:5
		selected_hart = hartsel_o[HartSelLen - 1:0];
		// Trace: design.sv:46660:5
		haltreq_o = 1'sb0;
		// Trace: design.sv:46661:5
		resumereq_o = 1'sb0;
		// Trace: design.sv:46662:5
		if (selected_hart <= sv2v_cast_FFD0D(NrHarts - 1)) begin
			// Trace: design.sv:46663:7
			haltreq_o[selected_hart] = dmcontrol_q[31];
			// Trace: design.sv:46664:7
			resumereq_o[selected_hart] = dmcontrol_q[30];
		end
	end
	// Trace: design.sv:46668:3
	assign dmactive_o = dmcontrol_q[0];
	// Trace: design.sv:46669:3
	assign cmd_o = command_q;
	// Trace: design.sv:46670:3
	assign cmd_valid_o = cmd_valid_q;
	// Trace: design.sv:46671:3
	assign progbuf_o = progbuf_q;
	// Trace: design.sv:46672:3
	assign data_o = data_q;
	// Trace: design.sv:46674:3
	assign resp_queue_pop = dmi_resp_ready_i & ~resp_queue_empty;
	// Trace: design.sv:46676:3
	assign ndmreset_o = dmcontrol_q[1];
	// Trace: design.sv:46679:3
	fifo_v2_264A2 #(.DEPTH(2)) i_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(~dmi_rst_ni),
		.testmode_i(testmode_i),
		.full_o(resp_queue_full),
		.empty_o(resp_queue_empty),
		.alm_full_o(),
		.alm_empty_o(),
		.data_i(resp_queue_data),
		.push_i(resp_queue_push),
		.data_o(dmi_resp_o[33-:32]),
		.pop_i(resp_queue_pop)
	);
	// Trace: design.sv:46698:3
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:46700:5
		if (!rst_ni) begin
			// Trace: design.sv:46701:7
			dmcontrol_q <= 1'sb0;
			// Trace: design.sv:46703:7
			cmderr_q <= 3'd0;
			// Trace: design.sv:46704:7
			command_q <= 1'sb0;
			// Trace: design.sv:46705:7
			cmd_valid_q <= 1'sb0;
			// Trace: design.sv:46706:7
			abstractauto_q <= 1'sb0;
			// Trace: design.sv:46707:7
			progbuf_q <= 1'sb0;
			// Trace: design.sv:46708:7
			data_q <= 1'sb0;
			// Trace: design.sv:46709:7
			sbcs_q <= 32'h00040000;
			// Trace: design.sv:46710:7
			sbaddr_q <= 1'sb0;
			// Trace: design.sv:46711:7
			sbdata_q <= 1'sb0;
			// Trace: design.sv:46712:7
			havereset_q <= 1'sb1;
		end
		else begin
			// Trace: design.sv:46714:7
			havereset_q <= SelectableHarts & havereset_d;
			// Trace: design.sv:46716:7
			if (!dmcontrol_q[0]) begin
				// Trace: design.sv:46717:9
				dmcontrol_q[31] <= 1'sb0;
				// Trace: design.sv:46718:9
				dmcontrol_q[30] <= 1'sb0;
				// Trace: design.sv:46719:9
				dmcontrol_q[29] <= 1'sb0;
				// Trace: design.sv:46720:9
				dmcontrol_q[28] <= 1'sb0;
				// Trace: design.sv:46721:9
				dmcontrol_q[27] <= 1'sb0;
				// Trace: design.sv:46722:9
				dmcontrol_q[26] <= 1'sb0;
				// Trace: design.sv:46723:9
				dmcontrol_q[25-:10] <= 1'sb0;
				// Trace: design.sv:46724:9
				dmcontrol_q[15-:10] <= 1'sb0;
				// Trace: design.sv:46725:9
				dmcontrol_q[5-:2] <= 1'sb0;
				// Trace: design.sv:46726:9
				dmcontrol_q[3] <= 1'sb0;
				// Trace: design.sv:46727:9
				dmcontrol_q[2] <= 1'sb0;
				// Trace: design.sv:46728:9
				dmcontrol_q[1] <= 1'sb0;
				// Trace: design.sv:46730:9
				dmcontrol_q[0] <= dmcontrol_d[0];
				// Trace: design.sv:46731:9
				cmderr_q <= 3'd0;
				// Trace: design.sv:46732:9
				command_q <= 1'sb0;
				// Trace: design.sv:46733:9
				cmd_valid_q <= 1'sb0;
				// Trace: design.sv:46734:9
				abstractauto_q <= 1'sb0;
				// Trace: design.sv:46735:9
				progbuf_q <= 1'sb0;
				// Trace: design.sv:46736:9
				data_q <= 1'sb0;
				// Trace: design.sv:46737:9
				sbcs_q <= 32'h00040000;
				// Trace: design.sv:46738:9
				sbaddr_q <= 1'sb0;
				// Trace: design.sv:46739:9
				sbdata_q <= 1'sb0;
			end
			else begin
				// Trace: design.sv:46741:9
				dmcontrol_q <= dmcontrol_d;
				// Trace: design.sv:46742:9
				cmderr_q <= cmderr_d;
				// Trace: design.sv:46743:9
				command_q <= command_d;
				// Trace: design.sv:46744:9
				cmd_valid_q <= cmd_valid_d;
				// Trace: design.sv:46745:9
				abstractauto_q <= abstractauto_d;
				// Trace: design.sv:46746:9
				progbuf_q <= progbuf_d;
				// Trace: design.sv:46747:9
				data_q <= data_d;
				// Trace: design.sv:46748:9
				sbcs_q <= sbcs_d;
				// Trace: design.sv:46749:9
				sbaddr_q <= sbaddr_d;
				// Trace: design.sv:46750:9
				sbdata_q <= sbdata_d;
			end
		end
	end
	initial _sv2v_0 = 0;
endmodule
module dmi_cdc (
	tck_i,
	trst_ni,
	jtag_dmi_req_i,
	jtag_dmi_ready_o,
	jtag_dmi_valid_i,
	jtag_dmi_cdc_clear_i,
	jtag_dmi_resp_o,
	jtag_dmi_valid_o,
	jtag_dmi_ready_i,
	clk_i,
	rst_ni,
	core_dmi_rst_no,
	core_dmi_req_o,
	core_dmi_valid_o,
	core_dmi_ready_i,
	core_dmi_resp_i,
	core_dmi_ready_o,
	core_dmi_valid_i
);
	// Trace: design.sv:46776:3
	input wire tck_i;
	// Trace: design.sv:46777:3
	input wire trst_ni;
	// Trace: design.sv:46778:3
	// removed localparam type dm_dtm_op_e
	// removed localparam type dm_dmi_req_t
	input wire [40:0] jtag_dmi_req_i;
	// Trace: design.sv:46779:3
	output wire jtag_dmi_ready_o;
	// Trace: design.sv:46780:3
	input wire jtag_dmi_valid_i;
	// Trace: design.sv:46781:3
	input wire jtag_dmi_cdc_clear_i;
	// Trace: design.sv:46785:3
	// removed localparam type dm_dmi_resp_t
	output wire [33:0] jtag_dmi_resp_o;
	// Trace: design.sv:46786:3
	output wire jtag_dmi_valid_o;
	// Trace: design.sv:46787:3
	input wire jtag_dmi_ready_i;
	// Trace: design.sv:46790:3
	input wire clk_i;
	// Trace: design.sv:46791:3
	input wire rst_ni;
	// Trace: design.sv:46793:3
	output wire core_dmi_rst_no;
	// Trace: design.sv:46794:3
	output wire [40:0] core_dmi_req_o;
	// Trace: design.sv:46795:3
	output wire core_dmi_valid_o;
	// Trace: design.sv:46796:3
	input wire core_dmi_ready_i;
	// Trace: design.sv:46798:3
	input wire [33:0] core_dmi_resp_i;
	// Trace: design.sv:46799:3
	output wire core_dmi_ready_o;
	// Trace: design.sv:46800:3
	input wire core_dmi_valid_i;
	// Trace: design.sv:46803:3
	wire core_clear_pending;
	// Trace: design.sv:46805:3
	cdc_2phase_clearable_88D17 i_cdc_req(
		.src_rst_ni(trst_ni),
		.src_clear_i(jtag_dmi_cdc_clear_i),
		.src_clk_i(tck_i),
		.src_clear_pending_o(),
		.src_data_i(jtag_dmi_req_i),
		.src_valid_i(jtag_dmi_valid_i),
		.src_ready_o(jtag_dmi_ready_o),
		.dst_rst_ni(rst_ni),
		.dst_clear_i(1'b0),
		.dst_clear_pending_o(core_clear_pending),
		.dst_clk_i(clk_i),
		.dst_data_o(core_dmi_req_o),
		.dst_valid_o(core_dmi_valid_o),
		.dst_ready_i(core_dmi_ready_i)
	);
	// Trace: design.sv:46827:3
	cdc_2phase_clearable_DC602 i_cdc_resp(
		.src_rst_ni(rst_ni),
		.src_clear_i(1'b0),
		.src_clear_pending_o(),
		.src_clk_i(clk_i),
		.src_data_i(core_dmi_resp_i),
		.src_valid_i(core_dmi_valid_i),
		.src_ready_o(core_dmi_ready_o),
		.dst_rst_ni(trst_ni),
		.dst_clear_i(jtag_dmi_cdc_clear_i),
		.dst_clear_pending_o(),
		.dst_clk_i(tck_i),
		.dst_data_o(jtag_dmi_resp_o),
		.dst_valid_o(jtag_dmi_valid_o),
		.dst_ready_i(jtag_dmi_ready_i)
	);
	// Trace: design.sv:46851:3
	reg core_clear_pending_q;
	// Trace: design.sv:46852:3
	reg core_dmi_rst_nq;
	// Trace: design.sv:46853:3
	wire clear_pending_rise_edge_detect;
	// Trace: design.sv:46855:3
	assign clear_pending_rise_edge_detect = !core_clear_pending_q && core_clear_pending;
	// Trace: design.sv:46857:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:46858:5
		if (!rst_ni) begin
			// Trace: design.sv:46859:7
			core_dmi_rst_nq <= 1'b1;
			// Trace: design.sv:46860:7
			core_clear_pending_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:46862:7
			core_dmi_rst_nq <= ~clear_pending_rise_edge_detect;
			// Trace: design.sv:46863:7
			core_clear_pending_q <= core_clear_pending;
		end
	// Trace: design.sv:46867:3
	assign core_dmi_rst_no = core_dmi_rst_nq;
endmodule
module dmi_jtag (
	clk_i,
	rst_ni,
	testmode_i,
	dmi_rst_no,
	dmi_req_o,
	dmi_req_valid_o,
	dmi_req_ready_i,
	dmi_resp_i,
	dmi_resp_ready_o,
	dmi_resp_valid_i,
	tck_i,
	tms_i,
	trst_ni,
	td_i,
	td_o,
	tdo_oe_o
);
	reg _sv2v_0;
	// Trace: design.sv:46889:13
	parameter [31:0] IdcodeValue = 32'h00000001;
	// Trace: design.sv:46891:3
	input wire clk_i;
	// Trace: design.sv:46892:3
	input wire rst_ni;
	// Trace: design.sv:46893:3
	input wire testmode_i;
	// Trace: design.sv:46897:3
	output wire dmi_rst_no;
	// Trace: design.sv:46898:3
	// removed localparam type dm_dtm_op_e
	// removed localparam type dm_dmi_req_t
	output wire [40:0] dmi_req_o;
	// Trace: design.sv:46899:3
	output wire dmi_req_valid_o;
	// Trace: design.sv:46900:3
	input wire dmi_req_ready_i;
	// Trace: design.sv:46902:3
	// removed localparam type dm_dmi_resp_t
	input wire [33:0] dmi_resp_i;
	// Trace: design.sv:46903:3
	output wire dmi_resp_ready_o;
	// Trace: design.sv:46904:3
	input wire dmi_resp_valid_i;
	// Trace: design.sv:46906:3
	input wire tck_i;
	// Trace: design.sv:46907:3
	input wire tms_i;
	// Trace: design.sv:46908:3
	input wire trst_ni;
	// Trace: design.sv:46909:3
	input wire td_i;
	// Trace: design.sv:46910:3
	output wire td_o;
	// Trace: design.sv:46911:3
	output wire tdo_oe_o;
	// Trace: design.sv:46914:3
	// removed localparam type dmi_error_e
	// Trace: design.sv:46918:3
	reg [1:0] error_d;
	reg [1:0] error_q;
	// Trace: design.sv:46920:3
	wire tck;
	// Trace: design.sv:46921:3
	wire jtag_dmi_clear;
	// Trace: design.sv:46923:3
	wire dmi_clear;
	// Trace: design.sv:46924:3
	wire update;
	// Trace: design.sv:46925:3
	wire capture;
	// Trace: design.sv:46926:3
	wire shift;
	// Trace: design.sv:46927:3
	wire tdi;
	// Trace: design.sv:46929:3
	wire dtmcs_select;
	// Trace: design.sv:46931:3
	// removed localparam type dm_dtmcs_t
	reg [31:0] dtmcs_q;
	assign dmi_clear = jtag_dmi_clear || ((dtmcs_select && update) && dtmcs_q[17]);
	// Trace: design.sv:46937:3
	reg [31:0] dtmcs_d;
	// Trace: design.sv:46939:3
	function automatic [30:0] sv2v_cast_31;
		input reg [30:0] inp;
		sv2v_cast_31 = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:46940:5
		dtmcs_d = dtmcs_q;
		// Trace: design.sv:46941:5
		if (capture) begin
			begin
				// Trace: design.sv:46942:7
				if (dtmcs_select)
					// Trace: design.sv:46943:9
					dtmcs_d = {20'h00001, error_q, 10'h071};
			end
		end
		if (shift) begin
			begin
				// Trace: design.sv:46957:7
				if (dtmcs_select)
					// Trace: design.sv:46957:25
					dtmcs_d = {tdi, sv2v_cast_31(dtmcs_q >> 1)};
			end
		end
	end
	// Trace: design.sv:46961:3
	always @(posedge tck or negedge trst_ni)
		// Trace: design.sv:46962:5
		if (!trst_ni)
			// Trace: design.sv:46963:7
			dtmcs_q <= 1'sb0;
		else
			// Trace: design.sv:46965:7
			dtmcs_q <= dtmcs_d;
	// Trace: design.sv:46973:3
	wire dmi_select;
	// Trace: design.sv:46974:3
	wire dmi_tdo;
	// Trace: design.sv:46976:3
	wire [40:0] dmi_req;
	// Trace: design.sv:46977:3
	wire dmi_req_ready;
	// Trace: design.sv:46978:3
	reg dmi_req_valid;
	// Trace: design.sv:46980:3
	wire [33:0] dmi_resp;
	// Trace: design.sv:46981:3
	wire dmi_resp_valid;
	// Trace: design.sv:46982:3
	wire dmi_resp_ready;
	// Trace: design.sv:46984:3
	// removed localparam type dmi_t
	// Trace: design.sv:46990:3
	// removed localparam type state_e
	// Trace: design.sv:46991:3
	reg [2:0] state_d;
	reg [2:0] state_q;
	// Trace: design.sv:46993:3
	reg [40:0] dr_d;
	reg [40:0] dr_q;
	// Trace: design.sv:46994:3
	reg [6:0] address_d;
	reg [6:0] address_q;
	// Trace: design.sv:46995:3
	reg [31:0] data_d;
	reg [31:0] data_q;
	// Trace: design.sv:46997:3
	wire [40:0] dmi;
	// Trace: design.sv:46998:3
	assign dmi = dr_q;
	// Trace: design.sv:46999:3
	assign dmi_req[40-:7] = address_q;
	// Trace: design.sv:47000:3
	assign dmi_req[31-:32] = data_q;
	// Trace: design.sv:47001:3
	assign dmi_req[33-:2] = (state_q == 3'd3 ? 2'h2 : 2'h1);
	// Trace: design.sv:47003:3
	assign dmi_resp_ready = 1'b1;
	// Trace: design.sv:47005:3
	reg error_dmi_busy;
	// Trace: design.sv:47007:3
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	always @(*) begin : p_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:47008:5
		error_dmi_busy = 1'b0;
		// Trace: design.sv:47010:5
		state_d = state_q;
		// Trace: design.sv:47011:5
		address_d = address_q;
		// Trace: design.sv:47012:5
		data_d = data_q;
		// Trace: design.sv:47013:5
		error_d = error_q;
		// Trace: design.sv:47015:5
		dmi_req_valid = 1'b0;
		// Trace: design.sv:47017:5
		if (dmi_clear) begin
			// Trace: design.sv:47018:7
			state_d = 3'd0;
			// Trace: design.sv:47019:7
			data_d = 1'sb0;
			// Trace: design.sv:47020:7
			error_d = 2'h0;
			// Trace: design.sv:47021:7
			address_d = 1'sb0;
		end
		else begin
			// Trace: design.sv:47023:7
			(* full_case, parallel_case *)
			case (state_q)
				3'd0:
					// Trace: design.sv:47026:11
					if ((dmi_select && update) && (error_q == 2'h0)) begin
						// Trace: design.sv:47028:13
						address_d = dmi[40-:7];
						// Trace: design.sv:47029:13
						data_d = dmi[33-:32];
						// Trace: design.sv:47030:13
						if (sv2v_cast_2(dmi[1-:2]) == 2'h1)
							// Trace: design.sv:47031:15
							state_d = 3'd1;
						else if (sv2v_cast_2(dmi[1-:2]) == 2'h2)
							// Trace: design.sv:47033:15
							state_d = 3'd3;
					end
				3'd1: begin
					// Trace: design.sv:47040:11
					dmi_req_valid = 1'b1;
					// Trace: design.sv:47041:11
					if (dmi_req_ready)
						// Trace: design.sv:47042:13
						state_d = 3'd2;
				end
				3'd2:
					// Trace: design.sv:47048:11
					if (dmi_resp_valid) begin
						// Trace: design.sv:47049:13
						data_d = dmi_resp[33-:32];
						// Trace: design.sv:47050:13
						state_d = 3'd0;
					end
				3'd3: begin
					// Trace: design.sv:47055:11
					dmi_req_valid = 1'b1;
					// Trace: design.sv:47057:11
					if (dmi_req_ready)
						// Trace: design.sv:47058:13
						state_d = 3'd4;
				end
				3'd4:
					// Trace: design.sv:47064:11
					if (dmi_resp_valid)
						// Trace: design.sv:47065:13
						state_d = 3'd0;
				default:
					// Trace: design.sv:47071:11
					if (dmi_resp_valid)
						// Trace: design.sv:47072:13
						state_d = 3'd0;
			endcase
			if (update && (state_q != 3'd0))
				// Trace: design.sv:47080:9
				error_dmi_busy = 1'b1;
			if (capture && |{state_q == 3'd1, state_q == 3'd2})
				// Trace: design.sv:47087:9
				error_dmi_busy = 1'b1;
			if (error_dmi_busy)
				// Trace: design.sv:47091:9
				error_d = 2'h3;
			if ((update && dtmcs_q[16]) && dtmcs_select)
				// Trace: design.sv:47095:9
				error_d = 2'h0;
		end
	end
	// Trace: design.sv:47101:3
	assign dmi_tdo = dr_q[0];
	// Trace: design.sv:47103:3
	always @(*) begin : p_shift
		if (_sv2v_0)
			;
		// Trace: design.sv:47104:5
		dr_d = dr_q;
		// Trace: design.sv:47105:5
		if (dmi_clear)
			// Trace: design.sv:47106:7
			dr_d = 1'sb0;
		else begin
			// Trace: design.sv:47108:7
			if (capture) begin
				begin
					// Trace: design.sv:47109:9
					if (dmi_select) begin
						begin
							// Trace: design.sv:47110:11
							if ((error_q == 2'h0) && !error_dmi_busy)
								// Trace: design.sv:47111:13
								dr_d = {address_q, data_q, 2'h0};
							else if ((error_q == 2'h3) || error_dmi_busy)
								// Trace: design.sv:47114:13
								dr_d = {address_q, data_q, 2'h3};
						end
					end
				end
			end
			if (shift) begin
				begin
					// Trace: design.sv:47120:9
					if (dmi_select)
						// Trace: design.sv:47121:11
						dr_d = {tdi, dr_q[40:1]};
				end
			end
		end
	end
	// Trace: design.sv:47127:3
	always @(posedge tck or negedge trst_ni)
		// Trace: design.sv:47128:5
		if (!trst_ni) begin
			// Trace: design.sv:47129:7
			dr_q <= 1'sb0;
			// Trace: design.sv:47130:7
			state_q <= 3'd0;
			// Trace: design.sv:47131:7
			address_q <= 1'sb0;
			// Trace: design.sv:47132:7
			data_q <= 1'sb0;
			// Trace: design.sv:47133:7
			error_q <= 2'h0;
		end
		else begin
			// Trace: design.sv:47135:7
			dr_q <= dr_d;
			// Trace: design.sv:47136:7
			state_q <= state_d;
			// Trace: design.sv:47137:7
			address_q <= address_d;
			// Trace: design.sv:47138:7
			data_q <= data_d;
			// Trace: design.sv:47139:7
			error_q <= error_d;
		end
	// Trace: design.sv:47146:3
	dmi_jtag_tap #(
		.IrLength(5),
		.IdcodeValue(IdcodeValue)
	) i_dmi_jtag_tap(
		.tck_i(tck_i),
		.tms_i(tms_i),
		.trst_ni(trst_ni),
		.td_i(td_i),
		.td_o(td_o),
		.tdo_oe_o(tdo_oe_o),
		.testmode_i(testmode_i),
		.tck_o(tck),
		.dmi_clear_o(jtag_dmi_clear),
		.update_o(update),
		.capture_o(capture),
		.shift_o(shift),
		.tdi_o(tdi),
		.dtmcs_select_o(dtmcs_select),
		.dtmcs_tdo_i(dtmcs_q[0]),
		.dmi_select_o(dmi_select),
		.dmi_tdo_i(dmi_tdo)
	);
	// Trace: design.sv:47172:3
	dmi_cdc i_dmi_cdc(
		.tck_i(tck),
		.trst_ni(trst_ni),
		.jtag_dmi_cdc_clear_i(dmi_clear),
		.jtag_dmi_req_i(dmi_req),
		.jtag_dmi_ready_o(dmi_req_ready),
		.jtag_dmi_valid_i(dmi_req_valid),
		.jtag_dmi_resp_o(dmi_resp),
		.jtag_dmi_valid_o(dmi_resp_valid),
		.jtag_dmi_ready_i(dmi_resp_ready),
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.core_dmi_rst_no(dmi_rst_no),
		.core_dmi_req_o(dmi_req_o),
		.core_dmi_valid_o(dmi_req_valid_o),
		.core_dmi_ready_i(dmi_req_ready_i),
		.core_dmi_resp_i(dmi_resp_i),
		.core_dmi_ready_o(dmi_resp_ready_o),
		.core_dmi_valid_i(dmi_resp_valid_i)
	);
	initial _sv2v_0 = 0;
endmodule
module dm_mem (
	clk_i,
	rst_ni,
	debug_req_o,
	hartsel_i,
	haltreq_i,
	resumereq_i,
	clear_resumeack_i,
	halted_o,
	resuming_o,
	progbuf_i,
	data_i,
	data_o,
	data_valid_o,
	cmd_valid_i,
	cmd_i,
	cmderror_valid_o,
	cmderror_o,
	cmdbusy_o,
	req_i,
	we_i,
	addr_i,
	wdata_i,
	be_i,
	rdata_o
);
	reg _sv2v_0;
	// Trace: design.sv:47215:13
	parameter [31:0] NrHarts = 1;
	// Trace: design.sv:47216:13
	parameter [31:0] BusWidth = 32;
	// Trace: design.sv:47217:13
	parameter [NrHarts - 1:0] SelectableHarts = {NrHarts {1'b1}};
	// Trace: design.sv:47218:13
	parameter [31:0] DmBaseAddress = 1'sb0;
	// Trace: design.sv:47220:3
	input wire clk_i;
	// Trace: design.sv:47221:3
	input wire rst_ni;
	// Trace: design.sv:47223:3
	output wire [NrHarts - 1:0] debug_req_o;
	// Trace: design.sv:47224:3
	input wire [19:0] hartsel_i;
	// Trace: design.sv:47226:3
	input wire [NrHarts - 1:0] haltreq_i;
	// Trace: design.sv:47227:3
	input wire [NrHarts - 1:0] resumereq_i;
	// Trace: design.sv:47228:3
	input wire clear_resumeack_i;
	// Trace: design.sv:47231:3
	output wire [NrHarts - 1:0] halted_o;
	// Trace: design.sv:47232:3
	output wire [NrHarts - 1:0] resuming_o;
	// Trace: design.sv:47234:3
	localparam [4:0] dm_ProgBufSize = 5'h08;
	input wire [255:0] progbuf_i;
	// Trace: design.sv:47236:3
	localparam [3:0] dm_DataCount = 4'h2;
	input wire [63:0] data_i;
	// Trace: design.sv:47237:3
	output reg [63:0] data_o;
	// Trace: design.sv:47238:3
	output reg data_valid_o;
	// Trace: design.sv:47240:3
	input wire cmd_valid_i;
	// Trace: design.sv:47241:3
	// removed localparam type dm_cmd_e
	// removed localparam type dm_command_t
	input wire [31:0] cmd_i;
	// Trace: design.sv:47242:3
	output reg cmderror_valid_o;
	// Trace: design.sv:47243:3
	// removed localparam type dm_cmderr_e
	output reg [2:0] cmderror_o;
	// Trace: design.sv:47244:3
	output reg cmdbusy_o;
	// Trace: design.sv:47248:3
	input wire req_i;
	// Trace: design.sv:47249:3
	input wire we_i;
	// Trace: design.sv:47250:3
	input wire [BusWidth - 1:0] addr_i;
	// Trace: design.sv:47251:3
	input wire [BusWidth - 1:0] wdata_i;
	// Trace: design.sv:47252:3
	input wire [(BusWidth / 8) - 1:0] be_i;
	// Trace: design.sv:47253:3
	output wire [BusWidth - 1:0] rdata_o;
	// Trace: design.sv:47255:3
	localparam [31:0] DbgAddressBits = 12;
	// Trace: design.sv:47256:3
	localparam [31:0] HartSelLen = (NrHarts == 1 ? 1 : $clog2(NrHarts));
	// Trace: design.sv:47257:3
	localparam [31:0] NrHartsAligned = 2 ** HartSelLen;
	// Trace: design.sv:47258:3
	localparam [31:0] MaxAar = (BusWidth == 64 ? 4 : 3);
	// Trace: design.sv:47259:3
	localparam [0:0] HasSndScratch = DmBaseAddress != 0;
	// Trace: design.sv:47261:3
	localparam [4:0] LoadBaseAddr = (DmBaseAddress == 0 ? 5'd0 : 5'd10);
	// Trace: design.sv:47263:3
	localparam [11:0] dm_DataAddr = 12'h380;
	localparam [11:0] DataBaseAddr = dm_DataAddr;
	// Trace: design.sv:47264:3
	localparam [11:0] DataEndAddr = 903;
	// Trace: design.sv:47265:3
	localparam [11:0] ProgBufBaseAddr = 864;
	// Trace: design.sv:47266:3
	localparam [11:0] ProgBufEndAddr = 895;
	// Trace: design.sv:47267:3
	localparam [11:0] AbstractCmdBaseAddr = ProgBufBaseAddr - 40;
	// Trace: design.sv:47268:3
	localparam [11:0] AbstractCmdEndAddr = ProgBufBaseAddr - 1;
	// Trace: design.sv:47270:3
	localparam [11:0] WhereToAddr = 'h300;
	// Trace: design.sv:47271:3
	localparam [11:0] FlagsBaseAddr = 'h400;
	// Trace: design.sv:47272:3
	localparam [11:0] FlagsEndAddr = 'h7ff;
	// Trace: design.sv:47274:3
	localparam [11:0] HaltedAddr = 'h100;
	// Trace: design.sv:47275:3
	localparam [11:0] GoingAddr = 'h104;
	// Trace: design.sv:47276:3
	localparam [11:0] ResumingAddr = 'h108;
	// Trace: design.sv:47277:3
	localparam [11:0] ExceptionAddr = 'h10c;
	// Trace: design.sv:47279:3
	wire [255:0] progbuf;
	// Trace: design.sv:47280:3
	reg [511:0] abstract_cmd;
	// Trace: design.sv:47281:3
	wire [NrHarts - 1:0] halted_d;
	reg [NrHarts - 1:0] halted_q;
	// Trace: design.sv:47282:3
	wire [NrHarts - 1:0] resuming_d;
	reg [NrHarts - 1:0] resuming_q;
	// Trace: design.sv:47283:3
	reg resume;
	reg go;
	reg going;
	// Trace: design.sv:47285:3
	reg exception;
	// Trace: design.sv:47286:3
	reg unsupported_command;
	// Trace: design.sv:47288:3
	wire [63:0] rom_rdata;
	// Trace: design.sv:47289:3
	reg [63:0] rdata_d;
	reg [63:0] rdata_q;
	// Trace: design.sv:47290:3
	reg word_enable32_q;
	// Trace: design.sv:47294:3
	wire [HartSelLen - 1:0] hartsel;
	wire [HartSelLen - 1:0] wdata_hartsel;
	// Trace: design.sv:47296:3
	assign hartsel = hartsel_i[HartSelLen - 1:0];
	// Trace: design.sv:47297:3
	assign wdata_hartsel = wdata_i[HartSelLen - 1:0];
	// Trace: design.sv:47299:3
	wire [NrHartsAligned - 1:0] resumereq_aligned;
	wire [NrHartsAligned - 1:0] haltreq_aligned;
	reg [NrHartsAligned - 1:0] halted_d_aligned;
	wire [NrHartsAligned - 1:0] halted_q_aligned;
	reg [NrHartsAligned - 1:0] halted_aligned;
	wire [NrHartsAligned - 1:0] resumereq_wdata_aligned;
	reg [NrHartsAligned - 1:0] resuming_d_aligned;
	wire [NrHartsAligned - 1:0] resuming_q_aligned;
	// Trace: design.sv:47304:3
	function automatic [NrHartsAligned - 1:0] sv2v_cast_DFF07;
		input reg [NrHartsAligned - 1:0] inp;
		sv2v_cast_DFF07 = inp;
	endfunction
	assign resumereq_aligned = sv2v_cast_DFF07(resumereq_i);
	// Trace: design.sv:47305:3
	assign haltreq_aligned = sv2v_cast_DFF07(haltreq_i);
	// Trace: design.sv:47306:3
	assign resumereq_wdata_aligned = sv2v_cast_DFF07(resumereq_i);
	// Trace: design.sv:47308:3
	assign halted_q_aligned = sv2v_cast_DFF07(halted_q);
	// Trace: design.sv:47309:3
	function automatic [NrHarts - 1:0] sv2v_cast_178F2;
		input reg [NrHarts - 1:0] inp;
		sv2v_cast_178F2 = inp;
	endfunction
	assign halted_d = sv2v_cast_178F2(halted_d_aligned);
	// Trace: design.sv:47310:3
	assign resuming_q_aligned = sv2v_cast_DFF07(resuming_q);
	// Trace: design.sv:47311:3
	assign resuming_d = sv2v_cast_178F2(resuming_d_aligned);
	// Trace: design.sv:47315:3
	wire fwd_rom_d;
	reg fwd_rom_q;
	// Trace: design.sv:47316:3
	// removed localparam type dm_ac_ar_cmd_t
	wire [23:0] ac_ar;
	// Trace: design.sv:47319:3
	function automatic [23:0] sv2v_cast_24;
		input reg [23:0] inp;
		sv2v_cast_24 = inp;
	endfunction
	assign ac_ar = sv2v_cast_24(cmd_i[23-:24]);
	// Trace: design.sv:47320:3
	assign debug_req_o = haltreq_i;
	// Trace: design.sv:47321:3
	assign halted_o = halted_q;
	// Trace: design.sv:47322:3
	assign resuming_o = resuming_q;
	// Trace: design.sv:47325:3
	assign progbuf = progbuf_i;
	// Trace: design.sv:47327:3
	// removed localparam type state_e
	// Trace: design.sv:47328:3
	reg [1:0] state_d;
	reg [1:0] state_q;
	// Trace: design.sv:47331:3
	always @(*) begin : p_hart_ctrl_queue
		if (_sv2v_0)
			;
		// Trace: design.sv:47332:5
		cmderror_valid_o = 1'b0;
		// Trace: design.sv:47333:5
		cmderror_o = 3'd0;
		// Trace: design.sv:47334:5
		state_d = state_q;
		// Trace: design.sv:47335:5
		go = 1'b0;
		// Trace: design.sv:47336:5
		resume = 1'b0;
		// Trace: design.sv:47337:5
		cmdbusy_o = 1'b1;
		// Trace: design.sv:47339:5
		(* full_case, parallel_case *)
		case (state_q)
			2'd0: begin
				// Trace: design.sv:47341:9
				cmdbusy_o = 1'b0;
				// Trace: design.sv:47342:9
				if ((cmd_valid_i && halted_q_aligned[hartsel]) && !unsupported_command)
					// Trace: design.sv:47344:11
					state_d = 2'd1;
				else if (cmd_valid_i) begin
					// Trace: design.sv:47347:11
					cmderror_valid_o = 1'b1;
					// Trace: design.sv:47348:11
					cmderror_o = 3'd4;
				end
				if (((resumereq_aligned[hartsel] && !resuming_q_aligned[hartsel]) && !haltreq_aligned[hartsel]) && halted_q_aligned[hartsel])
					// Trace: design.sv:47354:11
					state_d = 2'd2;
			end
			2'd1: begin
				// Trace: design.sv:47360:9
				cmdbusy_o = 1'b1;
				// Trace: design.sv:47361:9
				go = 1'b1;
				// Trace: design.sv:47363:9
				if (going)
					// Trace: design.sv:47364:13
					state_d = 2'd3;
			end
			2'd2: begin
				// Trace: design.sv:47369:9
				cmdbusy_o = 1'b1;
				// Trace: design.sv:47370:9
				resume = 1'b1;
				// Trace: design.sv:47371:9
				if (resuming_q_aligned[hartsel])
					// Trace: design.sv:47372:11
					state_d = 2'd0;
			end
			2'd3: begin
				// Trace: design.sv:47377:9
				cmdbusy_o = 1'b1;
				// Trace: design.sv:47378:9
				go = 1'b0;
				// Trace: design.sv:47380:9
				if (halted_aligned[hartsel])
					// Trace: design.sv:47381:11
					state_d = 2'd0;
			end
			default:
				;
		endcase
		if (unsupported_command && cmd_valid_i) begin
			// Trace: design.sv:47391:7
			cmderror_valid_o = 1'b1;
			// Trace: design.sv:47392:7
			cmderror_o = 3'd2;
		end
		if (exception) begin
			// Trace: design.sv:47396:7
			cmderror_valid_o = 1'b1;
			// Trace: design.sv:47397:7
			cmderror_o = 3'd3;
		end
	end
	// Trace: design.sv:47402:3
	wire [63:0] word_mux;
	// Trace: design.sv:47403:3
	assign word_mux = (fwd_rom_q ? rom_rdata : rdata_q);
	// Trace: design.sv:47405:3
	generate
		if (BusWidth == 64) begin : gen_word_mux64
			// Trace: design.sv:47406:5
			assign rdata_o = word_mux;
		end
		else begin : gen_word_mux32
			// Trace: design.sv:47408:5
			assign rdata_o = (word_enable32_q ? word_mux[32+:32] : word_mux[0+:32]);
		end
	endgenerate
	// Trace: design.sv:47412:3
	reg [63:0] data_bits;
	// Trace: design.sv:47413:3
	reg [63:0] rdata;
	// Trace: design.sv:47414:3
	localparam [63:0] dm_HaltAddress = 64'h0000000000000800;
	localparam [63:0] dm_ResumeAddress = 2052;
	function automatic [31:0] dm_jal;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:338:40
		input reg [4:0] rd;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:339:40
		input reg [20:0] imm;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:341:5
		dm_jal = {imm[20], imm[10:1], imm[11], imm[19:12], rd, 7'h6f};
	endfunction
	function automatic [20:0] sv2v_cast_21;
		input reg [20:0] inp;
		sv2v_cast_21 = inp;
	endfunction
	function automatic [$clog2(5'h08) - 1:0] sv2v_cast_63A1A;
		input reg [$clog2(5'h08) - 1:0] inp;
		sv2v_cast_63A1A = inp;
	endfunction
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [11:0] sv2v_cast_C1AAB;
		input reg [11:0] inp;
		sv2v_cast_C1AAB = inp;
	endfunction
	always @(*) begin : p_rw_logic
		if (_sv2v_0)
			;
		// Trace: design.sv:47416:5
		halted_d_aligned = sv2v_cast_DFF07(halted_q);
		// Trace: design.sv:47417:5
		resuming_d_aligned = sv2v_cast_DFF07(resuming_q);
		// Trace: design.sv:47418:5
		rdata_d = rdata_q;
		// Trace: design.sv:47420:5
		data_bits = data_i;
		// Trace: design.sv:47421:5
		rdata = 1'sb0;
		// Trace: design.sv:47424:5
		data_valid_o = 1'b0;
		// Trace: design.sv:47425:5
		exception = 1'b0;
		// Trace: design.sv:47426:5
		halted_aligned = 1'sb0;
		// Trace: design.sv:47427:5
		going = 1'b0;
		// Trace: design.sv:47430:5
		if (clear_resumeack_i)
			// Trace: design.sv:47431:7
			resuming_d_aligned[hartsel] = 1'b0;
		if (req_i) begin
			begin
				// Trace: design.sv:47436:7
				if (we_i) begin
					begin
						// Trace: design.sv:47437:9
						(* full_case, parallel_case *)
						if (addr_i[11:0] == HaltedAddr) begin
							// Trace: design.sv:47439:13
							halted_aligned[wdata_hartsel] = 1'b1;
							// Trace: design.sv:47440:13
							halted_d_aligned[wdata_hartsel] = 1'b1;
						end
						else if (addr_i[11:0] == GoingAddr)
							// Trace: design.sv:47443:13
							going = 1'b1;
						else if (addr_i[11:0] == ResumingAddr) begin
							// Trace: design.sv:47447:13
							halted_d_aligned[wdata_hartsel] = 1'b0;
							// Trace: design.sv:47449:13
							resuming_d_aligned[wdata_hartsel] = 1'b1;
						end
						else if (addr_i[11:0] == ExceptionAddr)
							// Trace: design.sv:47452:26
							exception = 1'b1;
						else if ((DataBaseAddr <= addr_i[11:0]) && (DataEndAddr >= addr_i[11:0])) begin
							// Trace: design.sv:47455:13
							data_valid_o = 1'b1;
							// Trace: design.sv:47456:13
							begin : sv2v_autoblock_1
								// Trace: design.sv:47456:18
								reg signed [31:0] i;
								// Trace: design.sv:47456:18
								for (i = 0; i < (BusWidth / 8); i = i + 1)
									begin
										// Trace: design.sv:47457:15
										if (be_i[i])
											// Trace: design.sv:47458:17
											data_bits[i * 8+:8] = wdata_i[i * 8+:8];
									end
							end
						end
					end
				end
				else
					// Trace: design.sv:47467:9
					(* full_case, parallel_case *)
					if (addr_i[11:0] == WhereToAddr) begin
						// Trace: design.sv:47471:13
						if (resumereq_wdata_aligned[wdata_hartsel])
							// Trace: design.sv:47472:15
							rdata_d = {32'b00000000000000000000000000000000, dm_jal(1'sb0, sv2v_cast_21(dm_ResumeAddress[11:0]) - sv2v_cast_21(WhereToAddr))};
						if (cmdbusy_o) begin
							begin
								// Trace: design.sv:47479:15
								if (((cmd_i[31-:8] == 8'h00) && !ac_ar[17]) && ac_ar[18])
									// Trace: design.sv:47481:17
									rdata_d = {32'b00000000000000000000000000000000, dm_jal(1'sb0, sv2v_cast_21(ProgBufBaseAddr) - sv2v_cast_21(WhereToAddr))};
								else
									// Trace: design.sv:47484:17
									rdata_d = {32'b00000000000000000000000000000000, dm_jal(1'sb0, sv2v_cast_21(AbstractCmdBaseAddr) - sv2v_cast_21(WhereToAddr))};
							end
						end
					end
					else if ((DataBaseAddr <= addr_i[11:0]) && (DataEndAddr >= addr_i[11:0]))
						// Trace: design.sv:47490:13
						rdata_d = {data_i[sv2v_cast_63A1A((addr_i[11:3] - DataBaseAddr[11:3]) + 1'b1) * 32+:32], data_i[sv2v_cast_63A1A(addr_i[11:3] - DataBaseAddr[11:3]) * 32+:32]};
					else if ((ProgBufBaseAddr <= addr_i[11:0]) && (ProgBufEndAddr >= addr_i[11:0]))
						// Trace: design.sv:47499:13
						rdata_d = progbuf[sv2v_cast_63A1A(addr_i[11:3] - ProgBufBaseAddr[11:3]) * 64+:64];
					else if ((AbstractCmdBaseAddr <= addr_i[11:0]) && (AbstractCmdEndAddr >= addr_i[11:0]))
						// Trace: design.sv:47506:13
						rdata_d = abstract_cmd[sv2v_cast_3(addr_i[11:3] - AbstractCmdBaseAddr[11:3]) * 64+:64];
					else if ((FlagsBaseAddr <= addr_i[11:0]) && (FlagsEndAddr >= addr_i[11:0])) begin
						// Trace: design.sv:47512:13
						if (({addr_i[11:3], 3'b000} - FlagsBaseAddr[11:0]) == (sv2v_cast_C1AAB(hartsel) & {{9 {1'b1}}, 3'b000}))
							// Trace: design.sv:47514:15
							rdata[(sv2v_cast_C1AAB(hartsel) & sv2v_cast_C1AAB(3'b111)) * 8+:8] = {6'b000000, resume, go};
						// Trace: design.sv:47516:13
						rdata_d = rdata;
					end
			end
		end
		// Trace: design.sv:47523:5
		data_o = data_bits;
	end
	// Trace: design.sv:47526:3
	// removed localparam type dm_csr_reg_t
	function automatic [31:0] dm_auipc;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:380:42
		input reg [4:0] rd;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:381:42
		input reg [20:0] imm;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:383:5
		dm_auipc = {imm[20], imm[10:1], imm[11], imm[19:12], rd, 7'h17};
	endfunction
	function automatic [31:0] dm_csrr;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:416:41
		input reg [11:0] csr;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:417:41
		input reg [4:0] dest;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:419:5
		dm_csrr = {csr, 8'h02, dest, 7'h73};
	endfunction
	function automatic [31:0] dm_csrw;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:410:41
		input reg [11:0] csr;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:411:41
		input reg [4:0] rs1;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:413:5
		dm_csrw = {csr, rs1, 15'h1073};
	endfunction
	function automatic [31:0] dm_ebreak;
		input reg _sv2v_unused;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:432:5
		dm_ebreak = 32'h00100073;
	endfunction
	function automatic [31:0] dm_float_load;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:394:47
		input reg [2:0] size;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:395:47
		input reg [4:0] dest;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:396:47
		input reg [4:0] base;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:397:47
		input reg [11:0] offset;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:399:5
		dm_float_load = {offset[11:0], base, size, dest, 7'b0000111};
	endfunction
	function automatic [31:0] dm_float_store;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:402:48
		input reg [2:0] size;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:403:48
		input reg [4:0] src;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:404:48
		input reg [4:0] base;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:405:48
		input reg [11:0] offset;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:407:5
		dm_float_store = {offset[11:5], src, base, size, offset[4:0], 7'b0100111};
	endfunction
	function automatic [31:0] dm_illegal;
		input reg _sv2v_unused;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:444:5
		dm_illegal = 32'h00000000;
	endfunction
	function automatic [31:0] dm_load;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:372:41
		input reg [2:0] size;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:373:41
		input reg [4:0] dest;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:374:41
		input reg [4:0] base;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:375:41
		input reg [11:0] offset;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:377:5
		dm_load = {offset[11:0], base, size, dest, 7'h03};
	endfunction
	function automatic [31:0] dm_nop;
		input reg _sv2v_unused;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:440:5
		dm_nop = 32'h00000013;
	endfunction
	function automatic [31:0] dm_slli;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:358:41
		input reg [4:0] rd;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:359:41
		input reg [4:0] rs1;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:360:41
		input reg [5:0] shamt;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:362:5
		dm_slli = {6'b000000, shamt[5:0], rs1, 3'h1, rd, 7'h13};
	endfunction
	function automatic [31:0] dm_srli;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:365:41
		input reg [4:0] rd;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:366:41
		input reg [4:0] rs1;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:367:41
		input reg [5:0] shamt;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:369:5
		dm_srli = {6'b000000, shamt[5:0], rs1, 3'h5, rd, 7'h13};
	endfunction
	function automatic [31:0] dm_store;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:386:42
		input reg [2:0] size;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:387:42
		input reg [4:0] src;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:388:42
		input reg [4:0] base;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:389:42
		input reg [11:0] offset;
		// Trace: ../src/pulp-platform.org__riscv_dbg_pkg_0/pulp_platform_riscv_dbg/src/dm_pkg.sv:391:5
		dm_store = {offset[11:5], src, base, size, offset[4:0], 7'h23};
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	always @(*) begin : p_abstract_cmd_rom
		if (_sv2v_0)
			;
		// Trace: design.sv:47528:5
		unsupported_command = 1'b0;
		// Trace: design.sv:47531:5
		abstract_cmd[31-:32] = dm_illegal(0);
		// Trace: design.sv:47533:5
		abstract_cmd[63-:32] = (HasSndScratch ? dm_auipc(5'd10, 1'sb0) : dm_nop(0));
		// Trace: design.sv:47535:5
		abstract_cmd[95-:32] = (HasSndScratch ? dm_srli(5'd10, 5'd10, 6'd12) : dm_nop(0));
		// Trace: design.sv:47536:5
		abstract_cmd[127-:32] = (HasSndScratch ? dm_slli(5'd10, 5'd10, 6'd12) : dm_nop(0));
		// Trace: design.sv:47537:5
		abstract_cmd[159-:32] = dm_nop(0);
		// Trace: design.sv:47538:5
		abstract_cmd[191-:32] = dm_nop(0);
		// Trace: design.sv:47539:5
		abstract_cmd[223-:32] = dm_nop(0);
		// Trace: design.sv:47540:5
		abstract_cmd[255-:32] = dm_nop(0);
		// Trace: design.sv:47541:5
		abstract_cmd[287-:32] = (HasSndScratch ? dm_csrr(12'h7b3, 5'd10) : dm_nop(0));
		// Trace: design.sv:47542:5
		abstract_cmd[319-:32] = dm_ebreak(0);
		// Trace: design.sv:47543:5
		abstract_cmd[320+:192] = 1'sb0;
		// Trace: design.sv:47546:5
		(* full_case, parallel_case *)
		case (cmd_i[31-:8])
			8'h00: begin
				// Trace: design.sv:47551:9
				if (((sv2v_cast_32(ac_ar[22-:3]) < MaxAar) && ac_ar[17]) && ac_ar[16]) begin
					// Trace: design.sv:47553:11
					abstract_cmd[31-:32] = (HasSndScratch ? dm_csrw(12'h7b3, 5'd10) : dm_nop(0));
					// Trace: design.sv:47555:11
					if (ac_ar[15:14] != {2 {1'sb0}}) begin
						// Trace: design.sv:47556:13
						abstract_cmd[31-:32] = dm_ebreak(0);
						// Trace: design.sv:47557:13
						unsupported_command = 1'b1;
					end
					else if (((HasSndScratch && ac_ar[12]) && !ac_ar[5]) && (ac_ar[4:0] == 5'd10)) begin
						// Trace: design.sv:47563:13
						abstract_cmd[159-:32] = dm_csrw(12'h7b2, 5'd8);
						// Trace: design.sv:47565:13
						abstract_cmd[191-:32] = dm_load(ac_ar[22-:3], 5'd8, LoadBaseAddr, dm_DataAddr);
						// Trace: design.sv:47567:13
						abstract_cmd[223-:32] = dm_csrw(12'h7b3, 5'd8);
						// Trace: design.sv:47569:13
						abstract_cmd[255-:32] = dm_csrr(12'h7b2, 5'd8);
					end
					else if (ac_ar[12]) begin
						begin
							// Trace: design.sv:47573:13
							if (ac_ar[5])
								// Trace: design.sv:47574:15
								abstract_cmd[159-:32] = dm_float_load(ac_ar[22-:3], ac_ar[4:0], LoadBaseAddr, dm_DataAddr);
							else
								// Trace: design.sv:47577:15
								abstract_cmd[159-:32] = dm_load(ac_ar[22-:3], ac_ar[4:0], LoadBaseAddr, dm_DataAddr);
						end
					end
					else begin
						// Trace: design.sv:47584:13
						abstract_cmd[159-:32] = dm_csrw(12'h7b2, 5'd8);
						// Trace: design.sv:47586:13
						abstract_cmd[191-:32] = dm_load(ac_ar[22-:3], 5'd8, LoadBaseAddr, dm_DataAddr);
						// Trace: design.sv:47588:13
						abstract_cmd[223-:32] = dm_csrw(ac_ar[11:0], 5'd8);
						// Trace: design.sv:47590:13
						abstract_cmd[255-:32] = dm_csrr(12'h7b2, 5'd8);
					end
				end
				else if (((sv2v_cast_32(ac_ar[22-:3]) < MaxAar) && ac_ar[17]) && !ac_ar[16]) begin
					// Trace: design.sv:47594:11
					abstract_cmd[31-:32] = (HasSndScratch ? dm_csrw(12'h7b3, LoadBaseAddr) : dm_nop(0));
					// Trace: design.sv:47598:11
					if (ac_ar[15:14] != {2 {1'sb0}}) begin
						// Trace: design.sv:47599:15
						abstract_cmd[31-:32] = dm_ebreak(0);
						// Trace: design.sv:47600:15
						unsupported_command = 1'b1;
					end
					else if (((HasSndScratch && ac_ar[12]) && !ac_ar[5]) && (ac_ar[4:0] == 5'd10)) begin
						// Trace: design.sv:47606:13
						abstract_cmd[159-:32] = dm_csrw(12'h7b2, 5'd8);
						// Trace: design.sv:47608:13
						abstract_cmd[191-:32] = dm_csrr(12'h7b3, 5'd8);
						// Trace: design.sv:47610:13
						abstract_cmd[223-:32] = dm_store(ac_ar[22-:3], 5'd8, LoadBaseAddr, dm_DataAddr);
						// Trace: design.sv:47612:13
						abstract_cmd[255-:32] = dm_csrr(12'h7b2, 5'd8);
					end
					else if (ac_ar[12]) begin
						begin
							// Trace: design.sv:47616:13
							if (ac_ar[5])
								// Trace: design.sv:47617:15
								abstract_cmd[159-:32] = dm_float_store(ac_ar[22-:3], ac_ar[4:0], LoadBaseAddr, dm_DataAddr);
							else
								// Trace: design.sv:47620:15
								abstract_cmd[159-:32] = dm_store(ac_ar[22-:3], ac_ar[4:0], LoadBaseAddr, dm_DataAddr);
						end
					end
					else begin
						// Trace: design.sv:47627:13
						abstract_cmd[159-:32] = dm_csrw(12'h7b2, 5'd8);
						// Trace: design.sv:47629:13
						abstract_cmd[191-:32] = dm_csrr(ac_ar[11:0], 5'd8);
						// Trace: design.sv:47631:13
						abstract_cmd[223-:32] = dm_store(ac_ar[22-:3], 5'd8, LoadBaseAddr, dm_DataAddr);
						// Trace: design.sv:47633:13
						abstract_cmd[255-:32] = dm_csrr(12'h7b2, 5'd8);
					end
				end
				else if ((sv2v_cast_32(ac_ar[22-:3]) >= MaxAar) || (ac_ar[19] == 1'b1)) begin
					// Trace: design.sv:47639:11
					abstract_cmd[31-:32] = dm_ebreak(0);
					// Trace: design.sv:47640:11
					unsupported_command = 1'b1;
				end
				if (ac_ar[18] && !unsupported_command)
					// Trace: design.sv:47649:11
					abstract_cmd[319-:32] = dm_nop(0);
			end
			default: begin
				// Trace: design.sv:47656:9
				abstract_cmd[31-:32] = dm_ebreak(0);
				// Trace: design.sv:47657:9
				unsupported_command = 1'b1;
			end
		endcase
	end
	// Trace: design.sv:47662:3
	wire [63:0] rom_addr;
	// Trace: design.sv:47663:3
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	assign rom_addr = sv2v_cast_64(addr_i);
	// Trace: design.sv:47671:3
	generate
		if (HasSndScratch) begin : gen_rom_snd_scratch
			// Trace: design.sv:47672:5
			debug_rom i_debug_rom(
				.clk_i(clk_i),
				.req_i(req_i),
				.addr_i(rom_addr),
				.rdata_o(rom_rdata)
			);
		end
		else begin : gen_rom_one_scratch
			// Trace: design.sv:47682:5
			debug_rom_one_scratch i_debug_rom(
				.clk_i(clk_i),
				.req_i(req_i),
				.addr_i(rom_addr),
				.rdata_o(rom_rdata)
			);
		end
	endgenerate
	// Trace: design.sv:47692:3
	assign fwd_rom_d = addr_i[11:0] >= dm_HaltAddress[11:0];
	// Trace: design.sv:47694:3
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:47695:5
		if (!rst_ni) begin
			// Trace: design.sv:47696:7
			fwd_rom_q <= 1'b0;
			// Trace: design.sv:47697:7
			rdata_q <= 1'sb0;
			// Trace: design.sv:47698:7
			state_q <= 2'd0;
			// Trace: design.sv:47699:7
			word_enable32_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:47701:7
			fwd_rom_q <= fwd_rom_d;
			// Trace: design.sv:47702:7
			rdata_q <= rdata_d;
			// Trace: design.sv:47703:7
			state_q <= state_d;
			// Trace: design.sv:47704:7
			word_enable32_q <= addr_i[2];
		end
	end
	// Trace: design.sv:47708:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:47709:5
		if (!rst_ni) begin
			// Trace: design.sv:47710:7
			halted_q <= 1'b0;
			// Trace: design.sv:47711:7
			resuming_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:47713:7
			halted_q <= SelectableHarts & halted_d;
			// Trace: design.sv:47714:7
			resuming_q <= SelectableHarts & resuming_d;
		end
	initial _sv2v_0 = 0;
endmodule
module dm_obi_top (
	clk_i,
	rst_ni,
	testmode_i,
	ndmreset_o,
	dmactive_o,
	debug_req_o,
	unavailable_i,
	hartinfo_i,
	slave_req_i,
	slave_gnt_o,
	slave_we_i,
	slave_addr_i,
	slave_be_i,
	slave_wdata_i,
	slave_aid_i,
	slave_rvalid_o,
	slave_rdata_o,
	slave_rid_o,
	master_req_o,
	master_addr_o,
	master_we_o,
	master_wdata_o,
	master_be_o,
	master_gnt_i,
	master_rvalid_i,
	master_err_i,
	master_other_err_i,
	master_rdata_i,
	dmi_rst_ni,
	dmi_req_valid_i,
	dmi_req_ready_o,
	dmi_req_i,
	dmi_resp_valid_o,
	dmi_resp_ready_i,
	dmi_resp_o
);
	// Trace: design.sv:47782:13
	parameter [31:0] IdWidth = 1;
	// Trace: design.sv:47783:13
	parameter [31:0] NrHarts = 1;
	// Trace: design.sv:47784:13
	parameter [31:0] BusWidth = 32;
	// Trace: design.sv:47785:13
	parameter [31:0] DmBaseAddress = 'h1000;
	// Trace: design.sv:47788:13
	parameter [NrHarts - 1:0] SelectableHarts = {NrHarts {1'b1}};
	// Trace: design.sv:47790:3
	input wire clk_i;
	// Trace: design.sv:47792:3
	input wire rst_ni;
	// Trace: design.sv:47793:3
	input wire testmode_i;
	// Trace: design.sv:47794:3
	output wire ndmreset_o;
	// Trace: design.sv:47795:3
	output wire dmactive_o;
	// Trace: design.sv:47796:3
	output wire [NrHarts - 1:0] debug_req_o;
	// Trace: design.sv:47798:3
	input wire [NrHarts - 1:0] unavailable_i;
	// Trace: design.sv:47799:3
	// removed localparam type dm_hartinfo_t
	input wire [(NrHarts * 32) - 1:0] hartinfo_i;
	// Trace: design.sv:47801:3
	input wire slave_req_i;
	// Trace: design.sv:47803:3
	output wire slave_gnt_o;
	// Trace: design.sv:47804:3
	input wire slave_we_i;
	// Trace: design.sv:47805:3
	input wire [BusWidth - 1:0] slave_addr_i;
	// Trace: design.sv:47806:3
	input wire [(BusWidth / 8) - 1:0] slave_be_i;
	// Trace: design.sv:47807:3
	input wire [BusWidth - 1:0] slave_wdata_i;
	// Trace: design.sv:47809:3
	input wire [IdWidth - 1:0] slave_aid_i;
	// Trace: design.sv:47811:3
	output wire slave_rvalid_o;
	// Trace: design.sv:47812:3
	output wire [BusWidth - 1:0] slave_rdata_o;
	// Trace: design.sv:47814:3
	output wire [IdWidth - 1:0] slave_rid_o;
	// Trace: design.sv:47816:3
	output wire master_req_o;
	// Trace: design.sv:47817:3
	output wire [BusWidth - 1:0] master_addr_o;
	// Trace: design.sv:47818:3
	output wire master_we_o;
	// Trace: design.sv:47819:3
	output wire [BusWidth - 1:0] master_wdata_o;
	// Trace: design.sv:47820:3
	output wire [(BusWidth / 8) - 1:0] master_be_o;
	// Trace: design.sv:47821:3
	input wire master_gnt_i;
	// Trace: design.sv:47822:3
	input wire master_rvalid_i;
	// Trace: design.sv:47823:3
	input wire master_err_i;
	// Trace: design.sv:47824:3
	input wire master_other_err_i;
	// Trace: design.sv:47825:3
	input wire [BusWidth - 1:0] master_rdata_i;
	// Trace: design.sv:47828:3
	input wire dmi_rst_ni;
	// Trace: design.sv:47829:3
	input wire dmi_req_valid_i;
	// Trace: design.sv:47830:3
	output wire dmi_req_ready_o;
	// Trace: design.sv:47831:3
	// removed localparam type dm_dtm_op_e
	// removed localparam type dm_dmi_req_t
	input wire [40:0] dmi_req_i;
	// Trace: design.sv:47833:3
	output wire dmi_resp_valid_o;
	// Trace: design.sv:47834:3
	input wire dmi_resp_ready_i;
	// Trace: design.sv:47835:3
	// removed localparam type dm_dmi_resp_t
	output wire [33:0] dmi_resp_o;
	// Trace: design.sv:47839:3
	reg slave_rvalid_q;
	// Trace: design.sv:47840:3
	reg [IdWidth - 1:0] slave_rid_q;
	// Trace: design.sv:47843:3
	dm_top #(
		.NrHarts(NrHarts),
		.BusWidth(BusWidth),
		.DmBaseAddress(DmBaseAddress),
		.SelectableHarts(SelectableHarts)
	) i_dm_top(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.testmode_i(testmode_i),
		.ndmreset_o(ndmreset_o),
		.dmactive_o(dmactive_o),
		.debug_req_o(debug_req_o),
		.unavailable_i(unavailable_i),
		.hartinfo_i(hartinfo_i),
		.slave_req_i(slave_req_i),
		.slave_we_i(slave_we_i),
		.slave_addr_i(slave_addr_i),
		.slave_be_i(slave_be_i),
		.slave_wdata_i(slave_wdata_i),
		.slave_rdata_o(slave_rdata_o),
		.master_req_o(master_req_o),
		.master_add_o(master_addr_o),
		.master_we_o(master_we_o),
		.master_wdata_o(master_wdata_o),
		.master_be_o(master_be_o),
		.master_gnt_i(master_gnt_i),
		.master_r_valid_i(master_rvalid_i),
		.master_r_err_i(master_err_i),
		.master_r_other_err_i(master_other_err_i),
		.master_r_rdata_i(master_rdata_i),
		.dmi_rst_ni(dmi_rst_ni),
		.dmi_req_valid_i(dmi_req_valid_i),
		.dmi_req_ready_o(dmi_req_ready_o),
		.dmi_req_i(dmi_req_i),
		.dmi_resp_valid_o(dmi_resp_valid_o),
		.dmi_resp_ready_i(dmi_resp_ready_i),
		.dmi_resp_o(dmi_resp_o)
	);
	// Trace: design.sv:47891:3
	always @(posedge clk_i or negedge rst_ni) begin : obi_regs
		// Trace: design.sv:47892:5
		if (!rst_ni) begin
			// Trace: design.sv:47893:7
			slave_rvalid_q <= 1'b0;
			// Trace: design.sv:47894:7
			slave_rid_q <= 'b0;
		end
		else
			// Trace: design.sv:47896:7
			if (slave_req_i && slave_gnt_o) begin
				// Trace: design.sv:47897:9
				slave_rvalid_q <= 1'b1;
				// Trace: design.sv:47898:9
				slave_rid_q <= slave_aid_i;
			end
			else
				// Trace: design.sv:47900:9
				slave_rvalid_q <= 1'b0;
	end
	// Trace: design.sv:47905:3
	assign slave_gnt_o = 1'b1;
	// Trace: design.sv:47906:3
	assign slave_rvalid_o = slave_rvalid_q;
	// Trace: design.sv:47907:3
	assign slave_rid_o = slave_rid_q;
endmodule
module dm_sba (
	clk_i,
	rst_ni,
	dmactive_i,
	master_req_o,
	master_add_o,
	master_we_o,
	master_wdata_o,
	master_be_o,
	master_gnt_i,
	master_r_valid_i,
	master_r_err_i,
	master_r_other_err_i,
	master_r_rdata_i,
	sbaddress_i,
	sbaddress_write_valid_i,
	sbreadonaddr_i,
	sbaddress_o,
	sbautoincrement_i,
	sbaccess_i,
	sbreadondata_i,
	sbdata_i,
	sbdata_read_valid_i,
	sbdata_write_valid_i,
	sbdata_o,
	sbdata_valid_o,
	sbbusy_o,
	sberror_valid_o,
	sberror_o
);
	reg _sv2v_0;
	// Trace: design.sv:47928:13
	parameter [31:0] BusWidth = 32;
	// Trace: design.sv:47929:13
	parameter [0:0] ReadByteEnable = 1;
	// Trace: design.sv:47931:3
	input wire clk_i;
	// Trace: design.sv:47932:3
	input wire rst_ni;
	// Trace: design.sv:47933:3
	input wire dmactive_i;
	// Trace: design.sv:47935:3
	output wire master_req_o;
	// Trace: design.sv:47936:3
	output wire [BusWidth - 1:0] master_add_o;
	// Trace: design.sv:47937:3
	output wire master_we_o;
	// Trace: design.sv:47938:3
	output wire [BusWidth - 1:0] master_wdata_o;
	// Trace: design.sv:47939:3
	output wire [(BusWidth / 8) - 1:0] master_be_o;
	// Trace: design.sv:47940:3
	input wire master_gnt_i;
	// Trace: design.sv:47941:3
	input wire master_r_valid_i;
	// Trace: design.sv:47942:3
	input wire master_r_err_i;
	// Trace: design.sv:47943:3
	input wire master_r_other_err_i;
	// Trace: design.sv:47944:3
	input wire [BusWidth - 1:0] master_r_rdata_i;
	// Trace: design.sv:47946:3
	input wire [BusWidth - 1:0] sbaddress_i;
	// Trace: design.sv:47947:3
	input wire sbaddress_write_valid_i;
	// Trace: design.sv:47949:3
	input wire sbreadonaddr_i;
	// Trace: design.sv:47950:3
	output wire [BusWidth - 1:0] sbaddress_o;
	// Trace: design.sv:47951:3
	input wire sbautoincrement_i;
	// Trace: design.sv:47952:3
	input wire [2:0] sbaccess_i;
	// Trace: design.sv:47954:3
	input wire sbreadondata_i;
	// Trace: design.sv:47955:3
	input wire [BusWidth - 1:0] sbdata_i;
	// Trace: design.sv:47956:3
	input wire sbdata_read_valid_i;
	// Trace: design.sv:47957:3
	input wire sbdata_write_valid_i;
	// Trace: design.sv:47959:3
	output wire [BusWidth - 1:0] sbdata_o;
	// Trace: design.sv:47960:3
	output wire sbdata_valid_o;
	// Trace: design.sv:47962:3
	output wire sbbusy_o;
	// Trace: design.sv:47963:3
	output reg sberror_valid_o;
	// Trace: design.sv:47964:3
	output reg [2:0] sberror_o;
	// Trace: design.sv:47967:3
	localparam signed [31:0] BeIdxWidth = $clog2(BusWidth / 8);
	// Trace: design.sv:47968:3
	// removed localparam type dm_sba_state_e
	reg [2:0] state_d;
	reg [2:0] state_q;
	// Trace: design.sv:47970:3
	reg [BusWidth - 1:0] address;
	// Trace: design.sv:47971:3
	reg req;
	// Trace: design.sv:47972:3
	wire gnt;
	// Trace: design.sv:47973:3
	reg we;
	// Trace: design.sv:47974:3
	reg [(BusWidth / 8) - 1:0] be;
	// Trace: design.sv:47975:3
	reg [(BusWidth / 8) - 1:0] be_mask;
	// Trace: design.sv:47976:3
	reg [BeIdxWidth - 1:0] be_idx;
	// Trace: design.sv:47978:3
	assign sbbusy_o = state_q != 3'd0;
	// Trace: design.sv:47980:3
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	always @(*) begin : p_be_mask
		if (_sv2v_0)
			;
		// Trace: design.sv:47981:5
		be_mask = 1'sb0;
		// Trace: design.sv:47984:5
		(* full_case, parallel_case *)
		case (sbaccess_i)
			3'b000:
				// Trace: design.sv:47986:9
				be_mask[be_idx] = 1'sb1;
			3'b001:
				// Trace: design.sv:47989:9
				be_mask[sv2v_cast_32_signed({be_idx[BeIdxWidth - 1:1], 1'b0})+:2] = 1'sb1;
			3'b010:
				// Trace: design.sv:47992:9
				if (BusWidth == 32'd64)
					// Trace: design.sv:47992:33
					be_mask[sv2v_cast_32_signed({be_idx[BeIdxWidth - 1], 2'h0})+:4] = 1'sb1;
				else
					// Trace: design.sv:47993:33
					be_mask = 1'sb1;
			3'b011:
				// Trace: design.sv:47995:15
				be_mask = 1'sb1;
			default:
				;
		endcase
	end
	// Trace: design.sv:48000:3
	wire [BusWidth - 1:0] sbaccess_mask;
	// Trace: design.sv:48001:3
	assign sbaccess_mask = {BusWidth {1'b1}} << sbaccess_i;
	// Trace: design.sv:48003:3
	reg addr_incr_en;
	// Trace: design.sv:48004:3
	wire [BusWidth - 1:0] addr_incr;
	// Trace: design.sv:48005:3
	function automatic [BusWidth - 1:0] sv2v_cast_8CBFF;
		input reg [BusWidth - 1:0] inp;
		sv2v_cast_8CBFF = inp;
	endfunction
	assign addr_incr = (addr_incr_en ? sv2v_cast_8CBFF(1'b1) << sbaccess_i : {BusWidth {1'sb0}});
	// Trace: design.sv:48006:3
	assign sbaddress_o = sbaddress_i + addr_incr;
	// Trace: design.sv:48009:3
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	always @(*) begin : p_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:48010:5
		req = 1'b0;
		// Trace: design.sv:48011:5
		address = sbaddress_i;
		// Trace: design.sv:48012:5
		we = 1'b0;
		// Trace: design.sv:48013:5
		be = 1'sb0;
		// Trace: design.sv:48014:5
		be_idx = sbaddress_i[BeIdxWidth - 1:0];
		// Trace: design.sv:48016:5
		sberror_o = 1'sb0;
		// Trace: design.sv:48017:5
		sberror_valid_o = 1'b0;
		// Trace: design.sv:48019:5
		addr_incr_en = 1'b0;
		// Trace: design.sv:48021:5
		state_d = state_q;
		// Trace: design.sv:48023:5
		(* full_case, parallel_case *)
		case (state_q)
			3'd0: begin
				// Trace: design.sv:48026:9
				if (sbaddress_write_valid_i && sbreadonaddr_i)
					// Trace: design.sv:48026:57
					state_d = 3'd1;
				if (sbdata_write_valid_i)
					// Trace: design.sv:48028:35
					state_d = 3'd2;
				if (sbdata_read_valid_i && sbreadondata_i)
					// Trace: design.sv:48030:52
					state_d = 3'd1;
			end
			3'd1: begin
				// Trace: design.sv:48034:9
				req = 1'b1;
				// Trace: design.sv:48035:9
				if (ReadByteEnable)
					// Trace: design.sv:48035:29
					be = be_mask;
				if (gnt)
					// Trace: design.sv:48036:18
					state_d = 3'd3;
			end
			3'd2: begin
				// Trace: design.sv:48040:9
				req = 1'b1;
				// Trace: design.sv:48041:9
				we = 1'b1;
				// Trace: design.sv:48042:9
				be = be_mask;
				// Trace: design.sv:48043:9
				if (gnt)
					// Trace: design.sv:48043:18
					state_d = 3'd4;
			end
			3'd3:
				// Trace: design.sv:48047:9
				if (sbdata_valid_o) begin
					// Trace: design.sv:48048:11
					state_d = 3'd0;
					// Trace: design.sv:48050:11
					addr_incr_en = sbautoincrement_i;
					// Trace: design.sv:48052:11
					if (master_r_other_err_i) begin
						// Trace: design.sv:48053:13
						sberror_valid_o = 1'b1;
						// Trace: design.sv:48054:13
						sberror_o = 3'd7;
					end
					else if (master_r_err_i) begin
						// Trace: design.sv:48057:13
						sberror_valid_o = 1'b1;
						// Trace: design.sv:48058:13
						sberror_o = 3'd2;
					end
				end
			3'd4:
				// Trace: design.sv:48064:9
				if (sbdata_valid_o) begin
					// Trace: design.sv:48065:11
					state_d = 3'd0;
					// Trace: design.sv:48067:11
					addr_incr_en = sbautoincrement_i;
					// Trace: design.sv:48069:11
					if (master_r_other_err_i) begin
						// Trace: design.sv:48070:13
						sberror_valid_o = 1'b1;
						// Trace: design.sv:48071:13
						sberror_o = 3'd7;
					end
					else if (master_r_err_i) begin
						// Trace: design.sv:48074:13
						sberror_valid_o = 1'b1;
						// Trace: design.sv:48075:13
						sberror_o = 3'd2;
					end
				end
			default:
				// Trace: design.sv:48080:16
				state_d = 3'd0;
		endcase
		if ((sv2v_cast_32(sbaccess_i) > BeIdxWidth) && (state_q != 3'd0)) begin
			// Trace: design.sv:48085:7
			req = 1'b0;
			// Trace: design.sv:48086:7
			state_d = 3'd0;
			// Trace: design.sv:48087:7
			sberror_valid_o = 1'b1;
			// Trace: design.sv:48088:7
			sberror_o = 3'd4;
		end
		if (|(sbaddress_i & ~sbaccess_mask) && (state_q != 3'd0)) begin
			// Trace: design.sv:48093:7
			req = 1'b0;
			// Trace: design.sv:48094:7
			state_d = 3'd0;
			// Trace: design.sv:48095:7
			sberror_valid_o = 1'b1;
			// Trace: design.sv:48096:7
			sberror_o = 3'd3;
		end
	end
	// Trace: design.sv:48101:3
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:48102:5
		if (!rst_ni)
			// Trace: design.sv:48103:7
			state_q <= 3'd0;
		else
			// Trace: design.sv:48105:7
			state_q <= state_d;
	end
	// Trace: design.sv:48109:3
	wire [BeIdxWidth - 1:0] be_idx_masked;
	// Trace: design.sv:48110:3
	function automatic [BeIdxWidth - 1:0] sv2v_cast_F03CB;
		input reg [BeIdxWidth - 1:0] inp;
		sv2v_cast_F03CB = inp;
	endfunction
	assign be_idx_masked = be_idx & sv2v_cast_F03CB(sbaccess_mask);
	// Trace: design.sv:48111:3
	assign master_req_o = req;
	// Trace: design.sv:48112:3
	assign master_add_o = address[BusWidth - 1:0];
	// Trace: design.sv:48113:3
	assign master_we_o = we;
	// Trace: design.sv:48114:3
	assign master_wdata_o = sbdata_i[BusWidth - 1:0] << (8 * be_idx_masked);
	// Trace: design.sv:48115:3
	assign master_be_o = be[(BusWidth / 8) - 1:0];
	// Trace: design.sv:48116:3
	assign gnt = master_gnt_i;
	// Trace: design.sv:48117:3
	assign sbdata_valid_o = master_r_valid_i;
	// Trace: design.sv:48118:3
	assign sbdata_o = master_r_rdata_i[BusWidth - 1:0] >> (8 * be_idx_masked);
	initial _sv2v_0 = 0;
endmodule
module dm_top (
	clk_i,
	rst_ni,
	testmode_i,
	ndmreset_o,
	dmactive_o,
	debug_req_o,
	unavailable_i,
	hartinfo_i,
	slave_req_i,
	slave_we_i,
	slave_addr_i,
	slave_be_i,
	slave_wdata_i,
	slave_rdata_o,
	master_req_o,
	master_add_o,
	master_we_o,
	master_wdata_o,
	master_be_o,
	master_gnt_i,
	master_r_valid_i,
	master_r_err_i,
	master_r_other_err_i,
	master_r_rdata_i,
	dmi_rst_ni,
	dmi_req_valid_i,
	dmi_req_ready_o,
	dmi_req_i,
	dmi_resp_valid_o,
	dmi_resp_ready_i,
	dmi_resp_o
);
	// Trace: design.sv:48141:13
	parameter [31:0] NrHarts = 1;
	// Trace: design.sv:48142:13
	parameter [31:0] BusWidth = 32;
	// Trace: design.sv:48143:13
	parameter [31:0] DmBaseAddress = 'h1000;
	// Trace: design.sv:48146:13
	parameter [NrHarts - 1:0] SelectableHarts = {NrHarts {1'b1}};
	// Trace: design.sv:48148:13
	parameter [0:0] ReadByteEnable = 1;
	// Trace: design.sv:48150:3
	input wire clk_i;
	// Trace: design.sv:48152:3
	input wire rst_ni;
	// Trace: design.sv:48153:3
	input wire testmode_i;
	// Trace: design.sv:48154:3
	output wire ndmreset_o;
	// Trace: design.sv:48155:3
	output wire dmactive_o;
	// Trace: design.sv:48156:3
	output wire [NrHarts - 1:0] debug_req_o;
	// Trace: design.sv:48158:3
	input wire [NrHarts - 1:0] unavailable_i;
	// Trace: design.sv:48159:3
	// removed localparam type dm_hartinfo_t
	input wire [(NrHarts * 32) - 1:0] hartinfo_i;
	// Trace: design.sv:48161:3
	input wire slave_req_i;
	// Trace: design.sv:48162:3
	input wire slave_we_i;
	// Trace: design.sv:48163:3
	input wire [BusWidth - 1:0] slave_addr_i;
	// Trace: design.sv:48164:3
	input wire [(BusWidth / 8) - 1:0] slave_be_i;
	// Trace: design.sv:48165:3
	input wire [BusWidth - 1:0] slave_wdata_i;
	// Trace: design.sv:48166:3
	output wire [BusWidth - 1:0] slave_rdata_o;
	// Trace: design.sv:48168:3
	output wire master_req_o;
	// Trace: design.sv:48169:3
	output wire [BusWidth - 1:0] master_add_o;
	// Trace: design.sv:48170:3
	output wire master_we_o;
	// Trace: design.sv:48171:3
	output wire [BusWidth - 1:0] master_wdata_o;
	// Trace: design.sv:48172:3
	output wire [(BusWidth / 8) - 1:0] master_be_o;
	// Trace: design.sv:48173:3
	input wire master_gnt_i;
	// Trace: design.sv:48174:3
	input wire master_r_valid_i;
	// Trace: design.sv:48175:3
	input wire master_r_err_i;
	// Trace: design.sv:48176:3
	input wire master_r_other_err_i;
	// Trace: design.sv:48177:3
	input wire [BusWidth - 1:0] master_r_rdata_i;
	// Trace: design.sv:48180:3
	input wire dmi_rst_ni;
	// Trace: design.sv:48183:3
	input wire dmi_req_valid_i;
	// Trace: design.sv:48184:3
	output wire dmi_req_ready_o;
	// Trace: design.sv:48185:3
	// removed localparam type dm_dtm_op_e
	// removed localparam type dm_dmi_req_t
	input wire [40:0] dmi_req_i;
	// Trace: design.sv:48187:3
	output wire dmi_resp_valid_o;
	// Trace: design.sv:48188:3
	input wire dmi_resp_ready_i;
	// Trace: design.sv:48189:3
	// removed localparam type dm_dmi_resp_t
	output wire [33:0] dmi_resp_o;
	// Trace: design.sv:48193:3
	wire [NrHarts - 1:0] halted;
	// Trace: design.sv:48195:3
	wire [NrHarts - 1:0] resumeack;
	// Trace: design.sv:48196:3
	wire [NrHarts - 1:0] haltreq;
	// Trace: design.sv:48197:3
	wire [NrHarts - 1:0] resumereq;
	// Trace: design.sv:48198:3
	wire clear_resumeack;
	// Trace: design.sv:48199:3
	wire cmd_valid;
	// Trace: design.sv:48200:3
	// removed localparam type dm_cmd_e
	// removed localparam type dm_command_t
	wire [31:0] cmd;
	// Trace: design.sv:48202:3
	wire cmderror_valid;
	// Trace: design.sv:48203:3
	// removed localparam type dm_cmderr_e
	wire [2:0] cmderror;
	// Trace: design.sv:48204:3
	wire cmdbusy;
	// Trace: design.sv:48205:3
	localparam [4:0] dm_ProgBufSize = 5'h08;
	wire [255:0] progbuf;
	// Trace: design.sv:48206:3
	localparam [3:0] dm_DataCount = 4'h2;
	wire [63:0] data_csrs_mem;
	// Trace: design.sv:48207:3
	wire [63:0] data_mem_csrs;
	// Trace: design.sv:48208:3
	wire data_valid;
	// Trace: design.sv:48209:3
	wire [19:0] hartsel;
	// Trace: design.sv:48211:3
	wire [BusWidth - 1:0] sbaddress_csrs_sba;
	// Trace: design.sv:48212:3
	wire [BusWidth - 1:0] sbaddress_sba_csrs;
	// Trace: design.sv:48213:3
	wire sbaddress_write_valid;
	// Trace: design.sv:48214:3
	wire sbreadonaddr;
	// Trace: design.sv:48215:3
	wire sbautoincrement;
	// Trace: design.sv:48216:3
	wire [2:0] sbaccess;
	// Trace: design.sv:48217:3
	wire sbreadondata;
	// Trace: design.sv:48218:3
	wire [BusWidth - 1:0] sbdata_write;
	// Trace: design.sv:48219:3
	wire sbdata_read_valid;
	// Trace: design.sv:48220:3
	wire sbdata_write_valid;
	// Trace: design.sv:48221:3
	wire [BusWidth - 1:0] sbdata_read;
	// Trace: design.sv:48222:3
	wire sbdata_valid;
	// Trace: design.sv:48223:3
	wire sbbusy;
	// Trace: design.sv:48224:3
	wire sberror_valid;
	// Trace: design.sv:48225:3
	wire [2:0] sberror;
	// Trace: design.sv:48228:3
	dm_csrs #(
		.NrHarts(NrHarts),
		.BusWidth(BusWidth),
		.SelectableHarts(SelectableHarts)
	) i_dm_csrs(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.testmode_i(testmode_i),
		.dmi_rst_ni(dmi_rst_ni),
		.dmi_req_valid_i(dmi_req_valid_i),
		.dmi_req_ready_o(dmi_req_ready_o),
		.dmi_req_i(dmi_req_i),
		.dmi_resp_valid_o(dmi_resp_valid_o),
		.dmi_resp_ready_i(dmi_resp_ready_i),
		.dmi_resp_o(dmi_resp_o),
		.ndmreset_o(ndmreset_o),
		.dmactive_o(dmactive_o),
		.hartsel_o(hartsel),
		.hartinfo_i(hartinfo_i),
		.halted_i(halted),
		.unavailable_i(unavailable_i),
		.resumeack_i(resumeack),
		.haltreq_o(haltreq),
		.resumereq_o(resumereq),
		.clear_resumeack_o(clear_resumeack),
		.cmd_valid_o(cmd_valid),
		.cmd_o(cmd),
		.cmderror_valid_i(cmderror_valid),
		.cmderror_i(cmderror),
		.cmdbusy_i(cmdbusy),
		.progbuf_o(progbuf),
		.data_i(data_mem_csrs),
		.data_valid_i(data_valid),
		.data_o(data_csrs_mem),
		.sbaddress_o(sbaddress_csrs_sba),
		.sbaddress_i(sbaddress_sba_csrs),
		.sbaddress_write_valid_o(sbaddress_write_valid),
		.sbreadonaddr_o(sbreadonaddr),
		.sbautoincrement_o(sbautoincrement),
		.sbaccess_o(sbaccess),
		.sbreadondata_o(sbreadondata),
		.sbdata_o(sbdata_write),
		.sbdata_read_valid_o(sbdata_read_valid),
		.sbdata_write_valid_o(sbdata_write_valid),
		.sbdata_i(sbdata_read),
		.sbdata_valid_i(sbdata_valid),
		.sbbusy_i(sbbusy),
		.sberror_valid_i(sberror_valid),
		.sberror_i(sberror)
	);
	// Trace: design.sv:48279:3
	dm_sba #(
		.BusWidth(BusWidth),
		.ReadByteEnable(ReadByteEnable)
	) i_dm_sba(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.dmactive_i(dmactive_o),
		.master_req_o(master_req_o),
		.master_add_o(master_add_o),
		.master_we_o(master_we_o),
		.master_wdata_o(master_wdata_o),
		.master_be_o(master_be_o),
		.master_gnt_i(master_gnt_i),
		.master_r_valid_i(master_r_valid_i),
		.master_r_err_i(master_r_err_i),
		.master_r_other_err_i(master_r_other_err_i),
		.master_r_rdata_i(master_r_rdata_i),
		.sbaddress_i(sbaddress_csrs_sba),
		.sbaddress_o(sbaddress_sba_csrs),
		.sbaddress_write_valid_i(sbaddress_write_valid),
		.sbreadonaddr_i(sbreadonaddr),
		.sbautoincrement_i(sbautoincrement),
		.sbaccess_i(sbaccess),
		.sbreadondata_i(sbreadondata),
		.sbdata_i(sbdata_write),
		.sbdata_read_valid_i(sbdata_read_valid),
		.sbdata_write_valid_i(sbdata_write_valid),
		.sbdata_o(sbdata_read),
		.sbdata_valid_o(sbdata_valid),
		.sbbusy_o(sbbusy),
		.sberror_valid_o(sberror_valid),
		.sberror_o(sberror)
	);
	// Trace: design.sv:48315:3
	dm_mem #(
		.NrHarts(NrHarts),
		.BusWidth(BusWidth),
		.SelectableHarts(SelectableHarts),
		.DmBaseAddress(DmBaseAddress)
	) i_dm_mem(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.debug_req_o(debug_req_o),
		.hartsel_i(hartsel),
		.haltreq_i(haltreq),
		.resumereq_i(resumereq),
		.clear_resumeack_i(clear_resumeack),
		.halted_o(halted),
		.resuming_o(resumeack),
		.cmd_valid_i(cmd_valid),
		.cmd_i(cmd),
		.cmderror_valid_o(cmderror_valid),
		.cmderror_o(cmderror),
		.cmdbusy_o(cmdbusy),
		.progbuf_i(progbuf),
		.data_i(data_csrs_mem),
		.data_o(data_mem_csrs),
		.data_valid_o(data_valid),
		.req_i(slave_req_i),
		.we_i(slave_we_i),
		.addr_i(slave_addr_i),
		.wdata_i(slave_wdata_i),
		.be_i(slave_be_i),
		.rdata_o(slave_rdata_o)
	);
endmodule
module dmi_jtag_tap (
	tck_i,
	tms_i,
	trst_ni,
	td_i,
	td_o,
	tdo_oe_o,
	testmode_i,
	tck_o,
	dmi_clear_o,
	update_o,
	capture_o,
	shift_o,
	tdi_o,
	dtmcs_select_o,
	dtmcs_tdo_i,
	dmi_select_o,
	dmi_tdo_i
);
	reg _sv2v_0;
	// Trace: design.sv:48367:13
	parameter [31:0] IrLength = 5;
	// Trace: design.sv:48369:13
	parameter [31:0] IdcodeValue = 32'h00000001;
	// Trace: design.sv:48375:3
	input wire tck_i;
	// Trace: design.sv:48376:3
	input wire tms_i;
	// Trace: design.sv:48377:3
	input wire trst_ni;
	// Trace: design.sv:48378:3
	input wire td_i;
	// Trace: design.sv:48379:3
	output reg td_o;
	// Trace: design.sv:48380:3
	output reg tdo_oe_o;
	// Trace: design.sv:48381:3
	input wire testmode_i;
	// Trace: design.sv:48383:3
	output wire tck_o;
	// Trace: design.sv:48385:3
	output wire dmi_clear_o;
	// Trace: design.sv:48386:3
	output wire update_o;
	// Trace: design.sv:48387:3
	output wire capture_o;
	// Trace: design.sv:48388:3
	output wire shift_o;
	// Trace: design.sv:48389:3
	output wire tdi_o;
	// Trace: design.sv:48390:3
	output reg dtmcs_select_o;
	// Trace: design.sv:48391:3
	input wire dtmcs_tdo_i;
	// Trace: design.sv:48393:3
	output reg dmi_select_o;
	// Trace: design.sv:48394:3
	input wire dmi_tdo_i;
	// Trace: design.sv:48397:3
	// removed localparam type tap_state_e
	// Trace: design.sv:48404:3
	reg [3:0] tap_state_q;
	reg [3:0] tap_state_d;
	// Trace: design.sv:48405:3
	reg update_dr;
	reg shift_dr;
	reg capture_dr;
	// Trace: design.sv:48407:3
	// removed localparam type ir_reg_e
	// Trace: design.sv:48420:3
	reg [IrLength - 1:0] jtag_ir_shift_d;
	reg [IrLength - 1:0] jtag_ir_shift_q;
	// Trace: design.sv:48422:3
	reg [IrLength - 1:0] jtag_ir_d;
	reg [IrLength - 1:0] jtag_ir_q;
	// Trace: design.sv:48423:3
	reg capture_ir;
	reg shift_ir;
	reg update_ir;
	reg test_logic_reset;
	// Trace: design.sv:48425:3
	function automatic [IrLength - 1:0] sv2v_cast_154DA;
		input reg [IrLength - 1:0] inp;
		sv2v_cast_154DA = inp;
	endfunction
	always @(*) begin : p_jtag
		if (_sv2v_0)
			;
		// Trace: design.sv:48426:5
		jtag_ir_shift_d = jtag_ir_shift_q;
		// Trace: design.sv:48427:5
		jtag_ir_d = jtag_ir_q;
		// Trace: design.sv:48430:5
		if (shift_ir)
			// Trace: design.sv:48431:7
			jtag_ir_shift_d = {td_i, jtag_ir_shift_q[IrLength - 1:1]};
		if (capture_ir)
			// Trace: design.sv:48436:7
			jtag_ir_shift_d = sv2v_cast_154DA(4'b0101);
		if (update_ir)
			// Trace: design.sv:48441:7
			jtag_ir_d = sv2v_cast_154DA(jtag_ir_shift_q);
		if (test_logic_reset)
			// Trace: design.sv:48446:7
			jtag_ir_d = sv2v_cast_154DA('h1);
	end
	// Trace: design.sv:48450:3
	always @(posedge tck_i or negedge trst_ni) begin : p_jtag_ir_reg
		// Trace: design.sv:48451:5
		if (!trst_ni) begin
			// Trace: design.sv:48452:7
			jtag_ir_shift_q <= 1'sb0;
			// Trace: design.sv:48453:7
			jtag_ir_q <= sv2v_cast_154DA('h1);
		end
		else begin
			// Trace: design.sv:48455:7
			jtag_ir_shift_q <= jtag_ir_shift_d;
			// Trace: design.sv:48456:7
			jtag_ir_q <= jtag_ir_d;
		end
	end
	// Trace: design.sv:48466:3
	reg [31:0] idcode_d;
	reg [31:0] idcode_q;
	// Trace: design.sv:48467:3
	reg idcode_select;
	// Trace: design.sv:48468:3
	reg bypass_select;
	// Trace: design.sv:48470:3
	reg bypass_d;
	reg bypass_q;
	// Trace: design.sv:48472:3
	function automatic [30:0] sv2v_cast_31;
		input reg [30:0] inp;
		sv2v_cast_31 = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:48473:5
		idcode_d = idcode_q;
		// Trace: design.sv:48474:5
		bypass_d = bypass_q;
		// Trace: design.sv:48476:5
		if (capture_dr) begin
			// Trace: design.sv:48477:7
			if (idcode_select)
				// Trace: design.sv:48477:26
				idcode_d = IdcodeValue;
			if (bypass_select)
				// Trace: design.sv:48478:26
				bypass_d = 1'b0;
		end
		if (shift_dr) begin
			// Trace: design.sv:48482:7
			if (idcode_select)
				// Trace: design.sv:48482:27
				idcode_d = {td_i, sv2v_cast_31(idcode_q >> 1)};
			if (bypass_select)
				// Trace: design.sv:48483:27
				bypass_d = td_i;
		end
	end
	// Trace: design.sv:48490:3
	always @(*) begin : p_data_reg_sel
		if (_sv2v_0)
			;
		// Trace: design.sv:48491:5
		dmi_select_o = 1'b0;
		// Trace: design.sv:48492:5
		dtmcs_select_o = 1'b0;
		// Trace: design.sv:48493:5
		idcode_select = 1'b0;
		// Trace: design.sv:48494:5
		bypass_select = 1'b0;
		// Trace: design.sv:48495:5
		(* full_case, parallel_case *)
		case (jtag_ir_q)
			sv2v_cast_154DA('h0):
				// Trace: design.sv:48496:18
				bypass_select = 1'b1;
			sv2v_cast_154DA('h1):
				// Trace: design.sv:48497:18
				idcode_select = 1'b1;
			sv2v_cast_154DA('h10):
				// Trace: design.sv:48498:18
				dtmcs_select_o = 1'b1;
			sv2v_cast_154DA('h11):
				// Trace: design.sv:48499:18
				dmi_select_o = 1'b1;
			sv2v_cast_154DA('h1f):
				// Trace: design.sv:48500:18
				bypass_select = 1'b1;
			default:
				// Trace: design.sv:48501:18
				bypass_select = 1'b1;
		endcase
	end
	// Trace: design.sv:48508:3
	reg tdo_mux;
	// Trace: design.sv:48510:3
	always @(*) begin : p_out_sel
		if (_sv2v_0)
			;
		// Trace: design.sv:48512:5
		if (shift_ir)
			// Trace: design.sv:48513:7
			tdo_mux = jtag_ir_shift_q[0];
		else
			// Trace: design.sv:48516:7
			(* full_case, parallel_case *)
			case (jtag_ir_q)
				sv2v_cast_154DA('h1):
					// Trace: design.sv:48517:25
					tdo_mux = idcode_q[0];
				sv2v_cast_154DA('h10):
					// Trace: design.sv:48518:25
					tdo_mux = dtmcs_tdo_i;
				sv2v_cast_154DA('h11):
					// Trace: design.sv:48519:25
					tdo_mux = dmi_tdo_i;
				default:
					// Trace: design.sv:48520:25
					tdo_mux = bypass_q;
			endcase
	end
	// Trace: design.sv:48528:3
	wire tck_n;
	wire tck_ni;
	// Trace: design.sv:48530:3
	cluster_clock_inverter i_tck_inv(
		.clk_i(tck_i),
		.clk_o(tck_ni)
	);
	// Trace: design.sv:48535:3
	pulp_clock_mux2 i_dft_tck_mux(
		.clk0_i(tck_ni),
		.clk1_i(tck_i),
		.clk_sel_i(testmode_i),
		.clk_o(tck_n)
	);
	// Trace: design.sv:48543:3
	always @(posedge tck_n or negedge trst_ni) begin : p_tdo_regs
		// Trace: design.sv:48544:5
		if (!trst_ni) begin
			// Trace: design.sv:48545:7
			td_o <= 1'b0;
			// Trace: design.sv:48546:7
			tdo_oe_o <= 1'b0;
		end
		else begin
			// Trace: design.sv:48548:7
			td_o <= tdo_mux;
			// Trace: design.sv:48549:7
			tdo_oe_o <= shift_ir | shift_dr;
		end
	end
	// Trace: design.sv:48556:3
	always @(*) begin : p_tap_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:48558:5
		test_logic_reset = 1'b0;
		// Trace: design.sv:48560:5
		capture_dr = 1'b0;
		// Trace: design.sv:48561:5
		shift_dr = 1'b0;
		// Trace: design.sv:48562:5
		update_dr = 1'b0;
		// Trace: design.sv:48564:5
		capture_ir = 1'b0;
		// Trace: design.sv:48565:5
		shift_ir = 1'b0;
		// Trace: design.sv:48567:5
		update_ir = 1'b0;
		// Trace: design.sv:48569:5
		(* full_case, parallel_case *)
		case (tap_state_q)
			4'd0: begin
				// Trace: design.sv:48571:9
				tap_state_d = (tms_i ? 4'd0 : 4'd1);
				// Trace: design.sv:48572:9
				test_logic_reset = 1'b1;
			end
			4'd1:
				// Trace: design.sv:48575:9
				tap_state_d = (tms_i ? 4'd2 : 4'd1);
			4'd2:
				// Trace: design.sv:48579:9
				tap_state_d = (tms_i ? 4'd9 : 4'd3);
			4'd3: begin
				// Trace: design.sv:48582:9
				capture_dr = 1'b1;
				// Trace: design.sv:48583:9
				tap_state_d = (tms_i ? 4'd5 : 4'd4);
			end
			4'd4: begin
				// Trace: design.sv:48586:9
				shift_dr = 1'b1;
				// Trace: design.sv:48587:9
				tap_state_d = (tms_i ? 4'd5 : 4'd4);
			end
			4'd5:
				// Trace: design.sv:48590:9
				tap_state_d = (tms_i ? 4'd8 : 4'd6);
			4'd6:
				// Trace: design.sv:48593:9
				tap_state_d = (tms_i ? 4'd7 : 4'd6);
			4'd7:
				// Trace: design.sv:48596:9
				tap_state_d = (tms_i ? 4'd8 : 4'd4);
			4'd8: begin
				// Trace: design.sv:48599:9
				update_dr = 1'b1;
				// Trace: design.sv:48600:9
				tap_state_d = (tms_i ? 4'd2 : 4'd1);
			end
			4'd9:
				// Trace: design.sv:48604:9
				tap_state_d = (tms_i ? 4'd0 : 4'd10);
			4'd10: begin
				// Trace: design.sv:48611:9
				capture_ir = 1'b1;
				// Trace: design.sv:48612:9
				tap_state_d = (tms_i ? 4'd12 : 4'd11);
			end
			4'd11: begin
				// Trace: design.sv:48619:9
				shift_ir = 1'b1;
				// Trace: design.sv:48620:9
				tap_state_d = (tms_i ? 4'd12 : 4'd11);
			end
			4'd12:
				// Trace: design.sv:48623:9
				tap_state_d = (tms_i ? 4'd15 : 4'd13);
			4'd13:
				// Trace: design.sv:48627:9
				tap_state_d = (tms_i ? 4'd14 : 4'd13);
			4'd14:
				// Trace: design.sv:48630:9
				tap_state_d = (tms_i ? 4'd15 : 4'd11);
			4'd15: begin
				// Trace: design.sv:48637:9
				update_ir = 1'b1;
				// Trace: design.sv:48638:9
				tap_state_d = (tms_i ? 4'd2 : 4'd1);
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:48644:3
	always @(posedge tck_i or negedge trst_ni) begin : p_regs
		// Trace: design.sv:48645:5
		if (!trst_ni) begin
			// Trace: design.sv:48646:7
			tap_state_q <= 4'd1;
			// Trace: design.sv:48647:7
			idcode_q <= IdcodeValue;
			// Trace: design.sv:48648:7
			bypass_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:48650:7
			tap_state_q <= tap_state_d;
			// Trace: design.sv:48651:7
			idcode_q <= idcode_d;
			// Trace: design.sv:48652:7
			bypass_q <= bypass_d;
		end
	end
	// Trace: design.sv:48658:3
	assign tck_o = tck_i;
	// Trace: design.sv:48659:3
	assign tdi_o = td_i;
	// Trace: design.sv:48660:3
	assign update_o = update_dr;
	// Trace: design.sv:48661:3
	assign shift_o = shift_dr;
	// Trace: design.sv:48662:3
	assign capture_o = capture_dr;
	// Trace: design.sv:48663:3
	assign dmi_clear_o = test_logic_reset;
	initial _sv2v_0 = 0;
endmodule
// removed package "fpnew_pkg"
module fpnew_cast_multi_2E827_EA7A2 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	reg _sv2v_0;
	// Trace: design.sv:49179:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: design.sv:49180:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtConfig = 1'sb1;
	// Trace: design.sv:49182:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: design.sv:49183:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: design.sv:49184:38
	// removed localparam type TagType
	// Trace: design.sv:49185:38
	// removed localparam type AuxType
	// Trace: design.sv:49187:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:34
		input reg signed [31:0] a;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:41
		input reg signed [31:0] b;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:296:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:308:48
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:309:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:5
			begin : sv2v_autoblock_1
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:312:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	function automatic [1:0] sv2v_cast_CDB06;
		input reg [1:0] inp;
		sv2v_cast_CDB06 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:88:45
		input reg [1:0] ifmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:89:5
		(* full_case, parallel_case *)
		case (ifmt)
			sv2v_cast_CDB06(0): fpnew_pkg_int_width = 8;
			sv2v_cast_CDB06(1): fpnew_pkg_int_width = 16;
			sv2v_cast_CDB06(2): fpnew_pkg_int_width = 32;
			sv2v_cast_CDB06(3): fpnew_pkg_int_width = 64;
			default: begin
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:96:9
				$fatal(1, "Invalid INT format supplied");
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:100:9
				fpnew_pkg_int_width = sv2v_cast_CDB06(0);
			end
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:355:49
		input reg [0:3] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:356:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:357:5
			begin : sv2v_autoblock_2
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:357:10
				reg signed [31:0] ifmt;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:357:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:358:7
						if (cfg[ifmt])
							// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:358:22
							res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_CDB06(ifmt)));
					end
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_maximum(fpnew_pkg_max_fp_width(FpFmtConfig), fpnew_pkg_max_int_width(IntFmtConfig));
	// Trace: design.sv:49189:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: design.sv:49191:3
	input wire clk_i;
	// Trace: design.sv:49192:3
	input wire rst_ni;
	// Trace: design.sv:49194:3
	input wire [WIDTH - 1:0] operands_i;
	// Trace: design.sv:49195:3
	input wire [4:0] is_boxed_i;
	// Trace: design.sv:49196:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:49197:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:49198:3
	input wire op_mod_i;
	// Trace: design.sv:49199:3
	input wire [2:0] src_fmt_i;
	// Trace: design.sv:49200:3
	input wire [2:0] dst_fmt_i;
	// Trace: design.sv:49201:3
	input wire [1:0] int_fmt_i;
	// Trace: design.sv:49202:3
	input wire tag_i;
	// Trace: design.sv:49203:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: design.sv:49205:3
	input wire in_valid_i;
	// Trace: design.sv:49206:3
	output wire in_ready_o;
	// Trace: design.sv:49207:3
	input wire flush_i;
	// Trace: design.sv:49209:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: design.sv:49210:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: design.sv:49211:3
	output wire extension_bit_o;
	// Trace: design.sv:49212:3
	output wire tag_o;
	// Trace: design.sv:49213:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: design.sv:49215:3
	output wire out_valid_o;
	// Trace: design.sv:49216:3
	input wire out_ready_i;
	// Trace: design.sv:49218:3
	output wire busy_o;
	// Trace: design.sv:49224:3
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	// Trace: design.sv:49225:3
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	// Trace: design.sv:49227:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:326:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:327:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:331:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:332:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:340:49
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:341:5
		reg [63:0] res;
		begin
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:342:5
			res = 1'sb0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:343:5
			begin : sv2v_autoblock_3
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:343:10
				reg [31:0] fmt;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:343:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:345:9
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt))));
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:346:9
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_5D882(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	// Trace: design.sv:49229:3
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	// Trace: design.sv:49230:3
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	// Trace: design.sv:49231:3
	localparam [31:0] SUPER_BIAS = (2 ** (SUPER_EXP_BITS - 1)) - 1;
	// Trace: design.sv:49234:3
	localparam [31:0] INT_MAN_WIDTH = fpnew_pkg_maximum(SUPER_MAN_BITS + 1, MAX_INT_WIDTH);
	// Trace: design.sv:49236:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(INT_MAN_WIDTH);
	// Trace: design.sv:49239:3
	localparam [31:0] INT_EXP_WIDTH = fpnew_pkg_maximum($clog2(MAX_INT_WIDTH), fpnew_pkg_maximum(SUPER_EXP_BITS, $clog2(SUPER_BIAS + SUPER_MAN_BITS))) + 1;
	// Trace: design.sv:49242:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: design.sv:49247:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: design.sv:49252:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: design.sv:49262:3
	wire [WIDTH - 1:0] operands_q;
	// Trace: design.sv:49263:3
	wire [4:0] is_boxed_q;
	// Trace: design.sv:49264:3
	wire op_mod_q;
	// Trace: design.sv:49265:3
	wire [2:0] src_fmt_q;
	// Trace: design.sv:49266:3
	wire [2:0] dst_fmt_q;
	// Trace: design.sv:49267:3
	wire [1:0] int_fmt_q;
	// Trace: design.sv:49270:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * WIDTH) + ((NUM_INP_REGS * WIDTH) - 1) : ((NUM_INP_REGS + 1) * WIDTH) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * WIDTH : 0)] inp_pipe_operands_q;
	// Trace: design.sv:49271:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)] inp_pipe_is_boxed_q;
	// Trace: design.sv:49272:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: design.sv:49273:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: design.sv:49274:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: design.sv:49275:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	// Trace: design.sv:49276:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: design.sv:49277:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] inp_pipe_int_fmt_q;
	// Trace: design.sv:49278:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: design.sv:49279:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: design.sv:49280:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: design.sv:49282:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: design.sv:49285:3
	wire [WIDTH * 1:1] sv2v_tmp_933AE;
	assign sv2v_tmp_933AE = operands_i;
	always @(*) inp_pipe_operands_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * WIDTH+:WIDTH] = sv2v_tmp_933AE;
	// Trace: design.sv:49286:3
	wire [5:1] sv2v_tmp_7038A;
	assign sv2v_tmp_7038A = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS] = sv2v_tmp_7038A;
	// Trace: design.sv:49287:3
	wire [3:1] sv2v_tmp_AA272;
	assign sv2v_tmp_AA272 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_AA272;
	// Trace: design.sv:49288:3
	wire [4:1] sv2v_tmp_14A3A;
	assign sv2v_tmp_14A3A = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_14A3A;
	// Trace: design.sv:49289:3
	wire [1:1] sv2v_tmp_72E02;
	assign sv2v_tmp_72E02 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_72E02;
	// Trace: design.sv:49290:3
	wire [3:1] sv2v_tmp_8EF42;
	assign sv2v_tmp_8EF42 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_8EF42;
	// Trace: design.sv:49291:3
	wire [3:1] sv2v_tmp_B0F12;
	assign sv2v_tmp_B0F12 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_B0F12;
	// Trace: design.sv:49292:3
	wire [2:1] sv2v_tmp_C9BC4;
	assign sv2v_tmp_C9BC4 = int_fmt_i;
	always @(*) inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_C9BC4;
	// Trace: design.sv:49293:3
	wire [1:1] sv2v_tmp_DE624;
	assign sv2v_tmp_DE624 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_DE624;
	// Trace: design.sv:49294:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_7E5D6;
	assign sv2v_tmp_7E5D6 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_7E5D6;
	// Trace: design.sv:49295:3
	wire [1:1] sv2v_tmp_CFC25;
	assign sv2v_tmp_CFC25 = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_CFC25;
	// Trace: design.sv:49297:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: design.sv:49299:3
	genvar _gv_i_69;
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_533F1;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_533F1 = inp;
	endfunction
	generate
		for (_gv_i_69 = 0; _gv_i_69 < NUM_INP_REGS; _gv_i_69 = _gv_i_69 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_69;
			// Trace: design.sv:49301:5
			wire reg_ena;
			// Trace: design.sv:49305:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:49307:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:49307:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:49307:485
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:49307:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:49307:715
						inp_pipe_valid_q[i + 1] <= 1'b0;
					else if (inp_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:49307:867
						inp_pipe_valid_q[i + 1] <= inp_pipe_valid_q[i];
			// Trace: design.sv:49309:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:49311:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49311:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49311:265
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49311:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49311:552
						inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * WIDTH+:WIDTH];
			// Trace: macro expansion of FFL at design.sv:49312:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49312:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49312:265
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49312:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49312:552
						inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS+:NUM_FORMATS];
			// Trace: macro expansion of FFL at design.sv:49313:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49313:180
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49313:277
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at design.sv:49313:467
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49313:564
						inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:49314:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49314:182
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49314:279
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_4CD2E(0);
				else
					// Trace: macro expansion of FFL at design.sv:49314:469
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49314:566
						inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
			// Trace: macro expansion of FFL at design.sv:49315:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49315:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49315:265
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49315:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49315:552
						inp_pipe_op_mod_q[i + 1] <= inp_pipe_op_mod_q[i];
			// Trace: macro expansion of FFL at design.sv:49316:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49316:192
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49316:289
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_5D882(0);
				else
					// Trace: macro expansion of FFL at design.sv:49316:479
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49316:576
						inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:49317:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49317:192
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49317:289
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_5D882(0);
				else
					// Trace: macro expansion of FFL at design.sv:49317:479
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49317:576
						inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:49318:96
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49318:193
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49318:290
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_CDB06(0);
				else
					// Trace: macro expansion of FFL at design.sv:49318:480
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49318:577
						inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:49319:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49319:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49319:275
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:49319:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49319:562
						inp_pipe_tag_q[i + 1] <= inp_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:49320:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49320:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49320:275
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_533F1(1'sb0);
				else
					// Trace: macro expansion of FFL at design.sv:49320:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49320:562
						inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
		end
	endgenerate
	// Trace: design.sv:49323:3
	assign operands_q = inp_pipe_operands_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * WIDTH+:WIDTH];
	// Trace: design.sv:49324:3
	assign is_boxed_q = inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS];
	// Trace: design.sv:49325:3
	assign op_mod_q = inp_pipe_op_mod_q[NUM_INP_REGS];
	// Trace: design.sv:49326:3
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: design.sv:49327:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: design.sv:49328:3
	assign int_fmt_q = inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	// Trace: design.sv:49333:3
	wire src_is_int;
	wire dst_is_int;
	// Trace: design.sv:49335:3
	assign src_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_4CD2E(12);
	// Trace: design.sv:49336:3
	assign dst_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_4CD2E(11);
	// Trace: design.sv:49338:3
	wire [INT_MAN_WIDTH - 1:0] encoded_mant;
	// Trace: design.sv:49340:3
	wire [4:0] fmt_sign;
	// Trace: design.sv:49341:3
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_exponent;
	// Trace: design.sv:49342:3
	wire [(NUM_FORMATS * INT_MAN_WIDTH) - 1:0] fmt_mantissa;
	// Trace: design.sv:49343:3
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_shift_compensation;
	// Trace: design.sv:49345:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [39:0] info;
	// Trace: design.sv:49347:3
	reg [(NUM_INT_FORMATS * INT_MAN_WIDTH) - 1:0] ifmt_input_val;
	// Trace: design.sv:49348:3
	wire int_sign;
	// Trace: design.sv:49349:3
	wire [INT_MAN_WIDTH - 1:0] int_value;
	wire [INT_MAN_WIDTH - 1:0] int_mantissa;
	// Trace: design.sv:49352:3
	genvar _gv_fmt_1;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [0:0] sv2v_cast_1_signed;
		input reg signed [0:0] inp;
		sv2v_cast_1_signed = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_fmt_1 = 0; _gv_fmt_1 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_1 = _gv_fmt_1 + 1) begin : fmt_init_inputs
			localparam fmt = _gv_fmt_1;
			// Trace: design.sv:49354:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			// Trace: design.sv:49355:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:49356:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_5D882(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: design.sv:49360:7
				fpnew_classifier #(
					.FpFormat(sv2v_cast_5D882(fmt)),
					.NumOperands(1)
				) i_fpnew_classifier(
					.operands_i(operands_q[FP_WIDTH - 1:0]),
					.is_boxed_i(is_boxed_q[fmt]),
					.info_o(info[fmt * 8+:8])
				);
				// Trace: design.sv:49369:7
				assign fmt_sign[fmt] = operands_q[FP_WIDTH - 1];
				// Trace: design.sv:49370:7
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed({1'b0, operands_q[MAN_BITS+:EXP_BITS]});
				// Trace: design.sv:49371:7
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {info[(fmt * 8) + 7], operands_q[MAN_BITS - 1:0]};
				// Trace: design.sv:49373:7
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed((INT_MAN_WIDTH - 1) - MAN_BITS);
			end
			else begin : inactive_format
				// Trace: design.sv:49375:7
				assign info[fmt * 8+:8] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: design.sv:49376:7
				assign fmt_sign[fmt] = fpnew_pkg_DONT_CARE;
				// Trace: design.sv:49377:7
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
				// Trace: design.sv:49378:7
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				// Trace: design.sv:49379:7
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	// Trace: design.sv:49384:3
	genvar _gv_ifmt_1;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	generate
		for (_gv_ifmt_1 = 0; _gv_ifmt_1 < sv2v_cast_32_signed(NUM_INT_FORMATS); _gv_ifmt_1 = _gv_ifmt_1 + 1) begin : gen_sign_extend_int
			localparam ifmt = _gv_ifmt_1;
			// Trace: design.sv:49386:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_CDB06(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: design.sv:49389:7
				always @(*) begin : sign_ext_input
					if (_sv2v_0)
						;
					// Trace: design.sv:49391:9
					ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {sv2v_cast_1(operands_q[INT_WIDTH - 1] & ~op_mod_q)}};
					// Trace: design.sv:49392:9
					ifmt_input_val[(ifmt * INT_MAN_WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = operands_q[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				// Trace: design.sv:49395:7
				wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_F208D;
				assign sv2v_tmp_F208D = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_F208D;
			end
		end
	endgenerate
	// Trace: design.sv:49400:3
	assign int_value = ifmt_input_val[int_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	// Trace: design.sv:49401:3
	assign int_sign = int_value[INT_MAN_WIDTH - 1] & ~op_mod_q;
	// Trace: design.sv:49402:3
	assign int_mantissa = (int_sign ? $unsigned(-int_value) : int_value);
	// Trace: design.sv:49405:3
	assign encoded_mant = (src_is_int ? int_mantissa : fmt_mantissa[src_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
	// Trace: design.sv:49410:3
	wire signed [INT_EXP_WIDTH - 1:0] src_bias;
	// Trace: design.sv:49411:3
	wire signed [INT_EXP_WIDTH - 1:0] src_exp;
	// Trace: design.sv:49412:3
	wire signed [INT_EXP_WIDTH - 1:0] src_subnormal;
	// Trace: design.sv:49413:3
	wire signed [INT_EXP_WIDTH - 1:0] src_offset;
	// Trace: design.sv:49415:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:336:40
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:337:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	assign src_bias = $signed(fpnew_pkg_bias(src_fmt_q));
	// Trace: design.sv:49416:3
	assign src_exp = fmt_exponent[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: design.sv:49417:3
	assign src_subnormal = $signed({1'b0, info[(src_fmt_q * 8) + 6]});
	// Trace: design.sv:49418:3
	assign src_offset = fmt_shift_compensation[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: design.sv:49420:3
	wire input_sign;
	// Trace: design.sv:49421:3
	wire signed [INT_EXP_WIDTH - 1:0] input_exp;
	// Trace: design.sv:49422:3
	wire [INT_MAN_WIDTH - 1:0] input_mant;
	// Trace: design.sv:49423:3
	wire mant_is_zero;
	// Trace: design.sv:49425:3
	wire signed [INT_EXP_WIDTH - 1:0] fp_input_exp;
	// Trace: design.sv:49426:3
	wire signed [INT_EXP_WIDTH - 1:0] int_input_exp;
	// Trace: design.sv:49429:3
	wire [LZC_RESULT_WIDTH - 1:0] renorm_shamt;
	// Trace: design.sv:49430:3
	wire [LZC_RESULT_WIDTH:0] renorm_shamt_sgn;
	// Trace: design.sv:49433:3
	lzc #(
		.WIDTH(INT_MAN_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(encoded_mant),
		.cnt_o(renorm_shamt),
		.empty_o(mant_is_zero)
	);
	// Trace: design.sv:49441:3
	assign renorm_shamt_sgn = $signed({1'b0, renorm_shamt});
	// Trace: design.sv:49444:3
	assign input_sign = (src_is_int ? int_sign : fmt_sign[src_fmt_q]);
	// Trace: design.sv:49446:3
	assign input_mant = encoded_mant << renorm_shamt;
	// Trace: design.sv:49448:3
	assign fp_input_exp = $signed((((src_exp + src_subnormal) - src_bias) - renorm_shamt_sgn) + src_offset);
	// Trace: design.sv:49450:3
	assign int_input_exp = $signed((INT_MAN_WIDTH - 1) - renorm_shamt_sgn);
	// Trace: design.sv:49452:3
	assign input_exp = (src_is_int ? int_input_exp : fp_input_exp);
	// Trace: design.sv:49454:3
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp;
	// Trace: design.sv:49457:3
	assign destination_exp = input_exp + $signed(fpnew_pkg_bias(dst_fmt_q));
	// Trace: design.sv:49463:3
	wire input_sign_q;
	// Trace: design.sv:49464:3
	wire signed [INT_EXP_WIDTH - 1:0] input_exp_q;
	// Trace: design.sv:49465:3
	wire [INT_MAN_WIDTH - 1:0] input_mant_q;
	// Trace: design.sv:49466:3
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp_q;
	// Trace: design.sv:49467:3
	wire src_is_int_q;
	// Trace: design.sv:49468:3
	wire dst_is_int_q;
	// Trace: design.sv:49469:3
	wire [7:0] info_q;
	// Trace: design.sv:49470:3
	wire mant_is_zero_q;
	// Trace: design.sv:49471:3
	wire op_mod_q2;
	// Trace: design.sv:49472:3
	wire [2:0] rnd_mode_q;
	// Trace: design.sv:49473:3
	wire [2:0] src_fmt_q2;
	// Trace: design.sv:49474:3
	wire [2:0] dst_fmt_q2;
	// Trace: design.sv:49475:3
	wire [1:0] int_fmt_q2;
	// Trace: design.sv:49479:3
	reg [0:NUM_MID_REGS] mid_pipe_input_sign_q;
	// Trace: design.sv:49480:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_input_exp_q;
	// Trace: design.sv:49481:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_MAN_WIDTH) + ((NUM_MID_REGS * INT_MAN_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_MAN_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_MAN_WIDTH : 0)] mid_pipe_input_mant_q;
	// Trace: design.sv:49482:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_dest_exp_q;
	// Trace: design.sv:49483:3
	reg [0:NUM_MID_REGS] mid_pipe_src_is_int_q;
	// Trace: design.sv:49484:3
	reg [0:NUM_MID_REGS] mid_pipe_dst_is_int_q;
	// Trace: design.sv:49485:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 8) + ((NUM_MID_REGS * 8) - 1) : ((NUM_MID_REGS + 1) * 8) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 8 : 0)] mid_pipe_info_q;
	// Trace: design.sv:49486:3
	reg [0:NUM_MID_REGS] mid_pipe_mant_zero_q;
	// Trace: design.sv:49487:3
	reg [0:NUM_MID_REGS] mid_pipe_op_mod_q;
	// Trace: design.sv:49488:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: design.sv:49489:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_src_fmt_q;
	// Trace: design.sv:49490:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	// Trace: design.sv:49491:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] mid_pipe_int_fmt_q;
	// Trace: design.sv:49492:3
	reg [0:NUM_MID_REGS] mid_pipe_tag_q;
	// Trace: design.sv:49493:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	// Trace: design.sv:49494:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: design.sv:49496:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: design.sv:49499:3
	wire [1:1] sv2v_tmp_73C39;
	assign sv2v_tmp_73C39 = input_sign;
	always @(*) mid_pipe_input_sign_q[0] = sv2v_tmp_73C39;
	// Trace: design.sv:49500:3
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_D63AF;
	assign sv2v_tmp_D63AF = input_exp;
	always @(*) mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_D63AF;
	// Trace: design.sv:49501:3
	wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_CED01;
	assign sv2v_tmp_CED01 = input_mant;
	always @(*) mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_CED01;
	// Trace: design.sv:49502:3
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_5026E;
	assign sv2v_tmp_5026E = destination_exp;
	always @(*) mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_5026E;
	// Trace: design.sv:49503:3
	wire [1:1] sv2v_tmp_6F1F9;
	assign sv2v_tmp_6F1F9 = src_is_int;
	always @(*) mid_pipe_src_is_int_q[0] = sv2v_tmp_6F1F9;
	// Trace: design.sv:49504:3
	wire [1:1] sv2v_tmp_202B9;
	assign sv2v_tmp_202B9 = dst_is_int;
	always @(*) mid_pipe_dst_is_int_q[0] = sv2v_tmp_202B9;
	// Trace: design.sv:49505:3
	wire [8:1] sv2v_tmp_C577A;
	assign sv2v_tmp_C577A = info[src_fmt_q * 8+:8];
	always @(*) mid_pipe_info_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 8+:8] = sv2v_tmp_C577A;
	// Trace: design.sv:49506:3
	wire [1:1] sv2v_tmp_CCDAF;
	assign sv2v_tmp_CCDAF = mant_is_zero;
	always @(*) mid_pipe_mant_zero_q[0] = sv2v_tmp_CCDAF;
	// Trace: design.sv:49507:3
	wire [1:1] sv2v_tmp_0DC3D;
	assign sv2v_tmp_0DC3D = op_mod_q;
	always @(*) mid_pipe_op_mod_q[0] = sv2v_tmp_0DC3D;
	// Trace: design.sv:49508:3
	wire [3:1] sv2v_tmp_EC44B;
	assign sv2v_tmp_EC44B = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_EC44B;
	// Trace: design.sv:49509:3
	wire [3:1] sv2v_tmp_8D32D;
	assign sv2v_tmp_8D32D = src_fmt_q;
	always @(*) mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_8D32D;
	// Trace: design.sv:49510:3
	wire [3:1] sv2v_tmp_9DD7D;
	assign sv2v_tmp_9DD7D = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_9DD7D;
	// Trace: design.sv:49511:3
	wire [2:1] sv2v_tmp_5CA4B;
	assign sv2v_tmp_5CA4B = int_fmt_q;
	always @(*) mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_5CA4B;
	// Trace: design.sv:49512:3
	wire [1:1] sv2v_tmp_7259D;
	assign sv2v_tmp_7259D = inp_pipe_tag_q[NUM_INP_REGS];
	always @(*) mid_pipe_tag_q[0] = sv2v_tmp_7259D;
	// Trace: design.sv:49513:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_88919;
	assign sv2v_tmp_88919 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_88919;
	// Trace: design.sv:49514:3
	wire [1:1] sv2v_tmp_C7159;
	assign sv2v_tmp_C7159 = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_C7159;
	// Trace: design.sv:49516:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: design.sv:49519:3
	genvar _gv_i_70;
	generate
		for (_gv_i_70 = 0; _gv_i_70 < NUM_MID_REGS; _gv_i_70 = _gv_i_70 + 1) begin : gen_inside_pipeline
			localparam i = _gv_i_70;
			// Trace: design.sv:49521:5
			wire reg_ena;
			// Trace: design.sv:49525:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:49527:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:49527:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:49527:485
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:49527:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:49527:715
						mid_pipe_valid_q[i + 1] <= 1'b0;
					else if (mid_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:49527:867
						mid_pipe_valid_q[i + 1] <= mid_pipe_valid_q[i];
			// Trace: design.sv:49529:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:49531:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49531:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49531:269
					mid_pipe_input_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49531:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49531:556
						mid_pipe_input_sign_q[i + 1] <= mid_pipe_input_sign_q[i];
			// Trace: macro expansion of FFL at design.sv:49532:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49532:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49532:269
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49532:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49532:556
						mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
			// Trace: macro expansion of FFL at design.sv:49533:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49533:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49533:269
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49533:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49533:556
						mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_MAN_WIDTH+:INT_MAN_WIDTH];
			// Trace: macro expansion of FFL at design.sv:49534:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49534:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49534:269
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49534:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49534:556
						mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
			// Trace: macro expansion of FFL at design.sv:49535:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49535:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49535:269
					mid_pipe_src_is_int_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49535:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49535:556
						mid_pipe_src_is_int_q[i + 1] <= mid_pipe_src_is_int_q[i];
			// Trace: macro expansion of FFL at design.sv:49536:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49536:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49536:269
					mid_pipe_dst_is_int_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49536:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49536:556
						mid_pipe_dst_is_int_q[i + 1] <= mid_pipe_dst_is_int_q[i];
			// Trace: macro expansion of FFL at design.sv:49537:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49537:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49537:269
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49537:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49537:556
						mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= mid_pipe_info_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 8+:8];
			// Trace: macro expansion of FFL at design.sv:49538:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49538:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49538:269
					mid_pipe_mant_zero_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49538:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49538:556
						mid_pipe_mant_zero_q[i + 1] <= mid_pipe_mant_zero_q[i];
			// Trace: macro expansion of FFL at design.sv:49539:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49539:172
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49539:269
					mid_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49539:459
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49539:556
						mid_pipe_op_mod_q[i + 1] <= mid_pipe_op_mod_q[i];
			// Trace: macro expansion of FFL at design.sv:49540:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49540:184
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49540:281
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at design.sv:49540:471
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49540:568
						mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:49541:99
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49541:196
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49541:293
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_5D882(0);
				else
					// Trace: macro expansion of FFL at design.sv:49541:483
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49541:580
						mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:49542:99
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49542:196
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49542:293
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_5D882(0);
				else
					// Trace: macro expansion of FFL at design.sv:49542:483
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49542:580
						mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:49543:100
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49543:197
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49543:294
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_CDB06(0);
				else
					// Trace: macro expansion of FFL at design.sv:49543:484
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49543:581
						mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:49544:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49544:182
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49544:279
					mid_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:49544:469
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49544:566
						mid_pipe_tag_q[i + 1] <= mid_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:49545:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49545:182
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49545:279
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_533F1(1'sb0);
				else
					// Trace: macro expansion of FFL at design.sv:49545:469
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49545:566
						mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
		end
	endgenerate
	// Trace: design.sv:49548:3
	assign input_sign_q = mid_pipe_input_sign_q[NUM_MID_REGS];
	// Trace: design.sv:49549:3
	assign input_exp_q = mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: design.sv:49550:3
	assign input_mant_q = mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	// Trace: design.sv:49551:3
	assign destination_exp_q = mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: design.sv:49552:3
	assign src_is_int_q = mid_pipe_src_is_int_q[NUM_MID_REGS];
	// Trace: design.sv:49553:3
	assign dst_is_int_q = mid_pipe_dst_is_int_q[NUM_MID_REGS];
	// Trace: design.sv:49554:3
	assign info_q = mid_pipe_info_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 8+:8];
	// Trace: design.sv:49555:3
	assign mant_is_zero_q = mid_pipe_mant_zero_q[NUM_MID_REGS];
	// Trace: design.sv:49556:3
	assign op_mod_q2 = mid_pipe_op_mod_q[NUM_MID_REGS];
	// Trace: design.sv:49557:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: design.sv:49558:3
	assign src_fmt_q2 = mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: design.sv:49559:3
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: design.sv:49560:3
	assign int_fmt_q2 = mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	// Trace: design.sv:49565:3
	reg [INT_EXP_WIDTH - 1:0] final_exp;
	// Trace: design.sv:49567:3
	reg [2 * INT_MAN_WIDTH:0] preshift_mant;
	// Trace: design.sv:49568:3
	wire [2 * INT_MAN_WIDTH:0] destination_mant;
	// Trace: design.sv:49569:3
	wire [SUPER_MAN_BITS - 1:0] final_mant;
	// Trace: design.sv:49570:3
	wire [MAX_INT_WIDTH - 1:0] final_int;
	// Trace: design.sv:49572:3
	reg [$clog2(INT_MAN_WIDTH + 1) - 1:0] denorm_shamt;
	// Trace: design.sv:49574:3
	wire [1:0] fp_round_sticky_bits;
	wire [1:0] int_round_sticky_bits;
	wire [1:0] round_sticky_bits;
	// Trace: design.sv:49575:3
	reg of_before_round;
	reg uf_before_round;
	// Trace: design.sv:49579:3
	always @(*) begin : cast_value
		if (_sv2v_0)
			;
		// Trace: design.sv:49581:5
		final_exp = $unsigned(destination_exp_q);
		// Trace: design.sv:49582:5
		preshift_mant = 1'sb0;
		// Trace: design.sv:49583:5
		denorm_shamt = SUPER_MAN_BITS - fpnew_pkg_man_bits(dst_fmt_q2);
		// Trace: design.sv:49584:5
		of_before_round = 1'b0;
		// Trace: design.sv:49585:5
		uf_before_round = 1'b0;
		// Trace: design.sv:49588:5
		preshift_mant = input_mant_q << (INT_MAN_WIDTH + 1);
		// Trace: design.sv:49591:5
		if (dst_is_int_q) begin
			// Trace: design.sv:49593:7
			denorm_shamt = $unsigned((MAX_INT_WIDTH - 1) - input_exp_q);
			// Trace: design.sv:49595:7
			if (input_exp_q >= $signed((fpnew_pkg_int_width(int_fmt_q2) - 1) + op_mod_q2)) begin
				// Trace: design.sv:49596:9
				denorm_shamt = 1'sb0;
				// Trace: design.sv:49597:9
				of_before_round = 1'b1;
			end
			else if (input_exp_q < -1) begin
				// Trace: design.sv:49600:9
				denorm_shamt = MAX_INT_WIDTH + 1;
				// Trace: design.sv:49601:9
				uf_before_round = 1'b1;
			end
		end
		else
			// Trace: design.sv:49606:7
			if ((destination_exp_q >= ($signed(2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1)) || (~src_is_int_q && info_q[4])) begin
				// Trace: design.sv:49608:9
				final_exp = $unsigned((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 2);
				// Trace: design.sv:49609:9
				preshift_mant = 1'sb1;
				// Trace: design.sv:49610:9
				of_before_round = 1'b1;
			end
			else if ((destination_exp_q < 1) && (destination_exp_q >= -$signed(fpnew_pkg_man_bits(dst_fmt_q2)))) begin
				// Trace: design.sv:49614:9
				final_exp = 1'sb0;
				// Trace: design.sv:49615:9
				denorm_shamt = $unsigned((denorm_shamt + 1) - destination_exp_q);
				// Trace: design.sv:49616:9
				uf_before_round = 1'b1;
			end
			else if (destination_exp_q < -$signed(fpnew_pkg_man_bits(dst_fmt_q2))) begin
				// Trace: design.sv:49619:9
				final_exp = 1'sb0;
				// Trace: design.sv:49620:9
				denorm_shamt = $unsigned((denorm_shamt + 2) + fpnew_pkg_man_bits(dst_fmt_q2));
				// Trace: design.sv:49621:9
				uf_before_round = 1'b1;
			end
	end
	// Trace: design.sv:49626:3
	localparam NUM_FP_STICKY = ((2 * INT_MAN_WIDTH) - SUPER_MAN_BITS) - 1;
	// Trace: design.sv:49627:3
	localparam NUM_INT_STICKY = (2 * INT_MAN_WIDTH) - MAX_INT_WIDTH;
	// Trace: design.sv:49630:3
	assign destination_mant = preshift_mant >> denorm_shamt;
	// Trace: design.sv:49632:3
	assign {final_mant, fp_round_sticky_bits[1]} = destination_mant[(2 * INT_MAN_WIDTH) - 1-:SUPER_MAN_BITS + 1];
	// Trace: design.sv:49634:3
	assign {final_int, int_round_sticky_bits[1]} = destination_mant[2 * INT_MAN_WIDTH-:MAX_INT_WIDTH + 1];
	// Trace: design.sv:49636:3
	assign fp_round_sticky_bits[0] = |{destination_mant[NUM_FP_STICKY - 1:0]};
	// Trace: design.sv:49637:3
	assign int_round_sticky_bits[0] = |{destination_mant[NUM_INT_STICKY - 1:0]};
	// Trace: design.sv:49640:3
	assign round_sticky_bits = (dst_is_int_q ? int_round_sticky_bits : fp_round_sticky_bits);
	// Trace: design.sv:49645:3
	wire [WIDTH - 1:0] pre_round_abs;
	// Trace: design.sv:49646:3
	wire of_after_round;
	// Trace: design.sv:49647:3
	wire uf_after_round;
	// Trace: design.sv:49649:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_pre_round_abs;
	// Trace: design.sv:49650:3
	reg [4:0] fmt_of_after_round;
	// Trace: design.sv:49651:3
	reg [4:0] fmt_uf_after_round;
	// Trace: design.sv:49653:3
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_pre_round_abs;
	// Trace: design.sv:49655:3
	wire rounded_sign;
	// Trace: design.sv:49656:3
	wire [WIDTH - 1:0] rounded_abs;
	// Trace: design.sv:49657:3
	wire result_true_zero;
	// Trace: design.sv:49659:3
	wire [WIDTH - 1:0] rounded_int_res;
	// Trace: design.sv:49660:3
	wire rounded_int_res_zero;
	// Trace: design.sv:49664:3
	genvar _gv_fmt_2;
	generate
		for (_gv_fmt_2 = 0; _gv_fmt_2 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_2 = _gv_fmt_2 + 1) begin : gen_res_assemble
			localparam fmt = _gv_fmt_2;
			// Trace: design.sv:49666:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:49667:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_5D882(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: design.sv:49670:7
				always @(*) begin : assemble_result
					if (_sv2v_0)
						;
					// Trace: design.sv:49671:9
					fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = {final_exp[EXP_BITS - 1:0], final_mant[MAN_BITS - 1:0]};
				end
			end
			else begin : inactive_format
				// Trace: design.sv:49674:7
				wire [WIDTH * 1:1] sv2v_tmp_DA55D;
				assign sv2v_tmp_DA55D = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = sv2v_tmp_DA55D;
			end
		end
	endgenerate
	// Trace: design.sv:49679:3
	genvar _gv_ifmt_2;
	generate
		for (_gv_ifmt_2 = 0; _gv_ifmt_2 < sv2v_cast_32_signed(NUM_INT_FORMATS); _gv_ifmt_2 = _gv_ifmt_2 + 1) begin : gen_int_res_sign_ext
			localparam ifmt = _gv_ifmt_2;
			// Trace: design.sv:49681:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_CDB06(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: design.sv:49684:7
				always @(*) begin : assemble_result
					if (_sv2v_0)
						;
					// Trace: design.sv:49686:9
					ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = {WIDTH {final_int[INT_WIDTH - 1]}};
					// Trace: design.sv:49687:9
					ifmt_pre_round_abs[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = final_int[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				// Trace: design.sv:49690:7
				wire [WIDTH * 1:1] sv2v_tmp_7C8AF;
				assign sv2v_tmp_7C8AF = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = sv2v_tmp_7C8AF;
			end
		end
	endgenerate
	// Trace: design.sv:49695:3
	assign pre_round_abs = (dst_is_int_q ? ifmt_pre_round_abs[int_fmt_q2 * WIDTH+:WIDTH] : fmt_pre_round_abs[dst_fmt_q2 * WIDTH+:WIDTH]);
	// Trace: design.sv:49697:3
	fpnew_rounding #(.AbsWidth(WIDTH)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(input_sign_q),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(1'b0),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_true_zero)
	);
	// Trace: design.sv:49710:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	// Trace: design.sv:49713:3
	genvar _gv_fmt_3;
	generate
		for (_gv_fmt_3 = 0; _gv_fmt_3 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_3 = _gv_fmt_3 + 1) begin : gen_sign_inject
			localparam fmt = _gv_fmt_3;
			// Trace: design.sv:49715:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			// Trace: design.sv:49716:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:49717:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_5D882(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: design.sv:49720:7
				always @(*) begin : post_process
					if (_sv2v_0)
						;
					// Trace: design.sv:49722:9
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					// Trace: design.sv:49723:9
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					// Trace: design.sv:49726:9
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: design.sv:49727:9
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = (src_is_int_q & mant_is_zero_q ? {FP_WIDTH * 1 {1'sb0}} : {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]});
				end
			end
			else begin : inactive_format
				// Trace: design.sv:49732:7
				wire [1:1] sv2v_tmp_4C394;
				assign sv2v_tmp_4C394 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4C394;
				// Trace: design.sv:49733:7
				wire [1:1] sv2v_tmp_5852E;
				assign sv2v_tmp_5852E = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_5852E;
				// Trace: design.sv:49734:7
				wire [WIDTH * 1:1] sv2v_tmp_F321A;
				assign sv2v_tmp_F321A = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_F321A;
			end
		end
	endgenerate
	// Trace: design.sv:49739:3
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	// Trace: design.sv:49740:3
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	// Trace: design.sv:49743:3
	assign rounded_int_res = (rounded_sign ? $unsigned(-rounded_abs) : rounded_abs);
	// Trace: design.sv:49744:3
	assign rounded_int_res_zero = rounded_int_res == {WIDTH {1'sb0}};
	// Trace: design.sv:49749:3
	wire [WIDTH - 1:0] fp_special_result;
	// Trace: design.sv:49750:3
	wire [4:0] fp_special_status;
	// Trace: design.sv:49751:3
	wire fp_result_is_special;
	// Trace: design.sv:49753:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	// Trace: design.sv:49756:3
	genvar _gv_fmt_4;
	generate
		for (_gv_fmt_4 = 0; _gv_fmt_4 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_4 = _gv_fmt_4 + 1) begin : gen_special_results
			localparam fmt = _gv_fmt_4;
			// Trace: design.sv:49758:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			// Trace: design.sv:49759:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:49760:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:49762:5
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			// Trace: design.sv:49763:5
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: design.sv:49766:7
				always @(*) begin : special_results
					// Trace: design.sv:49767:9
					reg [FP_WIDTH - 1:0] special_res;
					if (_sv2v_0)
						;
					// Trace: design.sv:49768:9
					special_res = (info_q[5] ? input_sign_q << (FP_WIDTH - 1) : {1'b0, QNAN_EXPONENT, QNAN_MANTISSA});
					// Trace: design.sv:49773:9
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: design.sv:49774:9
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: design.sv:49777:7
				wire [WIDTH * 1:1] sv2v_tmp_294DC;
				assign sv2v_tmp_294DC = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_294DC;
			end
		end
	endgenerate
	// Trace: design.sv:49782:3
	assign fp_result_is_special = ~src_is_int_q & ((info_q[5] | info_q[3]) | ~info_q[0]);
	// Trace: design.sv:49787:3
	assign fp_special_status = {info_q[2], 4'b0000};
	// Trace: design.sv:49790:3
	assign fp_special_result = fmt_special_result[dst_fmt_q2 * WIDTH+:WIDTH];
	// Trace: design.sv:49795:3
	wire [WIDTH - 1:0] int_special_result;
	// Trace: design.sv:49796:3
	wire [4:0] int_special_status;
	// Trace: design.sv:49797:3
	wire int_result_is_special;
	// Trace: design.sv:49799:3
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_special_result;
	// Trace: design.sv:49802:3
	genvar _gv_ifmt_3;
	generate
		for (_gv_ifmt_3 = 0; _gv_ifmt_3 < sv2v_cast_32_signed(NUM_INT_FORMATS); _gv_ifmt_3 = _gv_ifmt_3 + 1) begin : gen_special_results_int
			localparam ifmt = _gv_ifmt_3;
			// Trace: design.sv:49804:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_CDB06(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: design.sv:49807:7
				always @(*) begin : special_results
					// Trace: design.sv:49808:9
					reg [INT_WIDTH - 1:0] special_res;
					if (_sv2v_0)
						;
					// Trace: design.sv:49811:9
					special_res[INT_WIDTH - 2:0] = 1'sb1;
					// Trace: design.sv:49812:9
					special_res[INT_WIDTH - 1] = op_mod_q2;
					// Trace: design.sv:49815:9
					if (input_sign_q && !info_q[3])
						// Trace: design.sv:49816:11
						special_res = ~special_res;
					// Trace: design.sv:49819:9
					ifmt_special_result[ifmt * WIDTH+:WIDTH] = {WIDTH {special_res[INT_WIDTH - 1]}};
					// Trace: design.sv:49820:9
					ifmt_special_result[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: design.sv:49823:7
				wire [WIDTH * 1:1] sv2v_tmp_577FA;
				assign sv2v_tmp_577FA = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_special_result[ifmt * WIDTH+:WIDTH] = sv2v_tmp_577FA;
			end
		end
	endgenerate
	// Trace: design.sv:49828:3
	assign int_result_is_special = (((info_q[3] | info_q[4]) | of_before_round) | ~info_q[0]) | ((input_sign_q & op_mod_q2) & ~rounded_int_res_zero);
	// Trace: design.sv:49833:3
	assign int_special_status = 5'b10000;
	// Trace: design.sv:49836:3
	assign int_special_result = ifmt_special_result[int_fmt_q2 * WIDTH+:WIDTH];
	// Trace: design.sv:49841:3
	wire [4:0] int_regular_status;
	wire [4:0] fp_regular_status;
	// Trace: design.sv:49843:3
	wire [WIDTH - 1:0] fp_result;
	wire [WIDTH - 1:0] int_result;
	// Trace: design.sv:49844:3
	wire [4:0] fp_status;
	wire [4:0] int_status;
	// Trace: design.sv:49846:3
	assign fp_regular_status[4] = src_is_int_q & (of_before_round | of_after_round);
	// Trace: design.sv:49847:3
	assign fp_regular_status[3] = 1'b0;
	// Trace: design.sv:49848:3
	assign fp_regular_status[2] = ~src_is_int_q & (~info_q[4] & (of_before_round | of_after_round));
	// Trace: design.sv:49849:3
	assign fp_regular_status[1] = uf_after_round & fp_regular_status[0];
	// Trace: design.sv:49850:3
	assign fp_regular_status[0] = (src_is_int_q ? |fp_round_sticky_bits : |fp_round_sticky_bits | (~info_q[4] & (of_before_round | of_after_round)));
	// Trace: design.sv:49852:3
	assign int_regular_status = {4'b0000, |int_round_sticky_bits};
	// Trace: design.sv:49854:3
	assign fp_result = (fp_result_is_special ? fp_special_result : fmt_result[dst_fmt_q2 * WIDTH+:WIDTH]);
	// Trace: design.sv:49855:3
	assign fp_status = (fp_result_is_special ? fp_special_status : fp_regular_status);
	// Trace: design.sv:49856:3
	assign int_result = (int_result_is_special ? int_special_result : rounded_int_res);
	// Trace: design.sv:49857:3
	assign int_status = (int_result_is_special ? int_special_status : int_regular_status);
	// Trace: design.sv:49860:3
	wire [WIDTH - 1:0] result_d;
	// Trace: design.sv:49861:3
	wire [4:0] status_d;
	// Trace: design.sv:49862:3
	wire extension_bit;
	// Trace: design.sv:49865:3
	assign result_d = (dst_is_int_q ? int_result : fp_result);
	// Trace: design.sv:49866:3
	assign status_d = (dst_is_int_q ? int_status : fp_status);
	// Trace: design.sv:49869:3
	assign extension_bit = (dst_is_int_q ? int_result[WIDTH - 1] : 1'b1);
	// Trace: design.sv:49875:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: design.sv:49876:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: design.sv:49877:3
	reg [0:NUM_OUT_REGS] out_pipe_ext_bit_q;
	// Trace: design.sv:49878:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: design.sv:49879:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: design.sv:49880:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: design.sv:49882:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: design.sv:49885:3
	wire [WIDTH * 1:1] sv2v_tmp_6C5BE;
	assign sv2v_tmp_6C5BE = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6C5BE;
	// Trace: design.sv:49886:3
	wire [5:1] sv2v_tmp_D9FFA;
	assign sv2v_tmp_D9FFA = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_D9FFA;
	// Trace: design.sv:49887:3
	wire [1:1] sv2v_tmp_F04C7;
	assign sv2v_tmp_F04C7 = extension_bit;
	always @(*) out_pipe_ext_bit_q[0] = sv2v_tmp_F04C7;
	// Trace: design.sv:49888:3
	wire [1:1] sv2v_tmp_1CCC3;
	assign sv2v_tmp_1CCC3 = mid_pipe_tag_q[NUM_MID_REGS];
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_1CCC3;
	// Trace: design.sv:49889:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_6EDB0;
	assign sv2v_tmp_6EDB0 = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_6EDB0;
	// Trace: design.sv:49890:3
	wire [1:1] sv2v_tmp_E45E7;
	assign sv2v_tmp_E45E7 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_E45E7;
	// Trace: design.sv:49892:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: design.sv:49894:3
	genvar _gv_i_71;
	generate
		for (_gv_i_71 = 0; _gv_i_71 < NUM_OUT_REGS; _gv_i_71 = _gv_i_71 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_71;
			// Trace: design.sv:49896:5
			wire reg_ena;
			// Trace: design.sv:49900:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:49902:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:49902:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:49902:485
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:49902:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:49902:715
						out_pipe_valid_q[i + 1] <= 1'b0;
					else if (out_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:49902:867
						out_pipe_valid_q[i + 1] <= out_pipe_valid_q[i];
			// Trace: design.sv:49904:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:49906:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49906:166
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49906:263
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49906:453
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49906:550
						out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH];
			// Trace: macro expansion of FFL at design.sv:49907:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49907:166
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49907:263
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49907:453
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49907:550
						out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5];
			// Trace: macro expansion of FFL at design.sv:49908:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49908:166
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49908:263
					out_pipe_ext_bit_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:49908:453
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49908:550
						out_pipe_ext_bit_q[i + 1] <= out_pipe_ext_bit_q[i];
			// Trace: macro expansion of FFL at design.sv:49909:79
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49909:176
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49909:273
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:49909:463
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49909:560
						out_pipe_tag_q[i + 1] <= out_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:49910:79
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:49910:176
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:49910:273
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_533F1(1'sb0);
				else
					// Trace: macro expansion of FFL at design.sv:49910:463
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:49910:560
						out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
		end
	endgenerate
	// Trace: design.sv:49913:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: design.sv:49915:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: design.sv:49916:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: design.sv:49917:3
	assign extension_bit_o = out_pipe_ext_bit_q[NUM_OUT_REGS];
	// Trace: design.sv:49918:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: design.sv:49919:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: design.sv:49920:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: design.sv:49921:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
	initial _sv2v_0 = 0;
endmodule
module fpnew_classifier (
	operands_i,
	is_boxed_i,
	info_o
);
	reg _sv2v_0;
	// Trace: design.sv:49939:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_5D882(0);
	// Trace: design.sv:49940:13
	parameter [31:0] NumOperands = 1;
	// Trace: design.sv:49942:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: design.sv:49944:3
	input wire [(NumOperands * WIDTH) - 1:0] operands_i;
	// Trace: design.sv:49945:3
	input wire [NumOperands - 1:0] is_boxed_i;
	// Trace: design.sv:49946:3
	// removed localparam type fpnew_pkg_fp_info_t
	output reg [(NumOperands * 8) - 1:0] info_o;
	// Trace: design.sv:49949:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:326:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:327:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: design.sv:49950:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:331:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:332:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: design.sv:49953:3
	// removed localparam type fp_t
	// Trace: design.sv:49960:3
	genvar _gv_op_1;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_op_1 = 0; _gv_op_1 < sv2v_cast_32_signed(NumOperands); _gv_op_1 = _gv_op_1 + 1) begin : gen_num_values
			localparam op = _gv_op_1;
			// Trace: design.sv:49962:5
			reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] value;
			// Trace: design.sv:49963:5
			reg is_boxed;
			// Trace: design.sv:49964:5
			reg is_normal;
			// Trace: design.sv:49965:5
			reg is_inf;
			// Trace: design.sv:49966:5
			reg is_nan;
			// Trace: design.sv:49967:5
			reg is_signalling;
			// Trace: design.sv:49968:5
			reg is_quiet;
			// Trace: design.sv:49969:5
			reg is_zero;
			// Trace: design.sv:49970:5
			reg is_subnormal;
			// Trace: design.sv:49975:5
			always @(*) begin : classify_input
				if (_sv2v_0)
					;
				// Trace: design.sv:49976:7
				value = operands_i[op * WIDTH+:WIDTH];
				// Trace: design.sv:49977:7
				is_boxed = is_boxed_i[op];
				// Trace: design.sv:49978:7
				is_normal = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] != {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] != {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}});
				// Trace: design.sv:49979:7
				is_zero = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && (value[MAN_BITS - 1-:MAN_BITS] == {MAN_BITS * 1 {1'sb0}});
				// Trace: design.sv:49980:7
				is_subnormal = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && !is_zero;
				// Trace: design.sv:49981:7
				is_inf = is_boxed && ((value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}}) && (value[MAN_BITS - 1-:MAN_BITS] == {MAN_BITS * 1 {1'sb0}}));
				// Trace: design.sv:49982:7
				is_nan = !is_boxed || ((value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}}) && (value[MAN_BITS - 1-:MAN_BITS] != {MAN_BITS * 1 {1'sb0}}));
				// Trace: design.sv:49983:7
				is_signalling = (is_boxed && is_nan) && (value[(MAN_BITS - 1) - ((MAN_BITS - 1) - (MAN_BITS - 1))] == 1'b0);
				// Trace: design.sv:49984:7
				is_quiet = is_nan && !is_signalling;
				// Trace: design.sv:49986:7
				info_o[(op * 8) + 7] = is_normal;
				// Trace: design.sv:49987:7
				info_o[(op * 8) + 6] = is_subnormal;
				// Trace: design.sv:49988:7
				info_o[(op * 8) + 5] = is_zero;
				// Trace: design.sv:49989:7
				info_o[(op * 8) + 4] = is_inf;
				// Trace: design.sv:49990:7
				info_o[(op * 8) + 3] = is_nan;
				// Trace: design.sv:49991:7
				info_o[(op * 8) + 2] = is_signalling;
				// Trace: design.sv:49992:7
				info_o[(op * 8) + 1] = is_quiet;
				// Trace: design.sv:49993:7
				info_o[op * 8] = is_boxed;
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module fpnew_divsqrt_multi_E225A_955F4 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	dst_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	reg _sv2v_0;
	// Trace: design.sv:50015:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: design.sv:50017:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: design.sv:50018:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd1;
	// Trace: design.sv:50019:38
	// removed localparam type TagType
	// Trace: design.sv:50020:38
	// removed localparam type AuxType
	// Trace: design.sv:50022:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:34
		input reg signed [31:0] a;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:41
		input reg signed [31:0] b;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:296:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:308:48
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:309:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:5
			begin : sv2v_autoblock_1
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:312:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: design.sv:50023:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: design.sv:50025:3
	input wire clk_i;
	// Trace: design.sv:50026:3
	input wire rst_ni;
	// Trace: design.sv:50028:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: design.sv:50029:3
	input wire [9:0] is_boxed_i;
	// Trace: design.sv:50030:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:50031:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:50032:3
	input wire [2:0] dst_fmt_i;
	// Trace: design.sv:50033:3
	input wire tag_i;
	// Trace: design.sv:50034:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: design.sv:50036:3
	input wire in_valid_i;
	// Trace: design.sv:50037:3
	output wire in_ready_o;
	// Trace: design.sv:50038:3
	input wire flush_i;
	// Trace: design.sv:50040:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: design.sv:50041:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: design.sv:50042:3
	output wire extension_bit_o;
	// Trace: design.sv:50043:3
	output wire tag_o;
	// Trace: design.sv:50044:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: design.sv:50046:3
	output wire out_valid_o;
	// Trace: design.sv:50047:3
	input wire out_ready_i;
	// Trace: design.sv:50049:3
	output wire busy_o;
	// Trace: design.sv:50056:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: design.sv:50061:3
	localparam NUM_OUT_REGS = ((PipeConfig == 2'd1) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: design.sv:50071:3
	wire [(2 * WIDTH) - 1:0] operands_q;
	// Trace: design.sv:50072:3
	wire [2:0] rnd_mode_q;
	// Trace: design.sv:50073:3
	wire [3:0] op_q;
	// Trace: design.sv:50074:3
	wire [2:0] dst_fmt_q;
	// Trace: design.sv:50075:3
	wire in_valid_q;
	// Trace: design.sv:50078:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: design.sv:50079:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: design.sv:50080:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: design.sv:50081:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: design.sv:50082:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: design.sv:50083:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: design.sv:50084:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: design.sv:50086:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: design.sv:50089:3
	wire [2 * WIDTH:1] sv2v_tmp_44D18;
	assign sv2v_tmp_44D18 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_44D18;
	// Trace: design.sv:50090:3
	wire [3:1] sv2v_tmp_27FE8;
	assign sv2v_tmp_27FE8 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_27FE8;
	// Trace: design.sv:50091:3
	wire [4:1] sv2v_tmp_72726;
	assign sv2v_tmp_72726 = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_72726;
	// Trace: design.sv:50092:3
	wire [3:1] sv2v_tmp_014AE;
	assign sv2v_tmp_014AE = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_014AE;
	// Trace: design.sv:50093:3
	wire [1:1] sv2v_tmp_DE624;
	assign sv2v_tmp_DE624 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_DE624;
	// Trace: design.sv:50094:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_42C02;
	assign sv2v_tmp_42C02 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_42C02;
	// Trace: design.sv:50095:3
	wire [1:1] sv2v_tmp_CFC25;
	assign sv2v_tmp_CFC25 = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_CFC25;
	// Trace: design.sv:50097:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: design.sv:50099:3
	genvar _gv_i_72;
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_533F1;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_533F1 = inp;
	endfunction
	generate
		for (_gv_i_72 = 0; _gv_i_72 < NUM_INP_REGS; _gv_i_72 = _gv_i_72 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_72;
			// Trace: design.sv:50101:5
			wire reg_ena;
			// Trace: design.sv:50105:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:50107:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:50107:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:50107:485
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:50107:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:50107:715
						inp_pipe_valid_q[i + 1] <= 1'b0;
					else if (inp_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:50107:867
						inp_pipe_valid_q[i + 1] <= inp_pipe_valid_q[i];
			// Trace: design.sv:50109:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:50111:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50111:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50111:265
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50111:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50111:552
						inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2];
			// Trace: macro expansion of FFL at design.sv:50112:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50112:180
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50112:277
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at design.sv:50112:467
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50112:564
						inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:50113:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50113:182
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50113:279
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_4CD2E(0);
				else
					// Trace: macro expansion of FFL at design.sv:50113:469
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50113:566
						inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
			// Trace: macro expansion of FFL at design.sv:50114:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50114:192
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50114:289
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_5D882(0);
				else
					// Trace: macro expansion of FFL at design.sv:50114:479
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50114:576
						inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:50115:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50115:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50115:275
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:50115:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50115:562
						inp_pipe_tag_q[i + 1] <= inp_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:50116:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50116:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50116:275
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_533F1(1'sb0);
				else
					// Trace: macro expansion of FFL at design.sv:50116:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50116:562
						inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
		end
	endgenerate
	// Trace: design.sv:50119:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2];
	// Trace: design.sv:50120:3
	assign rnd_mode_q = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	// Trace: design.sv:50121:3
	assign op_q = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
	// Trace: design.sv:50122:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: design.sv:50123:3
	assign in_valid_q = inp_pipe_valid_q[NUM_INP_REGS];
	// Trace: design.sv:50128:3
	reg [1:0] divsqrt_fmt;
	// Trace: design.sv:50129:3
	reg [127:0] divsqrt_operands;
	// Trace: design.sv:50130:3
	reg input_is_fp8;
	// Trace: design.sv:50133:3
	always @(*) begin : translate_fmt
		if (_sv2v_0)
			;
		// Trace: design.sv:50134:5
		(* full_case, parallel_case *)
		case (dst_fmt_q)
			sv2v_cast_5D882('d0):
				// Trace: design.sv:50135:27
				divsqrt_fmt = 2'b00;
			sv2v_cast_5D882('d1):
				// Trace: design.sv:50136:27
				divsqrt_fmt = 2'b01;
			sv2v_cast_5D882('d2):
				// Trace: design.sv:50137:27
				divsqrt_fmt = 2'b10;
			sv2v_cast_5D882('d4):
				// Trace: design.sv:50138:27
				divsqrt_fmt = 2'b11;
			default:
				// Trace: design.sv:50139:27
				divsqrt_fmt = 2'b10;
		endcase
		// Trace: design.sv:50143:5
		input_is_fp8 = FpFmtConfig[sv2v_cast_5D882('d3)] & (dst_fmt_q == sv2v_cast_5D882('d3));
		// Trace: design.sv:50146:5
		divsqrt_operands[0+:64] = (input_is_fp8 ? operands_q[0+:WIDTH] << 8 : operands_q[0+:WIDTH]);
		// Trace: design.sv:50147:5
		divsqrt_operands[64+:64] = (input_is_fp8 ? operands_q[WIDTH+:WIDTH] << 8 : operands_q[WIDTH+:WIDTH]);
	end
	// Trace: design.sv:50153:3
	reg in_ready;
	// Trace: design.sv:50154:3
	wire div_valid;
	wire sqrt_valid;
	// Trace: design.sv:50155:3
	wire unit_ready;
	wire unit_done;
	// Trace: design.sv:50156:3
	wire op_starting;
	// Trace: design.sv:50157:3
	reg out_valid;
	wire out_ready;
	// Trace: design.sv:50158:3
	reg hold_result;
	// Trace: design.sv:50159:3
	reg data_is_held;
	// Trace: design.sv:50160:3
	reg unit_busy;
	// Trace: design.sv:50162:3
	// removed localparam type fsm_state_e
	// Trace: design.sv:50163:3
	reg [1:0] state_q;
	reg [1:0] state_d;
	// Trace: design.sv:50166:3
	assign inp_pipe_ready[NUM_INP_REGS] = in_ready;
	// Trace: design.sv:50169:3
	assign div_valid = ((in_valid_q & (op_q == sv2v_cast_4CD2E(4))) & in_ready) & ~flush_i;
	// Trace: design.sv:50170:3
	assign sqrt_valid = ((in_valid_q & (op_q != sv2v_cast_4CD2E(4))) & in_ready) & ~flush_i;
	// Trace: design.sv:50171:3
	assign op_starting = div_valid | sqrt_valid;
	// Trace: design.sv:50174:3
	always @(*) begin : flag_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:50176:5
		in_ready = 1'b0;
		// Trace: design.sv:50177:5
		out_valid = 1'b0;
		// Trace: design.sv:50178:5
		hold_result = 1'b0;
		// Trace: design.sv:50179:5
		data_is_held = 1'b0;
		// Trace: design.sv:50180:5
		unit_busy = 1'b0;
		// Trace: design.sv:50181:5
		state_d = state_q;
		// Trace: design.sv:50183:5
		(* full_case, parallel_case *)
		case (state_q)
			2'd0: begin
				// Trace: design.sv:50186:9
				in_ready = 1'b1;
				// Trace: design.sv:50187:9
				if (in_valid_q && unit_ready)
					// Trace: design.sv:50188:11
					state_d = 2'd1;
			end
			2'd1: begin
				// Trace: design.sv:50193:9
				unit_busy = 1'b1;
				// Trace: design.sv:50195:9
				if (unit_done) begin
					// Trace: design.sv:50196:11
					out_valid = 1'b1;
					// Trace: design.sv:50198:11
					if (out_ready) begin
						// Trace: design.sv:50199:13
						state_d = 2'd0;
						// Trace: design.sv:50200:13
						if (in_valid_q && unit_ready) begin
							// Trace: design.sv:50201:15
							in_ready = 1'b1;
							// Trace: design.sv:50202:15
							state_d = 2'd1;
						end
					end
					else begin
						// Trace: design.sv:50206:13
						hold_result = 1'b1;
						// Trace: design.sv:50207:13
						state_d = 2'd2;
					end
				end
			end
			2'd2: begin
				// Trace: design.sv:50213:9
				unit_busy = 1'b1;
				// Trace: design.sv:50214:9
				data_is_held = 1'b1;
				// Trace: design.sv:50215:9
				out_valid = 1'b1;
				// Trace: design.sv:50217:9
				if (out_ready) begin
					// Trace: design.sv:50218:11
					state_d = 2'd0;
					// Trace: design.sv:50219:11
					if (in_valid_q && unit_ready) begin
						// Trace: design.sv:50220:13
						in_ready = 1'b1;
						// Trace: design.sv:50221:13
						state_d = 2'd1;
					end
				end
			end
			default:
				// Trace: design.sv:50226:16
				state_d = 2'd0;
		endcase
		if (flush_i) begin
			// Trace: design.sv:50231:7
			unit_busy = 1'b0;
			// Trace: design.sv:50232:7
			out_valid = 1'b0;
			// Trace: design.sv:50233:7
			state_d = 2'd0;
		end
	end
	// Trace: macro expansion of FF at design.sv:50238:30
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at design.sv:50238:118
		if (!rst_ni)
			// Trace: macro expansion of FF at design.sv:50238:206
			state_q <= 2'd0;
		else
			// Trace: macro expansion of FF at design.sv:50238:378
			state_q <= state_d;
	// Trace: design.sv:50241:3
	reg result_is_fp8_q;
	// Trace: design.sv:50242:3
	reg result_tag_q;
	// Trace: design.sv:50243:3
	reg [AuxType_AUX_BITS - 1:0] result_aux_q;
	// Trace: macro expansion of FFL at design.sv:50246:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at design.sv:50246:167
		if (!rst_ni)
			// Trace: macro expansion of FFL at design.sv:50246:264
			result_is_fp8_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at design.sv:50246:454
			if (op_starting)
				// Trace: macro expansion of FFL at design.sv:50246:551
				result_is_fp8_q <= input_is_fp8;
	// Trace: macro expansion of FFL at design.sv:50247:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at design.sv:50247:167
		if (!rst_ni)
			// Trace: macro expansion of FFL at design.sv:50247:264
			result_tag_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at design.sv:50247:454
			if (op_starting)
				// Trace: macro expansion of FFL at design.sv:50247:551
				result_tag_q <= inp_pipe_tag_q[NUM_INP_REGS];
	// Trace: macro expansion of FFL at design.sv:50248:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at design.sv:50248:167
		if (!rst_ni)
			// Trace: macro expansion of FFL at design.sv:50248:264
			result_aux_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at design.sv:50248:454
			if (op_starting)
				// Trace: macro expansion of FFL at design.sv:50248:551
				result_aux_q <= inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: design.sv:50253:3
	wire [63:0] unit_result;
	// Trace: design.sv:50254:3
	wire [WIDTH - 1:0] adjusted_result;
	reg [WIDTH - 1:0] held_result_q;
	// Trace: design.sv:50255:3
	wire [4:0] unit_status;
	reg [4:0] held_status_q;
	// Trace: design.sv:50257:3
	div_sqrt_top_mvp i_divsqrt_lei(
		.Clk_CI(clk_i),
		.Rst_RBI(rst_ni),
		.Div_start_SI(div_valid),
		.Sqrt_start_SI(sqrt_valid),
		.Operand_a_DI(divsqrt_operands[0+:64]),
		.Operand_b_DI(divsqrt_operands[64+:64]),
		.RM_SI(rnd_mode_q),
		.Precision_ctl_SI(1'sb0),
		.Format_sel_SI(divsqrt_fmt),
		.Kill_SI(flush_i),
		.Result_DO(unit_result),
		.Fflags_SO(unit_status),
		.Ready_SO(unit_ready),
		.Done_SO(unit_done)
	);
	// Trace: design.sv:50275:3
	assign adjusted_result = (result_is_fp8_q ? unit_result >> 8 : unit_result);
	// Trace: macro expansion of FFLNR at design.sv:50278:58
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at design.sv:50278:100
		if (hold_result)
			// Trace: macro expansion of FFLNR at design.sv:50278:142
			held_result_q <= adjusted_result;
	// Trace: macro expansion of FFLNR at design.sv:50279:58
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at design.sv:50279:100
		if (hold_result)
			// Trace: macro expansion of FFLNR at design.sv:50279:142
			held_status_q <= unit_status;
	// Trace: design.sv:50284:3
	wire [WIDTH - 1:0] result_d;
	// Trace: design.sv:50285:3
	wire [4:0] status_d;
	// Trace: design.sv:50287:3
	assign result_d = (data_is_held ? held_result_q : adjusted_result);
	// Trace: design.sv:50288:3
	assign status_d = (data_is_held ? held_status_q : unit_status);
	// Trace: design.sv:50294:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: design.sv:50295:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: design.sv:50296:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: design.sv:50297:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: design.sv:50298:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: design.sv:50300:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: design.sv:50303:3
	wire [WIDTH * 1:1] sv2v_tmp_8E412;
	assign sv2v_tmp_8E412 = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_8E412;
	// Trace: design.sv:50304:3
	wire [5:1] sv2v_tmp_F3F80;
	assign sv2v_tmp_F3F80 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_F3F80;
	// Trace: design.sv:50305:3
	wire [1:1] sv2v_tmp_AFEEA;
	assign sv2v_tmp_AFEEA = result_tag_q;
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_AFEEA;
	// Trace: design.sv:50306:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_03F4C;
	assign sv2v_tmp_03F4C = result_aux_q;
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_03F4C;
	// Trace: design.sv:50307:3
	wire [1:1] sv2v_tmp_F96BC;
	assign sv2v_tmp_F96BC = out_valid;
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_F96BC;
	// Trace: design.sv:50309:3
	assign out_ready = out_pipe_ready[0];
	// Trace: design.sv:50311:3
	genvar _gv_i_73;
	generate
		for (_gv_i_73 = 0; _gv_i_73 < NUM_OUT_REGS; _gv_i_73 = _gv_i_73 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_73;
			// Trace: design.sv:50313:5
			wire reg_ena;
			// Trace: design.sv:50317:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:50319:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:50319:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:50319:485
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:50319:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:50319:715
						out_pipe_valid_q[i + 1] <= 1'b0;
					else if (out_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:50319:867
						out_pipe_valid_q[i + 1] <= out_pipe_valid_q[i];
			// Trace: design.sv:50321:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:50323:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50323:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50323:261
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50323:451
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50323:548
						out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH];
			// Trace: macro expansion of FFL at design.sv:50324:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50324:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50324:261
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50324:451
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50324:548
						out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5];
			// Trace: macro expansion of FFL at design.sv:50325:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50325:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50325:271
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:50325:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50325:558
						out_pipe_tag_q[i + 1] <= out_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:50326:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50326:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50326:271
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_533F1(1'sb0);
				else
					// Trace: macro expansion of FFL at design.sv:50326:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50326:558
						out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
		end
	endgenerate
	// Trace: design.sv:50329:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: design.sv:50331:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: design.sv:50332:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: design.sv:50333:3
	assign extension_bit_o = 1'b1;
	// Trace: design.sv:50334:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: design.sv:50335:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: design.sv:50336:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: design.sv:50337:3
	assign busy_o = |{inp_pipe_valid_q, unit_busy, out_pipe_valid_q};
	initial _sv2v_0 = 0;
endmodule
module fpnew_fma_EA93F (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	reg _sv2v_0;
	// Trace: design.sv:50357:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_5D882(0);
	// Trace: design.sv:50358:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: design.sv:50359:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: design.sv:50360:38
	// removed localparam type TagType
	// Trace: design.sv:50361:38
	// removed localparam type AuxType
	// Trace: design.sv:50363:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: design.sv:50365:3
	input wire clk_i;
	// Trace: design.sv:50366:3
	input wire rst_ni;
	// Trace: design.sv:50368:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: design.sv:50369:3
	input wire [2:0] is_boxed_i;
	// Trace: design.sv:50370:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:50371:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:50372:3
	input wire op_mod_i;
	// Trace: design.sv:50373:3
	input wire tag_i;
	// Trace: design.sv:50374:3
	input wire aux_i;
	// Trace: design.sv:50376:3
	input wire in_valid_i;
	// Trace: design.sv:50377:3
	output wire in_ready_o;
	// Trace: design.sv:50378:3
	input wire flush_i;
	// Trace: design.sv:50380:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: design.sv:50381:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: design.sv:50382:3
	output wire extension_bit_o;
	// Trace: design.sv:50383:3
	output wire tag_o;
	// Trace: design.sv:50384:3
	output wire aux_o;
	// Trace: design.sv:50386:3
	output wire out_valid_o;
	// Trace: design.sv:50387:3
	input wire out_ready_i;
	// Trace: design.sv:50389:3
	output wire busy_o;
	// Trace: design.sv:50395:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:326:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:327:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: design.sv:50396:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:331:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:332:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: design.sv:50397:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:336:40
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:337:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	localparam [31:0] BIAS = fpnew_pkg_bias(FpFormat);
	// Trace: design.sv:50399:3
	localparam [31:0] PRECISION_BITS = MAN_BITS + 1;
	// Trace: design.sv:50401:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: design.sv:50402:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: design.sv:50406:3
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:34
		input reg signed [31:0] a;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:41
		input reg signed [31:0] b;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:296:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	localparam [31:0] EXP_WIDTH = $unsigned(fpnew_pkg_maximum(EXP_BITS + 2, LZC_RESULT_WIDTH));
	// Trace: design.sv:50408:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 3);
	// Trace: design.sv:50410:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: design.sv:50415:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: design.sv:50420:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: design.sv:50429:3
	// removed localparam type fp_t
	// Trace: design.sv:50439:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: design.sv:50440:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_is_boxed_q;
	// Trace: design.sv:50441:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: design.sv:50442:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: design.sv:50443:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: design.sv:50444:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: design.sv:50445:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: design.sv:50446:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: design.sv:50448:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: design.sv:50451:3
	wire [3 * WIDTH:1] sv2v_tmp_15914;
	assign sv2v_tmp_15914 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_15914;
	// Trace: design.sv:50452:3
	wire [3:1] sv2v_tmp_3D994;
	assign sv2v_tmp_3D994 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_3D994;
	// Trace: design.sv:50453:3
	wire [3:1] sv2v_tmp_85314;
	assign sv2v_tmp_85314 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_85314;
	// Trace: design.sv:50454:3
	wire [4:1] sv2v_tmp_D905E;
	assign sv2v_tmp_D905E = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_D905E;
	// Trace: design.sv:50455:3
	wire [1:1] sv2v_tmp_72E02;
	assign sv2v_tmp_72E02 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_72E02;
	// Trace: design.sv:50456:3
	wire [1:1] sv2v_tmp_DE624;
	assign sv2v_tmp_DE624 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_DE624;
	// Trace: design.sv:50457:3
	wire [1:1] sv2v_tmp_683C4;
	assign sv2v_tmp_683C4 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_683C4;
	// Trace: design.sv:50458:3
	wire [1:1] sv2v_tmp_CFC25;
	assign sv2v_tmp_CFC25 = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_CFC25;
	// Trace: design.sv:50460:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: design.sv:50462:3
	genvar _gv_i_74;
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	generate
		for (_gv_i_74 = 0; _gv_i_74 < NUM_INP_REGS; _gv_i_74 = _gv_i_74 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_74;
			// Trace: design.sv:50464:5
			wire reg_ena;
			// Trace: design.sv:50468:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:50470:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:50470:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:50470:485
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:50470:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:50470:715
						inp_pipe_valid_q[i + 1] <= 1'b0;
					else if (inp_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:50470:867
						inp_pipe_valid_q[i + 1] <= inp_pipe_valid_q[i];
			// Trace: design.sv:50472:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:50474:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50474:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50474:265
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50474:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50474:552
						inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3];
			// Trace: macro expansion of FFL at design.sv:50475:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50475:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50475:265
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50475:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50475:552
						inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:50476:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50476:180
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50476:277
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at design.sv:50476:467
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50476:564
						inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:50477:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50477:182
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50477:279
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_4CD2E(0);
				else
					// Trace: macro expansion of FFL at design.sv:50477:469
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50477:566
						inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
			// Trace: macro expansion of FFL at design.sv:50478:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50478:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50478:265
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50478:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50478:552
						inp_pipe_op_mod_q[i + 1] <= inp_pipe_op_mod_q[i];
			// Trace: macro expansion of FFL at design.sv:50479:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50479:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50479:275
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:50479:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50479:562
						inp_pipe_tag_q[i + 1] <= inp_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:50480:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50480:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50480:275
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:50480:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50480:562
						inp_pipe_aux_q[i + 1] <= inp_pipe_aux_q[i];
		end
	endgenerate
	// Trace: design.sv:50486:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [23:0] info_q;
	// Trace: design.sv:50489:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(3)
	) i_class_inputs(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3]),
		.info_o(info_q)
	);
	// Trace: design.sv:50498:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_c;
	// Trace: design.sv:50499:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: design.sv:50513:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_51E93;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_51E93 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_78D38;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_78D38 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_89227;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_89227 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_D5F4C;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_D5F4C = inp;
	endfunction
	always @(*) begin : op_select
		if (_sv2v_0)
			;
		// Trace: design.sv:50516:5
		operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: design.sv:50517:5
		operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: design.sv:50518:5
		operand_c = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: design.sv:50519:5
		info_a = info_q[0+:8];
		// Trace: design.sv:50520:5
		info_b = info_q[8+:8];
		// Trace: design.sv:50521:5
		info_c = info_q[16+:8];
		// Trace: design.sv:50524:5
		operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] = operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: design.sv:50526:5
		(* full_case, parallel_case *)
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_4CD2E(0):
				;
			sv2v_cast_4CD2E(1):
				// Trace: design.sv:50528:26
				operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] = ~operand_a[1 + (EXP_BITS + (MAN_BITS - 1))];
			sv2v_cast_4CD2E(2): begin
				// Trace: design.sv:50530:9
				operand_a = {1'b0, sv2v_cast_51E93(BIAS), sv2v_cast_78D38(1'sb0)};
				// Trace: design.sv:50531:9
				info_a = 8'b10000001;
			end
			sv2v_cast_4CD2E(3): begin
				// Trace: design.sv:50534:9
				operand_c = {1'b1, sv2v_cast_89227(1'sb0), sv2v_cast_78D38(1'sb0)};
				// Trace: design.sv:50535:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: design.sv:50538:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
				// Trace: design.sv:50539:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
				// Trace: design.sv:50540:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
				// Trace: design.sv:50541:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: design.sv:50542:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: design.sv:50543:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: design.sv:50551:3
	wire any_operand_inf;
	// Trace: design.sv:50552:3
	wire any_operand_nan;
	// Trace: design.sv:50553:3
	wire signalling_nan;
	// Trace: design.sv:50554:3
	wire effective_subtraction;
	// Trace: design.sv:50555:3
	wire tentative_sign;
	// Trace: design.sv:50558:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: design.sv:50559:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: design.sv:50560:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: design.sv:50562:3
	assign effective_subtraction = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]) ^ operand_c[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: design.sv:50564:3
	assign tentative_sign = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: design.sv:50569:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result;
	// Trace: design.sv:50570:3
	reg [4:0] special_status;
	// Trace: design.sv:50571:3
	reg result_is_special;
	// Trace: design.sv:50573:3
	always @(*) begin : special_cases
		if (_sv2v_0)
			;
		// Trace: design.sv:50575:5
		special_result = {1'b0, sv2v_cast_89227(1'sb1), sv2v_cast_D5F4C(2 ** (MAN_BITS - 1))};
		// Trace: design.sv:50576:5
		special_status = 1'sb0;
		// Trace: design.sv:50577:5
		result_is_special = 1'b0;
		// Trace: design.sv:50583:5
		if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
			// Trace: design.sv:50584:7
			result_is_special = 1'b1;
			// Trace: design.sv:50585:7
			special_status[4] = 1'b1;
		end
		else if (any_operand_nan) begin
			// Trace: design.sv:50588:7
			result_is_special = 1'b1;
			// Trace: design.sv:50589:7
			special_status[4] = signalling_nan;
		end
		else if (any_operand_inf) begin
			// Trace: design.sv:50592:7
			result_is_special = 1'b1;
			// Trace: design.sv:50594:7
			if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
				// Trace: design.sv:50595:9
				special_status[4] = 1'b1;
			else if (info_a[4] || info_b[4])
				// Trace: design.sv:50599:9
				special_result = {operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_89227(1'sb1), sv2v_cast_78D38(1'sb0)};
			else if (info_c[4])
				// Trace: design.sv:50603:9
				special_result = {operand_c[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_89227(1'sb1), sv2v_cast_78D38(1'sb0)};
		end
	end
	// Trace: design.sv:50611:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: design.sv:50612:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: design.sv:50613:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: design.sv:50616:3
	assign exponent_a = $signed({1'b0, operand_a[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: design.sv:50617:3
	assign exponent_b = $signed({1'b0, operand_b[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: design.sv:50618:3
	assign exponent_c = $signed({1'b0, operand_c[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: design.sv:50622:3
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	// Trace: design.sv:50624:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(BIAS) : $signed((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - $signed(BIAS)));
	// Trace: design.sv:50630:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: design.sv:50632:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	// Trace: design.sv:50635:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: design.sv:50637:3
	always @(*) begin : addend_shift_amount
		if (_sv2v_0)
			;
		// Trace: design.sv:50639:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: design.sv:50640:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: design.sv:50643:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: design.sv:50646:7
			addend_shamt = 0;
	end
	// Trace: design.sv:50652:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: design.sv:50653:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: design.sv:50654:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: design.sv:50657:3
	assign mantissa_a = {info_a[7], operand_a[MAN_BITS - 1-:MAN_BITS]};
	// Trace: design.sv:50658:3
	assign mantissa_b = {info_b[7], operand_b[MAN_BITS - 1-:MAN_BITS]};
	// Trace: design.sv:50659:3
	assign mantissa_c = {info_c[7], operand_c[MAN_BITS - 1-:MAN_BITS]};
	// Trace: design.sv:50662:3
	assign product = mantissa_a * mantissa_b;
	// Trace: design.sv:50667:3
	assign product_shifted = product << 2;
	// Trace: design.sv:50672:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: design.sv:50673:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: design.sv:50674:3
	wire sticky_before_add;
	// Trace: design.sv:50675:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: design.sv:50676:3
	wire inject_carry_in;
	// Trace: design.sv:50686:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: design.sv:50689:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: design.sv:50693:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: design.sv:50694:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: design.sv:50699:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	// Trace: design.sv:50700:3
	wire sum_carry;
	// Trace: design.sv:50701:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: design.sv:50702:3
	wire final_sign;
	// Trace: design.sv:50705:3
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: design.sv:50706:3
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	// Trace: design.sv:50709:3
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	// Trace: design.sv:50712:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: design.sv:50720:3
	wire effective_subtraction_q;
	// Trace: design.sv:50721:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: design.sv:50722:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: design.sv:50723:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: design.sv:50724:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: design.sv:50725:3
	wire sticky_before_add_q;
	// Trace: design.sv:50726:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: design.sv:50727:3
	wire final_sign_q;
	// Trace: design.sv:50728:3
	wire [2:0] rnd_mode_q;
	// Trace: design.sv:50729:3
	wire result_is_special_q;
	// Trace: design.sv:50730:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result_q;
	// Trace: design.sv:50731:3
	wire [4:0] special_status_q;
	// Trace: design.sv:50733:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: design.sv:50734:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: design.sv:50735:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: design.sv:50736:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: design.sv:50737:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: design.sv:50738:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: design.sv:50739:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: design.sv:50740:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: design.sv:50741:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: design.sv:50742:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: design.sv:50743:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: design.sv:50744:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: design.sv:50745:3
	reg [0:NUM_MID_REGS] mid_pipe_tag_q;
	// Trace: design.sv:50746:3
	reg [0:NUM_MID_REGS] mid_pipe_aux_q;
	// Trace: design.sv:50747:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: design.sv:50749:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: design.sv:50752:3
	wire [1:1] sv2v_tmp_301F1;
	assign sv2v_tmp_301F1 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_301F1;
	// Trace: design.sv:50753:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_27C8D;
	assign sv2v_tmp_27C8D = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_27C8D;
	// Trace: design.sv:50754:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_DEAE0;
	assign sv2v_tmp_DEAE0 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_DEAE0;
	// Trace: design.sv:50755:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_530A2;
	assign sv2v_tmp_530A2 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_530A2;
	// Trace: design.sv:50756:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_12F7F;
	assign sv2v_tmp_12F7F = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_12F7F;
	// Trace: design.sv:50757:3
	wire [1:1] sv2v_tmp_6A24C;
	assign sv2v_tmp_6A24C = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6A24C;
	// Trace: design.sv:50758:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_A48E2;
	assign sv2v_tmp_A48E2 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_A48E2;
	// Trace: design.sv:50759:3
	wire [1:1] sv2v_tmp_9C379;
	assign sv2v_tmp_9C379 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_9C379;
	// Trace: design.sv:50760:3
	wire [3:1] sv2v_tmp_C990F;
	assign sv2v_tmp_C990F = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_C990F;
	// Trace: design.sv:50761:3
	wire [1:1] sv2v_tmp_08378;
	assign sv2v_tmp_08378 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_08378;
	// Trace: design.sv:50762:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_8913F;
	assign sv2v_tmp_8913F = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_8913F;
	// Trace: design.sv:50763:3
	wire [5:1] sv2v_tmp_9D338;
	assign sv2v_tmp_9D338 = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_9D338;
	// Trace: design.sv:50764:3
	wire [1:1] sv2v_tmp_7259D;
	assign sv2v_tmp_7259D = inp_pipe_tag_q[NUM_INP_REGS];
	always @(*) mid_pipe_tag_q[0] = sv2v_tmp_7259D;
	// Trace: design.sv:50765:3
	wire [1:1] sv2v_tmp_8CE3D;
	assign sv2v_tmp_8CE3D = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) mid_pipe_aux_q[0] = sv2v_tmp_8CE3D;
	// Trace: design.sv:50766:3
	wire [1:1] sv2v_tmp_C7159;
	assign sv2v_tmp_C7159 = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_C7159;
	// Trace: design.sv:50768:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: design.sv:50771:3
	genvar _gv_i_75;
	generate
		for (_gv_i_75 = 0; _gv_i_75 < NUM_MID_REGS; _gv_i_75 = _gv_i_75 + 1) begin : gen_inside_pipeline
			localparam i = _gv_i_75;
			// Trace: design.sv:50773:5
			wire reg_ena;
			// Trace: design.sv:50777:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:50779:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:50779:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:50779:485
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:50779:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:50779:715
						mid_pipe_valid_q[i + 1] <= 1'b0;
					else if (mid_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:50779:867
						mid_pipe_valid_q[i + 1] <= mid_pipe_valid_q[i];
			// Trace: design.sv:50781:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:50783:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50783:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50783:271
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50783:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50783:558
						mid_pipe_eff_sub_q[i + 1] <= mid_pipe_eff_sub_q[i];
			// Trace: macro expansion of FFL at design.sv:50784:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50784:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50784:271
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50784:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50784:558
						mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH];
			// Trace: macro expansion of FFL at design.sv:50785:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50785:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50785:271
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50785:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50785:558
						mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH];
			// Trace: macro expansion of FFL at design.sv:50786:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50786:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50786:271
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50786:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50786:558
						mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH];
			// Trace: macro expansion of FFL at design.sv:50787:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50787:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50787:271
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50787:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50787:558
						mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
			// Trace: macro expansion of FFL at design.sv:50788:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50788:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50788:271
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50788:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50788:558
						mid_pipe_sticky_q[i + 1] <= mid_pipe_sticky_q[i];
			// Trace: macro expansion of FFL at design.sv:50789:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50789:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50789:271
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50789:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50789:558
						mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
			// Trace: macro expansion of FFL at design.sv:50790:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50790:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50790:271
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50790:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50790:558
						mid_pipe_final_sign_q[i + 1] <= mid_pipe_final_sign_q[i];
			// Trace: macro expansion of FFL at design.sv:50791:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50791:186
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50791:283
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at design.sv:50791:473
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50791:570
						mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:50792:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50792:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50792:271
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50792:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50792:558
						mid_pipe_res_is_spec_q[i + 1] <= mid_pipe_res_is_spec_q[i];
			// Trace: macro expansion of FFL at design.sv:50793:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50793:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50793:271
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50793:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50793:558
						mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
			// Trace: macro expansion of FFL at design.sv:50794:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50794:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50794:271
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50794:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50794:558
						mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5];
			// Trace: macro expansion of FFL at design.sv:50795:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50795:184
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50795:281
					mid_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:50795:471
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50795:568
						mid_pipe_tag_q[i + 1] <= mid_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:50796:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50796:184
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50796:281
					mid_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:50796:471
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50796:568
						mid_pipe_aux_q[i + 1] <= mid_pipe_aux_q[i];
		end
	endgenerate
	// Trace: design.sv:50799:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: design.sv:50800:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: design.sv:50801:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: design.sv:50802:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: design.sv:50803:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: design.sv:50804:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: design.sv:50805:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: design.sv:50806:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: design.sv:50807:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: design.sv:50808:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: design.sv:50809:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: design.sv:50810:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: design.sv:50815:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: design.sv:50816:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: design.sv:50817:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: design.sv:50818:3
	wire lzc_zeroes;
	// Trace: design.sv:50820:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: design.sv:50821:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: design.sv:50823:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: design.sv:50824:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: design.sv:50825:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: design.sv:50826:3
	wire sticky_after_norm;
	// Trace: design.sv:50828:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: design.sv:50830:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: design.sv:50833:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: design.sv:50842:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: design.sv:50845:3
	always @(*) begin : norm_shift_amount
		if (_sv2v_0)
			;
		// Trace: design.sv:50847:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: design.sv:50849:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: design.sv:50851:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: design.sv:50852:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: design.sv:50856:9
					norm_shamt = $unsigned(($signed(PRECISION_BITS) + 2) + exponent_product_q);
					// Trace: design.sv:50857:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: design.sv:50861:7
			norm_shamt = addend_shamt_q;
			// Trace: design.sv:50862:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: design.sv:50867:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: design.sv:50871:3
	always @(*) begin : small_norm
		if (_sv2v_0)
			;
		// Trace: design.sv:50873:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: design.sv:50874:5
		final_exponent = normalized_exponent;
		// Trace: design.sv:50877:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: design.sv:50878:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: design.sv:50879:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: design.sv:50885:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: design.sv:50886:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: design.sv:50889:7
			final_exponent = 1'sb0;
	end
	// Trace: design.sv:50894:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: design.sv:50899:3
	wire pre_round_sign;
	// Trace: design.sv:50900:3
	wire [EXP_BITS - 1:0] pre_round_exponent;
	// Trace: design.sv:50901:3
	wire [MAN_BITS - 1:0] pre_round_mantissa;
	// Trace: design.sv:50902:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] pre_round_abs;
	// Trace: design.sv:50903:3
	wire [1:0] round_sticky_bits;
	// Trace: design.sv:50905:3
	wire of_before_round;
	wire of_after_round;
	// Trace: design.sv:50906:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: design.sv:50907:3
	wire result_zero;
	// Trace: design.sv:50909:3
	wire rounded_sign;
	// Trace: design.sv:50910:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] rounded_abs;
	// Trace: design.sv:50913:3
	assign of_before_round = final_exponent >= ((2 ** EXP_BITS) - 1);
	// Trace: design.sv:50914:3
	assign uf_before_round = final_exponent == 0;
	// Trace: design.sv:50917:3
	assign pre_round_sign = final_sign_q;
	// Trace: design.sv:50918:3
	assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : $unsigned(final_exponent[EXP_BITS - 1:0]));
	// Trace: design.sv:50919:3
	assign pre_round_mantissa = (of_before_round ? {MAN_BITS {1'sb1}} : final_mantissa[MAN_BITS:1]);
	// Trace: design.sv:50920:3
	assign pre_round_abs = {pre_round_exponent, pre_round_mantissa};
	// Trace: design.sv:50923:3
	assign round_sticky_bits = (of_before_round ? 2'b11 : {final_mantissa[0], sticky_after_norm});
	// Trace: design.sv:50926:3
	fpnew_rounding #(.AbsWidth(EXP_BITS + MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: design.sv:50940:3
	assign uf_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
	// Trace: design.sv:50941:3
	assign of_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
	// Trace: design.sv:50946:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: design.sv:50947:3
	wire [4:0] regular_status;
	// Trace: design.sv:50950:3
	assign regular_result = {rounded_sign, rounded_abs};
	// Trace: design.sv:50951:3
	assign regular_status[4] = 1'b0;
	// Trace: design.sv:50952:3
	assign regular_status[3] = 1'b0;
	// Trace: design.sv:50953:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: design.sv:50954:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: design.sv:50955:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: design.sv:50958:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: design.sv:50959:3
	wire [4:0] status_d;
	// Trace: design.sv:50962:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: design.sv:50963:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: design.sv:50969:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: design.sv:50970:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: design.sv:50971:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: design.sv:50972:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: design.sv:50973:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: design.sv:50975:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: design.sv:50978:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_4232B;
	assign sv2v_tmp_4232B = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_4232B;
	// Trace: design.sv:50979:3
	wire [5:1] sv2v_tmp_07934;
	assign sv2v_tmp_07934 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_07934;
	// Trace: design.sv:50980:3
	wire [1:1] sv2v_tmp_1CCC3;
	assign sv2v_tmp_1CCC3 = mid_pipe_tag_q[NUM_MID_REGS];
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_1CCC3;
	// Trace: design.sv:50981:3
	wire [1:1] sv2v_tmp_F4A83;
	assign sv2v_tmp_F4A83 = mid_pipe_aux_q[NUM_MID_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_F4A83;
	// Trace: design.sv:50982:3
	wire [1:1] sv2v_tmp_E45E7;
	assign sv2v_tmp_E45E7 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_E45E7;
	// Trace: design.sv:50984:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: design.sv:50986:3
	genvar _gv_i_76;
	generate
		for (_gv_i_76 = 0; _gv_i_76 < NUM_OUT_REGS; _gv_i_76 = _gv_i_76 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_76;
			// Trace: design.sv:50988:5
			wire reg_ena;
			// Trace: design.sv:50992:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:50994:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:50994:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:50994:485
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:50994:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:50994:715
						out_pipe_valid_q[i + 1] <= 1'b0;
					else if (out_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:50994:867
						out_pipe_valid_q[i + 1] <= out_pipe_valid_q[i];
			// Trace: design.sv:50996:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:50998:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50998:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50998:261
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50998:451
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50998:548
						out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
			// Trace: macro expansion of FFL at design.sv:50999:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:50999:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:50999:261
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:50999:451
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:50999:548
						out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5];
			// Trace: macro expansion of FFL at design.sv:51000:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51000:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51000:271
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:51000:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51000:558
						out_pipe_tag_q[i + 1] <= out_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:51001:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51001:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51001:271
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:51001:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51001:558
						out_pipe_aux_q[i + 1] <= out_pipe_aux_q[i];
		end
	endgenerate
	// Trace: design.sv:51004:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: design.sv:51006:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: design.sv:51007:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: design.sv:51008:3
	assign extension_bit_o = 1'b1;
	// Trace: design.sv:51009:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: design.sv:51010:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: design.sv:51011:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: design.sv:51012:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
	initial _sv2v_0 = 0;
endmodule
module fpnew_fma_multi_B5D6B_A0513 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	reg _sv2v_0;
	// Trace: design.sv:51032:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: design.sv:51033:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: design.sv:51034:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: design.sv:51035:38
	// removed localparam type TagType
	// Trace: design.sv:51036:38
	// removed localparam type AuxType
	// Trace: design.sv:51038:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:34
		input reg signed [31:0] a;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:41
		input reg signed [31:0] b;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:296:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:308:48
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:309:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:5
			begin : sv2v_autoblock_1
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:312:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: design.sv:51039:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: design.sv:51041:3
	input wire clk_i;
	// Trace: design.sv:51042:3
	input wire rst_ni;
	// Trace: design.sv:51044:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: design.sv:51045:3
	input wire [14:0] is_boxed_i;
	// Trace: design.sv:51046:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:51047:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:51048:3
	input wire op_mod_i;
	// Trace: design.sv:51049:3
	input wire [2:0] src_fmt_i;
	// Trace: design.sv:51050:3
	input wire [2:0] dst_fmt_i;
	// Trace: design.sv:51051:3
	input wire tag_i;
	// Trace: design.sv:51052:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: design.sv:51054:3
	input wire in_valid_i;
	// Trace: design.sv:51055:3
	output wire in_ready_o;
	// Trace: design.sv:51056:3
	input wire flush_i;
	// Trace: design.sv:51058:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: design.sv:51059:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: design.sv:51060:3
	output wire extension_bit_o;
	// Trace: design.sv:51061:3
	output wire tag_o;
	// Trace: design.sv:51062:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: design.sv:51064:3
	output wire out_valid_o;
	// Trace: design.sv:51065:3
	input wire out_ready_i;
	// Trace: design.sv:51067:3
	output wire busy_o;
	// Trace: design.sv:51074:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:326:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:327:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:331:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:332:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:340:49
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:341:5
		reg [63:0] res;
		begin
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:342:5
			res = 1'sb0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:343:5
			begin : sv2v_autoblock_2
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:343:10
				reg [31:0] fmt;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:343:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:345:9
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt))));
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:346:9
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_5D882(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	// Trace: design.sv:51076:3
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	// Trace: design.sv:51077:3
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	// Trace: design.sv:51080:3
	localparam [31:0] PRECISION_BITS = SUPER_MAN_BITS + 1;
	// Trace: design.sv:51082:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: design.sv:51083:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: design.sv:51087:3
	localparam [31:0] EXP_WIDTH = fpnew_pkg_maximum(SUPER_EXP_BITS + 2, LZC_RESULT_WIDTH);
	// Trace: design.sv:51089:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 3);
	// Trace: design.sv:51091:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: design.sv:51096:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: design.sv:51101:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: design.sv:51110:3
	// removed localparam type fp_t
	// Trace: design.sv:51120:3
	wire [(3 * WIDTH) - 1:0] operands_q;
	// Trace: design.sv:51121:3
	wire [2:0] src_fmt_q;
	// Trace: design.sv:51122:3
	wire [2:0] dst_fmt_q;
	// Trace: design.sv:51125:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: design.sv:51126:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)) + 1) * 3) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)) + 1) * 3) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3 : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3)] inp_pipe_is_boxed_q;
	// Trace: design.sv:51127:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: design.sv:51128:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: design.sv:51129:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: design.sv:51130:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	// Trace: design.sv:51131:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: design.sv:51132:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: design.sv:51133:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: design.sv:51134:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: design.sv:51136:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: design.sv:51139:3
	wire [3 * WIDTH:1] sv2v_tmp_2F660;
	assign sv2v_tmp_2F660 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_2F660;
	// Trace: design.sv:51140:3
	wire [15:1] sv2v_tmp_F6596;
	assign sv2v_tmp_F6596 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] = sv2v_tmp_F6596;
	// Trace: design.sv:51141:3
	wire [3:1] sv2v_tmp_D6AA0;
	assign sv2v_tmp_D6AA0 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_D6AA0;
	// Trace: design.sv:51142:3
	wire [4:1] sv2v_tmp_99256;
	assign sv2v_tmp_99256 = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_99256;
	// Trace: design.sv:51143:3
	wire [1:1] sv2v_tmp_72E02;
	assign sv2v_tmp_72E02 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_72E02;
	// Trace: design.sv:51144:3
	wire [3:1] sv2v_tmp_97D9E;
	assign sv2v_tmp_97D9E = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_97D9E;
	// Trace: design.sv:51145:3
	wire [3:1] sv2v_tmp_C878E;
	assign sv2v_tmp_C878E = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_C878E;
	// Trace: design.sv:51146:3
	wire [1:1] sv2v_tmp_DE624;
	assign sv2v_tmp_DE624 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_DE624;
	// Trace: design.sv:51147:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_BFBB2;
	assign sv2v_tmp_BFBB2 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_BFBB2;
	// Trace: design.sv:51148:3
	wire [1:1] sv2v_tmp_CFC25;
	assign sv2v_tmp_CFC25 = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_CFC25;
	// Trace: design.sv:51150:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: design.sv:51152:3
	genvar _gv_i_77;
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_533F1;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_533F1 = inp;
	endfunction
	generate
		for (_gv_i_77 = 0; _gv_i_77 < NUM_INP_REGS; _gv_i_77 = _gv_i_77 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_77;
			// Trace: design.sv:51154:5
			wire reg_ena;
			// Trace: design.sv:51158:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:51160:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:51160:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:51160:485
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:51160:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:51160:715
						inp_pipe_valid_q[i + 1] <= 1'b0;
					else if (inp_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:51160:867
						inp_pipe_valid_q[i + 1] <= inp_pipe_valid_q[i];
			// Trace: design.sv:51162:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:51164:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51164:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51164:265
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51164:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51164:552
						inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3];
			// Trace: macro expansion of FFL at design.sv:51165:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51165:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51165:265
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51165:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51165:552
						inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15];
			// Trace: macro expansion of FFL at design.sv:51166:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51166:180
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51166:277
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at design.sv:51166:467
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51166:564
						inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:51167:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51167:182
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51167:279
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_4CD2E(0);
				else
					// Trace: macro expansion of FFL at design.sv:51167:469
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51167:566
						inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
			// Trace: macro expansion of FFL at design.sv:51168:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51168:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51168:265
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51168:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51168:552
						inp_pipe_op_mod_q[i + 1] <= inp_pipe_op_mod_q[i];
			// Trace: macro expansion of FFL at design.sv:51169:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51169:192
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51169:289
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_5D882(0);
				else
					// Trace: macro expansion of FFL at design.sv:51169:479
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51169:576
						inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:51170:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51170:192
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51170:289
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_5D882(0);
				else
					// Trace: macro expansion of FFL at design.sv:51170:479
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51170:576
						inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:51171:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51171:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51171:275
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:51171:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51171:562
						inp_pipe_tag_q[i + 1] <= inp_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:51172:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51172:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51172:275
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_533F1(1'sb0);
				else
					// Trace: macro expansion of FFL at design.sv:51172:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51172:562
						inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
		end
	endgenerate
	// Trace: design.sv:51175:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3];
	// Trace: design.sv:51176:3
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: design.sv:51177:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: design.sv:51182:3
	wire [14:0] fmt_sign;
	// Trace: design.sv:51183:3
	wire signed [(15 * SUPER_EXP_BITS) - 1:0] fmt_exponent;
	// Trace: design.sv:51184:3
	wire [(15 * SUPER_MAN_BITS) - 1:0] fmt_mantissa;
	// Trace: design.sv:51186:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [119:0] info_q;
	// Trace: design.sv:51189:3
	genvar _gv_fmt_5;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	function automatic signed [SUPER_EXP_BITS - 1:0] sv2v_cast_994BB_signed;
		input reg signed [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_994BB_signed = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_3FC64;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_3FC64 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_fmt_5 = 0; _gv_fmt_5 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_5 = _gv_fmt_5 + 1) begin : fmt_init_inputs
			localparam fmt = _gv_fmt_5;
			// Trace: design.sv:51191:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51192:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51193:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_5D882(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: design.sv:51196:7
				wire [(3 * FP_WIDTH) - 1:0] trimmed_ops;
				// Trace: design.sv:51199:7
				fpnew_classifier #(
					.FpFormat(sv2v_cast_5D882(fmt)),
					.NumOperands(3)
				) i_fpnew_classifier(
					.operands_i(trimmed_ops),
					.is_boxed_i(inp_pipe_is_boxed_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1))) * 3+:3]),
					.info_o(info_q[8 * (fmt * 3)+:24])
				);
				genvar _gv_op_2;
				for (_gv_op_2 = 0; _gv_op_2 < 3; _gv_op_2 = _gv_op_2 + 1) begin : gen_operands
					localparam op = _gv_op_2;
					// Trace: design.sv:51208:9
					assign trimmed_ops[op * fpnew_pkg_fp_width(sv2v_cast_5D882(_gv_fmt_5))+:fpnew_pkg_fp_width(sv2v_cast_5D882(_gv_fmt_5))] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH];
					// Trace: design.sv:51209:9
					assign fmt_sign[(fmt * 3) + op] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)];
					// Trace: design.sv:51210:9
					assign fmt_exponent[((fmt * 3) + op) * SUPER_EXP_BITS+:SUPER_EXP_BITS] = $signed({1'b0, operands_q[(op * WIDTH) + MAN_BITS+:EXP_BITS]});
					// Trace: design.sv:51211:9
					assign fmt_mantissa[((fmt * 3) + op) * SUPER_MAN_BITS+:SUPER_MAN_BITS] = {info_q[(((fmt * 3) + op) * 8) + 7], operands_q[(op * WIDTH) + (MAN_BITS - 1)-:MAN_BITS]} << (SUPER_MAN_BITS - MAN_BITS);
				end
			end
			else begin : inactive_format
				// Trace: design.sv:51215:7
				assign info_q[8 * (fmt * 3)+:24] = {3 {sv2v_cast_8(fpnew_pkg_DONT_CARE)}};
				// Trace: design.sv:51216:7
				assign fmt_sign[fmt * 3+:3] = fpnew_pkg_DONT_CARE;
				// Trace: design.sv:51217:7
				assign fmt_exponent[SUPER_EXP_BITS * (fmt * 3)+:SUPER_EXP_BITS * 3] = {3 {sv2v_cast_994BB_signed(fpnew_pkg_DONT_CARE)}};
				// Trace: design.sv:51218:7
				assign fmt_mantissa[SUPER_MAN_BITS * (fmt * 3)+:SUPER_MAN_BITS * 3] = {3 {sv2v_cast_3FC64(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	// Trace: design.sv:51222:3
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_a;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_b;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_c;
	// Trace: design.sv:51223:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: design.sv:51237:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:336:40
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:337:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_994BB;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_994BB = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_2F96C;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_2F96C = inp;
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_1FC93;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_1FC93 = inp;
	endfunction
	always @(*) begin : op_select
		if (_sv2v_0)
			;
		// Trace: design.sv:51240:5
		operand_a = {fmt_sign[src_fmt_q * 3], fmt_exponent[(src_fmt_q * 3) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[(src_fmt_q * 3) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: design.sv:51241:5
		operand_b = {fmt_sign[(src_fmt_q * 3) + 1], fmt_exponent[((src_fmt_q * 3) + 1) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((src_fmt_q * 3) + 1) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: design.sv:51242:5
		operand_c = {fmt_sign[(dst_fmt_q * 3) + 2], fmt_exponent[((dst_fmt_q * 3) + 2) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((dst_fmt_q * 3) + 2) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: design.sv:51243:5
		info_a = info_q[(src_fmt_q * 3) * 8+:8];
		// Trace: design.sv:51244:5
		info_b = info_q[((src_fmt_q * 3) + 1) * 8+:8];
		// Trace: design.sv:51245:5
		info_c = info_q[((dst_fmt_q * 3) + 2) * 8+:8];
		// Trace: design.sv:51248:5
		operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: design.sv:51250:5
		(* full_case, parallel_case *)
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_4CD2E(0):
				;
			sv2v_cast_4CD2E(1):
				// Trace: design.sv:51252:26
				operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = ~operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
			sv2v_cast_4CD2E(2): begin
				// Trace: design.sv:51254:9
				operand_a = {1'b0, sv2v_cast_994BB(fpnew_pkg_bias(src_fmt_q)), sv2v_cast_2F96C(1'sb0)};
				// Trace: design.sv:51255:9
				info_a = 8'b10000001;
			end
			sv2v_cast_4CD2E(3): begin
				// Trace: design.sv:51258:9
				operand_c = {1'b1, sv2v_cast_1FC93(1'sb0), sv2v_cast_2F96C(1'sb0)};
				// Trace: design.sv:51259:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: design.sv:51262:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_994BB(fpnew_pkg_DONT_CARE), sv2v_cast_3FC64(fpnew_pkg_DONT_CARE)};
				// Trace: design.sv:51263:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_994BB(fpnew_pkg_DONT_CARE), sv2v_cast_3FC64(fpnew_pkg_DONT_CARE)};
				// Trace: design.sv:51264:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_994BB(fpnew_pkg_DONT_CARE), sv2v_cast_3FC64(fpnew_pkg_DONT_CARE)};
				// Trace: design.sv:51265:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: design.sv:51266:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: design.sv:51267:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: design.sv:51275:3
	wire any_operand_inf;
	// Trace: design.sv:51276:3
	wire any_operand_nan;
	// Trace: design.sv:51277:3
	wire signalling_nan;
	// Trace: design.sv:51278:3
	wire effective_subtraction;
	// Trace: design.sv:51279:3
	wire tentative_sign;
	// Trace: design.sv:51282:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: design.sv:51283:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: design.sv:51284:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: design.sv:51286:3
	assign effective_subtraction = (operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))]) ^ operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	// Trace: design.sv:51288:3
	assign tentative_sign = operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	// Trace: design.sv:51293:3
	wire [WIDTH - 1:0] special_result;
	// Trace: design.sv:51294:3
	wire [4:0] special_status;
	// Trace: design.sv:51295:3
	wire result_is_special;
	// Trace: design.sv:51297:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	// Trace: design.sv:51298:3
	reg [24:0] fmt_special_status;
	// Trace: design.sv:51299:3
	reg [4:0] fmt_result_is_special;
	// Trace: design.sv:51302:3
	genvar _gv_fmt_6;
	generate
		for (_gv_fmt_6 = 0; _gv_fmt_6 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_6 = _gv_fmt_6 + 1) begin : gen_special_results
			localparam fmt = _gv_fmt_6;
			// Trace: design.sv:51304:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51305:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51306:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51308:5
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			// Trace: design.sv:51309:5
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			// Trace: design.sv:51310:5
			localparam [MAN_BITS - 1:0] ZERO_MANTISSA = 1'sb0;
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: design.sv:51313:7
				always @(*) begin : special_results
					// Trace: design.sv:51314:9
					reg [FP_WIDTH - 1:0] special_res;
					if (_sv2v_0)
						;
					// Trace: design.sv:51317:9
					special_res = {1'b0, QNAN_EXPONENT, QNAN_MANTISSA};
					// Trace: design.sv:51318:9
					fmt_special_status[fmt * 5+:5] = 1'sb0;
					// Trace: design.sv:51319:9
					fmt_result_is_special[fmt] = 1'b0;
					// Trace: design.sv:51325:9
					if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
						// Trace: design.sv:51326:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: design.sv:51327:11
						fmt_special_status[(fmt * 5) + 4] = 1'b1;
					end
					else if (any_operand_nan) begin
						// Trace: design.sv:51330:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: design.sv:51331:11
						fmt_special_status[(fmt * 5) + 4] = signalling_nan;
					end
					else if (any_operand_inf) begin
						// Trace: design.sv:51334:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: design.sv:51336:11
						if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
							// Trace: design.sv:51337:13
							fmt_special_status[(fmt * 5) + 4] = 1'b1;
						else if (info_a[4] || info_b[4])
							// Trace: design.sv:51341:13
							special_res = {operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
						else if (info_c[4])
							// Trace: design.sv:51345:13
							special_res = {operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
					end
					// Trace: design.sv:51349:9
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: design.sv:51350:9
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: design.sv:51353:7
				wire [WIDTH * 1:1] sv2v_tmp_D05EE;
				assign sv2v_tmp_D05EE = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_D05EE;
				// Trace: design.sv:51354:7
				wire [5:1] sv2v_tmp_0AFA1;
				assign sv2v_tmp_0AFA1 = 1'sb0;
				always @(*) fmt_special_status[fmt * 5+:5] = sv2v_tmp_0AFA1;
				// Trace: design.sv:51355:7
				wire [1:1] sv2v_tmp_EE036;
				assign sv2v_tmp_EE036 = 1'b0;
				always @(*) fmt_result_is_special[fmt] = sv2v_tmp_EE036;
			end
		end
	endgenerate
	// Trace: design.sv:51360:3
	assign result_is_special = fmt_result_is_special[dst_fmt_q];
	// Trace: design.sv:51362:3
	assign special_status = fmt_special_status[dst_fmt_q * 5+:5];
	// Trace: design.sv:51364:3
	assign special_result = fmt_special_result[dst_fmt_q * WIDTH+:WIDTH];
	// Trace: design.sv:51369:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: design.sv:51370:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: design.sv:51371:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: design.sv:51374:3
	assign exponent_a = $signed({1'b0, operand_a[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: design.sv:51375:3
	assign exponent_b = $signed({1'b0, operand_b[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: design.sv:51376:3
	assign exponent_c = $signed({1'b0, operand_c[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: design.sv:51380:3
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	// Trace: design.sv:51382:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(fpnew_pkg_bias(dst_fmt_q)) : $signed(((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - (2 * $signed(fpnew_pkg_bias(src_fmt_q)))) + $signed(fpnew_pkg_bias(dst_fmt_q))));
	// Trace: design.sv:51389:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: design.sv:51391:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	// Trace: design.sv:51394:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: design.sv:51396:3
	always @(*) begin : addend_shift_amount
		if (_sv2v_0)
			;
		// Trace: design.sv:51398:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: design.sv:51399:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: design.sv:51402:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: design.sv:51405:7
			addend_shamt = 0;
	end
	// Trace: design.sv:51411:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: design.sv:51412:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: design.sv:51413:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: design.sv:51416:3
	assign mantissa_a = {info_a[7], operand_a[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: design.sv:51417:3
	assign mantissa_b = {info_b[7], operand_b[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: design.sv:51418:3
	assign mantissa_c = {info_c[7], operand_c[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: design.sv:51421:3
	assign product = mantissa_a * mantissa_b;
	// Trace: design.sv:51426:3
	assign product_shifted = product << 2;
	// Trace: design.sv:51431:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: design.sv:51432:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: design.sv:51433:3
	wire sticky_before_add;
	// Trace: design.sv:51434:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: design.sv:51435:3
	wire inject_carry_in;
	// Trace: design.sv:51445:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: design.sv:51448:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: design.sv:51451:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: design.sv:51452:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: design.sv:51457:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	// Trace: design.sv:51458:3
	wire sum_carry;
	// Trace: design.sv:51459:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: design.sv:51460:3
	wire final_sign;
	// Trace: design.sv:51463:3
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: design.sv:51464:3
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	// Trace: design.sv:51467:3
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	// Trace: design.sv:51470:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: design.sv:51478:3
	wire effective_subtraction_q;
	// Trace: design.sv:51479:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: design.sv:51480:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: design.sv:51481:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: design.sv:51482:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: design.sv:51483:3
	wire sticky_before_add_q;
	// Trace: design.sv:51484:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: design.sv:51485:3
	wire final_sign_q;
	// Trace: design.sv:51486:3
	wire [2:0] dst_fmt_q2;
	// Trace: design.sv:51487:3
	wire [2:0] rnd_mode_q;
	// Trace: design.sv:51488:3
	wire result_is_special_q;
	// Trace: design.sv:51489:3
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] special_result_q;
	// Trace: design.sv:51490:3
	wire [4:0] special_status_q;
	// Trace: design.sv:51492:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: design.sv:51493:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: design.sv:51494:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: design.sv:51495:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: design.sv:51496:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: design.sv:51497:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: design.sv:51498:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: design.sv:51499:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: design.sv:51500:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: design.sv:51501:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	// Trace: design.sv:51502:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: design.sv:51503:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) + ((NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: design.sv:51504:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: design.sv:51505:3
	reg [0:NUM_MID_REGS] mid_pipe_tag_q;
	// Trace: design.sv:51506:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	// Trace: design.sv:51507:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: design.sv:51509:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: design.sv:51512:3
	wire [1:1] sv2v_tmp_301F1;
	assign sv2v_tmp_301F1 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_301F1;
	// Trace: design.sv:51513:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_C29F5;
	assign sv2v_tmp_C29F5 = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_C29F5;
	// Trace: design.sv:51514:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_24DD8;
	assign sv2v_tmp_24DD8 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_24DD8;
	// Trace: design.sv:51515:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_6091A;
	assign sv2v_tmp_6091A = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_6091A;
	// Trace: design.sv:51516:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_CB467;
	assign sv2v_tmp_CB467 = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_CB467;
	// Trace: design.sv:51517:3
	wire [1:1] sv2v_tmp_6A24C;
	assign sv2v_tmp_6A24C = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6A24C;
	// Trace: design.sv:51518:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_6ABE6;
	assign sv2v_tmp_6ABE6 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_6ABE6;
	// Trace: design.sv:51519:3
	wire [1:1] sv2v_tmp_9C379;
	assign sv2v_tmp_9C379 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_9C379;
	// Trace: design.sv:51520:3
	wire [3:1] sv2v_tmp_68647;
	assign sv2v_tmp_68647 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_68647;
	// Trace: design.sv:51521:3
	wire [3:1] sv2v_tmp_59791;
	assign sv2v_tmp_59791 = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_59791;
	// Trace: design.sv:51522:3
	wire [1:1] sv2v_tmp_08378;
	assign sv2v_tmp_08378 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_08378;
	// Trace: design.sv:51523:3
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) * 1:1] sv2v_tmp_3E0BB;
	assign sv2v_tmp_3E0BB = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] = sv2v_tmp_3E0BB;
	// Trace: design.sv:51524:3
	wire [5:1] sv2v_tmp_80D24;
	assign sv2v_tmp_80D24 = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_80D24;
	// Trace: design.sv:51525:3
	wire [1:1] sv2v_tmp_7259D;
	assign sv2v_tmp_7259D = inp_pipe_tag_q[NUM_INP_REGS];
	always @(*) mid_pipe_tag_q[0] = sv2v_tmp_7259D;
	// Trace: design.sv:51526:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_B88C1;
	assign sv2v_tmp_B88C1 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_B88C1;
	// Trace: design.sv:51527:3
	wire [1:1] sv2v_tmp_C7159;
	assign sv2v_tmp_C7159 = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_C7159;
	// Trace: design.sv:51529:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: design.sv:51532:3
	genvar _gv_i_78;
	generate
		for (_gv_i_78 = 0; _gv_i_78 < NUM_MID_REGS; _gv_i_78 = _gv_i_78 + 1) begin : gen_inside_pipeline
			localparam i = _gv_i_78;
			// Trace: design.sv:51534:5
			wire reg_ena;
			// Trace: design.sv:51538:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:51540:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:51540:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:51540:485
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:51540:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:51540:715
						mid_pipe_valid_q[i + 1] <= 1'b0;
					else if (mid_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:51540:867
						mid_pipe_valid_q[i + 1] <= mid_pipe_valid_q[i];
			// Trace: design.sv:51542:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:51544:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51544:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51544:271
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51544:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51544:558
						mid_pipe_eff_sub_q[i + 1] <= mid_pipe_eff_sub_q[i];
			// Trace: macro expansion of FFL at design.sv:51545:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51545:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51545:271
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51545:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51545:558
						mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH];
			// Trace: macro expansion of FFL at design.sv:51546:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51546:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51546:271
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51546:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51546:558
						mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH];
			// Trace: macro expansion of FFL at design.sv:51547:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51547:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51547:271
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51547:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51547:558
						mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH];
			// Trace: macro expansion of FFL at design.sv:51548:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51548:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51548:271
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51548:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51548:558
						mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
			// Trace: macro expansion of FFL at design.sv:51549:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51549:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51549:271
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51549:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51549:558
						mid_pipe_sticky_q[i + 1] <= mid_pipe_sticky_q[i];
			// Trace: macro expansion of FFL at design.sv:51550:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51550:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51550:271
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51550:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51550:558
						mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
			// Trace: macro expansion of FFL at design.sv:51551:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51551:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51551:271
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51551:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51551:558
						mid_pipe_final_sign_q[i + 1] <= mid_pipe_final_sign_q[i];
			// Trace: macro expansion of FFL at design.sv:51552:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51552:186
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51552:283
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at design.sv:51552:473
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51552:570
						mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:51553:101
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51553:198
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51553:295
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_5D882(0);
				else
					// Trace: macro expansion of FFL at design.sv:51553:485
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51553:582
						mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
			// Trace: macro expansion of FFL at design.sv:51554:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51554:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51554:271
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51554:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51554:558
						mid_pipe_res_is_spec_q[i + 1] <= mid_pipe_res_is_spec_q[i];
			// Trace: macro expansion of FFL at design.sv:51555:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51555:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51555:271
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51555:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51555:558
						mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS];
			// Trace: macro expansion of FFL at design.sv:51556:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51556:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51556:271
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51556:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51556:558
						mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5];
			// Trace: macro expansion of FFL at design.sv:51557:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51557:184
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51557:281
					mid_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:51557:471
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51557:568
						mid_pipe_tag_q[i + 1] <= mid_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:51558:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51558:184
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51558:281
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_533F1(1'sb0);
				else
					// Trace: macro expansion of FFL at design.sv:51558:471
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51558:568
						mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
		end
	endgenerate
	// Trace: design.sv:51561:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: design.sv:51562:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: design.sv:51563:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: design.sv:51564:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: design.sv:51565:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: design.sv:51566:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: design.sv:51567:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: design.sv:51568:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: design.sv:51569:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: design.sv:51570:3
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: design.sv:51571:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: design.sv:51572:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS];
	// Trace: design.sv:51573:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: design.sv:51578:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: design.sv:51579:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: design.sv:51580:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: design.sv:51581:3
	wire lzc_zeroes;
	// Trace: design.sv:51583:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: design.sv:51584:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: design.sv:51586:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: design.sv:51587:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: design.sv:51588:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: design.sv:51589:3
	wire sticky_after_norm;
	// Trace: design.sv:51591:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: design.sv:51593:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: design.sv:51596:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: design.sv:51605:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: design.sv:51608:3
	always @(*) begin : norm_shift_amount
		if (_sv2v_0)
			;
		// Trace: design.sv:51610:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: design.sv:51612:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: design.sv:51614:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: design.sv:51615:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: design.sv:51619:9
					norm_shamt = $unsigned($signed((PRECISION_BITS + 2) + exponent_product_q));
					// Trace: design.sv:51620:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: design.sv:51624:7
			norm_shamt = addend_shamt_q;
			// Trace: design.sv:51625:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: design.sv:51630:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: design.sv:51634:3
	always @(*) begin : small_norm
		if (_sv2v_0)
			;
		// Trace: design.sv:51636:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: design.sv:51637:5
		final_exponent = normalized_exponent;
		// Trace: design.sv:51640:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: design.sv:51641:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: design.sv:51642:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: design.sv:51648:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: design.sv:51649:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: design.sv:51652:7
			final_exponent = 1'sb0;
	end
	// Trace: design.sv:51657:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: design.sv:51662:3
	wire pre_round_sign;
	// Trace: design.sv:51663:3
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] pre_round_abs;
	// Trace: design.sv:51664:3
	wire [1:0] round_sticky_bits;
	// Trace: design.sv:51666:3
	wire of_before_round;
	wire of_after_round;
	// Trace: design.sv:51667:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: design.sv:51669:3
	wire [(NUM_FORMATS * (SUPER_EXP_BITS + SUPER_MAN_BITS)) - 1:0] fmt_pre_round_abs;
	// Trace: design.sv:51670:3
	wire [9:0] fmt_round_sticky_bits;
	// Trace: design.sv:51672:3
	reg [4:0] fmt_of_after_round;
	// Trace: design.sv:51673:3
	reg [4:0] fmt_uf_after_round;
	// Trace: design.sv:51675:3
	wire rounded_sign;
	// Trace: design.sv:51676:3
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] rounded_abs;
	// Trace: design.sv:51677:3
	wire result_zero;
	// Trace: design.sv:51680:3
	assign of_before_round = final_exponent >= ((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1);
	// Trace: design.sv:51681:3
	assign uf_before_round = final_exponent == 0;
	// Trace: design.sv:51684:3
	genvar _gv_fmt_7;
	generate
		for (_gv_fmt_7 = 0; _gv_fmt_7 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_7 = _gv_fmt_7 + 1) begin : gen_res_assemble
			localparam fmt = _gv_fmt_7;
			// Trace: design.sv:51686:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51687:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51689:5
			wire [EXP_BITS - 1:0] pre_round_exponent;
			// Trace: design.sv:51690:5
			wire [MAN_BITS - 1:0] pre_round_mantissa;
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: design.sv:51694:7
				assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : final_exponent[EXP_BITS - 1:0]);
				// Trace: design.sv:51695:7
				assign pre_round_mantissa = (of_before_round ? {fpnew_pkg_man_bits(sv2v_cast_5D882(_gv_fmt_7)) {1'sb1}} : final_mantissa[SUPER_MAN_BITS-:MAN_BITS]);
				// Trace: design.sv:51697:7
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {pre_round_exponent, pre_round_mantissa};
				// Trace: design.sv:51700:7
				assign fmt_round_sticky_bits[(fmt * 2) + 1] = final_mantissa[SUPER_MAN_BITS - MAN_BITS] | of_before_round;
				if (MAN_BITS < SUPER_MAN_BITS) begin : narrow_sticky
					// Trace: design.sv:51705:9
					assign fmt_round_sticky_bits[fmt * 2] = (|final_mantissa[(SUPER_MAN_BITS - MAN_BITS) - 1:0] | sticky_after_norm) | of_before_round;
				end
				else begin : normal_sticky
					// Trace: design.sv:51708:9
					assign fmt_round_sticky_bits[fmt * 2] = sticky_after_norm | of_before_round;
				end
			end
			else begin : inactive_format
				// Trace: design.sv:51711:7
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {SUPER_EXP_BITS + SUPER_MAN_BITS {fpnew_pkg_DONT_CARE}};
				// Trace: design.sv:51712:7
				assign fmt_round_sticky_bits[fmt * 2+:2] = {2 {fpnew_pkg_DONT_CARE}};
			end
		end
	endgenerate
	// Trace: design.sv:51717:3
	assign pre_round_sign = final_sign_q;
	// Trace: design.sv:51718:3
	assign pre_round_abs = fmt_pre_round_abs[dst_fmt_q2 * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS];
	// Trace: design.sv:51721:3
	assign round_sticky_bits = fmt_round_sticky_bits[dst_fmt_q2 * 2+:2];
	// Trace: design.sv:51724:3
	fpnew_rounding #(.AbsWidth(SUPER_EXP_BITS + SUPER_MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: design.sv:51737:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	// Trace: design.sv:51739:3
	genvar _gv_fmt_8;
	generate
		for (_gv_fmt_8 = 0; _gv_fmt_8 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_8 = _gv_fmt_8 + 1) begin : gen_sign_inject
			localparam fmt = _gv_fmt_8;
			// Trace: design.sv:51741:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51742:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_5D882(fmt));
			// Trace: design.sv:51743:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_5D882(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: design.sv:51746:7
				always @(*) begin : post_process
					if (_sv2v_0)
						;
					// Trace: design.sv:51748:9
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					// Trace: design.sv:51749:9
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					// Trace: design.sv:51752:9
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: design.sv:51753:9
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]};
				end
			end
			else begin : inactive_format
				// Trace: design.sv:51756:7
				wire [1:1] sv2v_tmp_4C394;
				assign sv2v_tmp_4C394 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4C394;
				// Trace: design.sv:51757:7
				wire [1:1] sv2v_tmp_5852E;
				assign sv2v_tmp_5852E = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_5852E;
				// Trace: design.sv:51758:7
				wire [WIDTH * 1:1] sv2v_tmp_49668;
				assign sv2v_tmp_49668 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_49668;
			end
		end
	endgenerate
	// Trace: design.sv:51763:3
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	// Trace: design.sv:51764:3
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	// Trace: design.sv:51770:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: design.sv:51771:3
	wire [4:0] regular_status;
	// Trace: design.sv:51774:3
	assign regular_result = fmt_result[dst_fmt_q2 * WIDTH+:WIDTH];
	// Trace: design.sv:51775:3
	assign regular_status[4] = 1'b0;
	// Trace: design.sv:51776:3
	assign regular_status[3] = 1'b0;
	// Trace: design.sv:51777:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: design.sv:51778:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: design.sv:51779:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: design.sv:51782:3
	wire [WIDTH - 1:0] result_d;
	// Trace: design.sv:51783:3
	wire [4:0] status_d;
	// Trace: design.sv:51786:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: design.sv:51787:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: design.sv:51793:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: design.sv:51794:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: design.sv:51795:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: design.sv:51796:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: design.sv:51797:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: design.sv:51799:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: design.sv:51802:3
	wire [WIDTH * 1:1] sv2v_tmp_469C2;
	assign sv2v_tmp_469C2 = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_469C2;
	// Trace: design.sv:51803:3
	wire [5:1] sv2v_tmp_A6238;
	assign sv2v_tmp_A6238 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_A6238;
	// Trace: design.sv:51804:3
	wire [1:1] sv2v_tmp_1CCC3;
	assign sv2v_tmp_1CCC3 = mid_pipe_tag_q[NUM_MID_REGS];
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_1CCC3;
	// Trace: design.sv:51805:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_D2D68;
	assign sv2v_tmp_D2D68 = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_D2D68;
	// Trace: design.sv:51806:3
	wire [1:1] sv2v_tmp_E45E7;
	assign sv2v_tmp_E45E7 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_E45E7;
	// Trace: design.sv:51808:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: design.sv:51810:3
	genvar _gv_i_79;
	generate
		for (_gv_i_79 = 0; _gv_i_79 < NUM_OUT_REGS; _gv_i_79 = _gv_i_79 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_79;
			// Trace: design.sv:51812:5
			wire reg_ena;
			// Trace: design.sv:51816:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:51818:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:51818:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:51818:485
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:51818:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:51818:715
						out_pipe_valid_q[i + 1] <= 1'b0;
					else if (out_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:51818:867
						out_pipe_valid_q[i + 1] <= out_pipe_valid_q[i];
			// Trace: design.sv:51820:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:51822:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51822:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51822:261
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51822:451
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51822:548
						out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH];
			// Trace: macro expansion of FFL at design.sv:51823:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51823:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51823:261
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51823:451
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51823:548
						out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5];
			// Trace: macro expansion of FFL at design.sv:51824:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51824:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51824:271
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:51824:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51824:558
						out_pipe_tag_q[i + 1] <= out_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:51825:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51825:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51825:271
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_533F1(1'sb0);
				else
					// Trace: macro expansion of FFL at design.sv:51825:461
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51825:558
						out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
		end
	endgenerate
	// Trace: design.sv:51828:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: design.sv:51830:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: design.sv:51831:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: design.sv:51832:3
	assign extension_bit_o = 1'b1;
	// Trace: design.sv:51833:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: design.sv:51834:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: design.sv:51835:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: design.sv:51836:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
	initial _sv2v_0 = 0;
endmodule
module fpnew_noncomp_DE16F (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	class_mask_o,
	is_class_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	reg _sv2v_0;
	// Trace: design.sv:51856:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_5D882(0);
	// Trace: design.sv:51857:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: design.sv:51858:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: design.sv:51859:38
	// removed localparam type TagType
	// Trace: design.sv:51860:38
	// removed localparam type AuxType
	// Trace: design.sv:51862:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: design.sv:51864:3
	input wire clk_i;
	// Trace: design.sv:51865:3
	input wire rst_ni;
	// Trace: design.sv:51867:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: design.sv:51868:3
	input wire [1:0] is_boxed_i;
	// Trace: design.sv:51869:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:51870:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:51871:3
	input wire op_mod_i;
	// Trace: design.sv:51872:3
	input wire tag_i;
	// Trace: design.sv:51873:3
	input wire aux_i;
	// Trace: design.sv:51875:3
	input wire in_valid_i;
	// Trace: design.sv:51876:3
	output wire in_ready_o;
	// Trace: design.sv:51877:3
	input wire flush_i;
	// Trace: design.sv:51879:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: design.sv:51880:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: design.sv:51881:3
	output wire extension_bit_o;
	// Trace: design.sv:51882:3
	// removed localparam type fpnew_pkg_classmask_e
	output wire [9:0] class_mask_o;
	// Trace: design.sv:51883:3
	output wire is_class_o;
	// Trace: design.sv:51884:3
	output wire tag_o;
	// Trace: design.sv:51885:3
	output wire aux_o;
	// Trace: design.sv:51887:3
	output wire out_valid_o;
	// Trace: design.sv:51888:3
	input wire out_ready_i;
	// Trace: design.sv:51890:3
	output wire busy_o;
	// Trace: design.sv:51896:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:326:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:327:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: design.sv:51897:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:331:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:332:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: design.sv:51899:3
	localparam NUM_INP_REGS = ((PipeConfig == 2'd0) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: design.sv:51904:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: design.sv:51913:3
	// removed localparam type fp_t
	// Trace: design.sv:51923:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: design.sv:51924:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)] inp_pipe_is_boxed_q;
	// Trace: design.sv:51925:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: design.sv:51926:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: design.sv:51927:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: design.sv:51928:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: design.sv:51929:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: design.sv:51930:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: design.sv:51932:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: design.sv:51935:3
	wire [2 * WIDTH:1] sv2v_tmp_E768C;
	assign sv2v_tmp_E768C = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_E768C;
	// Trace: design.sv:51936:3
	wire [2:1] sv2v_tmp_9866C;
	assign sv2v_tmp_9866C = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2+:2] = sv2v_tmp_9866C;
	// Trace: design.sv:51937:3
	wire [3:1] sv2v_tmp_B26FC;
	assign sv2v_tmp_B26FC = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_B26FC;
	// Trace: design.sv:51938:3
	wire [4:1] sv2v_tmp_6E66E;
	assign sv2v_tmp_6E66E = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_6E66E;
	// Trace: design.sv:51939:3
	wire [1:1] sv2v_tmp_72E02;
	assign sv2v_tmp_72E02 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_72E02;
	// Trace: design.sv:51940:3
	wire [1:1] sv2v_tmp_DE624;
	assign sv2v_tmp_DE624 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_DE624;
	// Trace: design.sv:51941:3
	wire [1:1] sv2v_tmp_683C4;
	assign sv2v_tmp_683C4 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_683C4;
	// Trace: design.sv:51942:3
	wire [1:1] sv2v_tmp_CFC25;
	assign sv2v_tmp_CFC25 = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_CFC25;
	// Trace: design.sv:51944:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: design.sv:51946:3
	genvar _gv_i_80;
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	generate
		for (_gv_i_80 = 0; _gv_i_80 < NUM_INP_REGS; _gv_i_80 = _gv_i_80 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_80;
			// Trace: design.sv:51948:5
			wire reg_ena;
			// Trace: design.sv:51952:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:51954:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:51954:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:51954:485
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:51954:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:51954:715
						inp_pipe_valid_q[i + 1] <= 1'b0;
					else if (inp_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:51954:867
						inp_pipe_valid_q[i + 1] <= inp_pipe_valid_q[i];
			// Trace: design.sv:51956:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:51958:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51958:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51958:265
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51958:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51958:552
						inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2];
			// Trace: macro expansion of FFL at design.sv:51959:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51959:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51959:265
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51959:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51959:552
						inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2+:2];
			// Trace: macro expansion of FFL at design.sv:51960:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51960:180
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51960:277
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at design.sv:51960:467
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51960:564
						inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3];
			// Trace: macro expansion of FFL at design.sv:51961:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51961:182
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51961:279
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_4CD2E(0);
				else
					// Trace: macro expansion of FFL at design.sv:51961:469
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51961:566
						inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
			// Trace: macro expansion of FFL at design.sv:51962:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51962:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51962:265
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:51962:455
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51962:552
						inp_pipe_op_mod_q[i + 1] <= inp_pipe_op_mod_q[i];
			// Trace: macro expansion of FFL at design.sv:51963:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51963:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51963:275
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:51963:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51963:562
						inp_pipe_tag_q[i + 1] <= inp_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:51964:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:51964:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:51964:275
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:51964:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:51964:562
						inp_pipe_aux_q[i + 1] <= inp_pipe_aux_q[i];
		end
	endgenerate
	// Trace: design.sv:51970:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [15:0] info_q;
	// Trace: design.sv:51973:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(2)
	) i_class_a(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2+:2]),
		.info_o(info_q)
	);
	// Trace: design.sv:51982:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	// Trace: design.sv:51983:3
	wire [7:0] info_a;
	wire [7:0] info_b;
	// Trace: design.sv:51986:3
	assign operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	// Trace: design.sv:51987:3
	assign operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	// Trace: design.sv:51988:3
	assign info_a = info_q[0+:8];
	// Trace: design.sv:51989:3
	assign info_b = info_q[8+:8];
	// Trace: design.sv:51991:3
	wire any_operand_inf;
	// Trace: design.sv:51992:3
	wire any_operand_nan;
	// Trace: design.sv:51993:3
	wire signalling_nan;
	// Trace: design.sv:51996:3
	assign any_operand_inf = |{info_a[4], info_b[4]};
	// Trace: design.sv:51997:3
	assign any_operand_nan = |{info_a[3], info_b[3]};
	// Trace: design.sv:51998:3
	assign signalling_nan = |{info_a[2], info_b[2]};
	// Trace: design.sv:52000:3
	wire operands_equal;
	wire operand_a_smaller;
	// Trace: design.sv:52003:3
	assign operands_equal = (operand_a == operand_b) || (info_a[5] && info_b[5]);
	// Trace: design.sv:52005:3
	assign operand_a_smaller = (operand_a < operand_b) ^ (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] || operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]);
	// Trace: design.sv:52010:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] sgnj_result;
	// Trace: design.sv:52011:3
	wire [4:0] sgnj_status;
	// Trace: design.sv:52012:3
	wire sgnj_extension_bit;
	// Trace: design.sv:52016:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_8D8F7;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_8D8F7 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_D5F4C;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_D5F4C = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_51E93;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_51E93 = inp;
	endfunction
	always @(*) begin : sign_injections
		// Trace: design.sv:52017:5
		reg sign_a;
		reg sign_b;
		if (_sv2v_0)
			;
		// Trace: design.sv:52019:5
		sgnj_result = operand_a;
		// Trace: design.sv:52022:5
		if (!info_a[0])
			// Trace: design.sv:52022:27
			sgnj_result = {1'b0, sv2v_cast_8D8F7(1'sb1), sv2v_cast_D5F4C(2 ** (MAN_BITS - 1))};
		// Trace: design.sv:52025:5
		sign_a = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] & info_a[0];
		// Trace: design.sv:52026:5
		sign_b = operand_b[1 + (EXP_BITS + (MAN_BITS - 1))] & info_b[0];
		(* full_case, parallel_case *)
		case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
			3'b000:
				// Trace: design.sv:52030:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_b;
			3'b001:
				// Trace: design.sv:52031:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = ~sign_b;
			3'b010:
				// Trace: design.sv:52032:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_a ^ sign_b;
			3'b011:
				// Trace: design.sv:52033:23
				sgnj_result = operand_a;
			default:
				// Trace: design.sv:52034:16
				sgnj_result = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
		endcase
	end
	// Trace: design.sv:52038:3
	assign sgnj_status = 1'sb0;
	// Trace: design.sv:52041:3
	assign sgnj_extension_bit = (inp_pipe_op_mod_q[NUM_INP_REGS] ? sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] : 1'b1);
	// Trace: design.sv:52046:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] minmax_result;
	// Trace: design.sv:52047:3
	reg [4:0] minmax_status;
	// Trace: design.sv:52048:3
	wire minmax_extension_bit;
	// Trace: design.sv:52052:3
	always @(*) begin : min_max
		if (_sv2v_0)
			;
		// Trace: design.sv:52054:5
		minmax_status = 1'sb0;
		// Trace: design.sv:52057:5
		minmax_status[4] = signalling_nan;
		// Trace: design.sv:52060:5
		if (info_a[3] && info_b[3])
			// Trace: design.sv:52061:7
			minmax_result = {1'b0, sv2v_cast_8D8F7(1'sb1), sv2v_cast_D5F4C(2 ** (MAN_BITS - 1))};
		else if (info_a[3])
			// Trace: design.sv:52063:29
			minmax_result = operand_b;
		else if (info_b[3])
			// Trace: design.sv:52064:29
			minmax_result = operand_a;
		else
			// Trace: design.sv:52067:7
			(* full_case, parallel_case *)
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					// Trace: design.sv:52068:25
					minmax_result = (operand_a_smaller ? operand_a : operand_b);
				3'b001:
					// Trace: design.sv:52069:25
					minmax_result = (operand_a_smaller ? operand_b : operand_a);
				default:
					// Trace: design.sv:52070:18
					minmax_result = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
			endcase
	end
	// Trace: design.sv:52075:3
	assign minmax_extension_bit = 1'b1;
	// Trace: design.sv:52080:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] cmp_result;
	// Trace: design.sv:52081:3
	reg [4:0] cmp_status;
	// Trace: design.sv:52082:3
	wire cmp_extension_bit;
	// Trace: design.sv:52087:3
	always @(*) begin : comparisons
		if (_sv2v_0)
			;
		// Trace: design.sv:52089:5
		cmp_result = 1'sb0;
		// Trace: design.sv:52090:5
		cmp_status = 1'sb0;
		// Trace: design.sv:52093:5
		if (signalling_nan)
			// Trace: design.sv:52093:25
			cmp_status[4] = 1'b1;
		else
			// Trace: design.sv:52096:7
			(* full_case, parallel_case *)
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					// Trace: design.sv:52098:11
					if (any_operand_nan)
						// Trace: design.sv:52098:32
						cmp_status[4] = 1'b1;
					else
						// Trace: design.sv:52099:16
						cmp_result = (operand_a_smaller | operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b001:
					// Trace: design.sv:52102:11
					if (any_operand_nan)
						// Trace: design.sv:52102:32
						cmp_status[4] = 1'b1;
					else
						// Trace: design.sv:52103:16
						cmp_result = (operand_a_smaller & ~operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b010:
					// Trace: design.sv:52106:11
					if (any_operand_nan)
						// Trace: design.sv:52106:32
						cmp_result = inp_pipe_op_mod_q[NUM_INP_REGS];
					else
						// Trace: design.sv:52107:16
						cmp_result = operands_equal ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				default:
					// Trace: design.sv:52109:18
					cmp_result = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
			endcase
	end
	// Trace: design.sv:52114:3
	assign cmp_extension_bit = 1'b0;
	// Trace: design.sv:52119:3
	wire [4:0] class_status;
	// Trace: design.sv:52120:3
	wire class_extension_bit;
	// Trace: design.sv:52121:3
	reg [9:0] class_mask_d;
	// Trace: design.sv:52124:3
	always @(*) begin : classify
		if (_sv2v_0)
			;
		// Trace: design.sv:52125:5
		if (info_a[7])
			// Trace: design.sv:52126:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000010 : 10'b0001000000);
		else if (info_a[6])
			// Trace: design.sv:52128:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000100 : 10'b0000100000);
		else if (info_a[5])
			// Trace: design.sv:52130:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000001000 : 10'b0000010000);
		else if (info_a[4])
			// Trace: design.sv:52132:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000001 : 10'b0010000000);
		else if (info_a[3])
			// Trace: design.sv:52134:7
			class_mask_d = (info_a[2] ? 10'b0100000000 : 10'b1000000000);
		else
			// Trace: design.sv:52136:7
			class_mask_d = 10'b1000000000;
	end
	// Trace: design.sv:52140:3
	assign class_status = 1'sb0;
	// Trace: design.sv:52141:3
	assign class_extension_bit = 1'b0;
	// Trace: design.sv:52146:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: design.sv:52147:3
	reg [4:0] status_d;
	// Trace: design.sv:52148:3
	reg extension_bit_d;
	// Trace: design.sv:52149:3
	wire is_class_d;
	// Trace: design.sv:52152:3
	always @(*) begin : select_result
		if (_sv2v_0)
			;
		// Trace: design.sv:52153:5
		(* full_case, parallel_case *)
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_4CD2E(6): begin
				// Trace: design.sv:52155:9
				result_d = sgnj_result;
				// Trace: design.sv:52156:9
				status_d = sgnj_status;
				// Trace: design.sv:52157:9
				extension_bit_d = sgnj_extension_bit;
			end
			sv2v_cast_4CD2E(7): begin
				// Trace: design.sv:52160:9
				result_d = minmax_result;
				// Trace: design.sv:52161:9
				status_d = minmax_status;
				// Trace: design.sv:52162:9
				extension_bit_d = minmax_extension_bit;
			end
			sv2v_cast_4CD2E(8): begin
				// Trace: design.sv:52165:9
				result_d = cmp_result;
				// Trace: design.sv:52166:9
				status_d = cmp_status;
				// Trace: design.sv:52167:9
				extension_bit_d = cmp_extension_bit;
			end
			sv2v_cast_4CD2E(9): begin
				// Trace: design.sv:52170:9
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
				// Trace: design.sv:52171:9
				status_d = class_status;
				// Trace: design.sv:52172:9
				extension_bit_d = class_extension_bit;
			end
			default: begin
				// Trace: design.sv:52175:9
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
				// Trace: design.sv:52176:9
				status_d = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: design.sv:52177:9
				extension_bit_d = fpnew_pkg_DONT_CARE;
			end
		endcase
	end
	// Trace: design.sv:52182:3
	assign is_class_d = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_4CD2E(9);
	// Trace: design.sv:52188:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: design.sv:52189:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: design.sv:52190:3
	reg [0:NUM_OUT_REGS] out_pipe_extension_bit_q;
	// Trace: design.sv:52191:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 10) + ((NUM_OUT_REGS * 10) - 1) : ((NUM_OUT_REGS + 1) * 10) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 10 : 0)] out_pipe_class_mask_q;
	// Trace: design.sv:52192:3
	reg [0:NUM_OUT_REGS] out_pipe_is_class_q;
	// Trace: design.sv:52193:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: design.sv:52194:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: design.sv:52195:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: design.sv:52197:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: design.sv:52200:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_35063;
	assign sv2v_tmp_35063 = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_35063;
	// Trace: design.sv:52201:3
	wire [5:1] sv2v_tmp_036FC;
	assign sv2v_tmp_036FC = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_036FC;
	// Trace: design.sv:52202:3
	wire [1:1] sv2v_tmp_C9204;
	assign sv2v_tmp_C9204 = extension_bit_d;
	always @(*) out_pipe_extension_bit_q[0] = sv2v_tmp_C9204;
	// Trace: design.sv:52203:3
	wire [10:1] sv2v_tmp_0A406;
	assign sv2v_tmp_0A406 = class_mask_d;
	always @(*) out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 10+:10] = sv2v_tmp_0A406;
	// Trace: design.sv:52204:3
	wire [1:1] sv2v_tmp_C899A;
	assign sv2v_tmp_C899A = is_class_d;
	always @(*) out_pipe_is_class_q[0] = sv2v_tmp_C899A;
	// Trace: design.sv:52205:3
	wire [1:1] sv2v_tmp_13053;
	assign sv2v_tmp_13053 = inp_pipe_tag_q[NUM_INP_REGS];
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_13053;
	// Trace: design.sv:52206:3
	wire [1:1] sv2v_tmp_571F3;
	assign sv2v_tmp_571F3 = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_571F3;
	// Trace: design.sv:52207:3
	wire [1:1] sv2v_tmp_B2A17;
	assign sv2v_tmp_B2A17 = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_B2A17;
	// Trace: design.sv:52209:3
	assign inp_pipe_ready[NUM_INP_REGS] = out_pipe_ready[0];
	// Trace: design.sv:52211:3
	genvar _gv_i_81;
	generate
		for (_gv_i_81 = 0; _gv_i_81 < NUM_OUT_REGS; _gv_i_81 = _gv_i_81 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_81;
			// Trace: design.sv:52213:5
			wire reg_ena;
			// Trace: design.sv:52217:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at design.sv:52219:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at design.sv:52219:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:52219:485
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at design.sv:52219:637
					if (flush_i)
						// Trace: macro expansion of FFLARNC at design.sv:52219:715
						out_pipe_valid_q[i + 1] <= 1'b0;
					else if (out_pipe_ready[i])
						// Trace: macro expansion of FFLARNC at design.sv:52219:867
						out_pipe_valid_q[i + 1] <= out_pipe_valid_q[i];
			// Trace: design.sv:52221:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at design.sv:52223:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:52223:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:52223:275
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:52223:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:52223:562
						out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
			// Trace: macro expansion of FFL at design.sv:52224:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:52224:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:52224:275
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:52224:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:52224:562
						out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5];
			// Trace: macro expansion of FFL at design.sv:52225:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:52225:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:52225:275
					out_pipe_extension_bit_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:52225:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:52225:562
						out_pipe_extension_bit_q[i + 1] <= out_pipe_extension_bit_q[i];
			// Trace: macro expansion of FFL at design.sv:52226:94
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:52226:191
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:52226:288
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= 10'b1000000000;
				else
					// Trace: macro expansion of FFL at design.sv:52226:478
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:52226:575
						out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 10+:10];
			// Trace: macro expansion of FFL at design.sv:52227:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:52227:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:52227:275
					out_pipe_is_class_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at design.sv:52227:465
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:52227:562
						out_pipe_is_class_q[i + 1] <= out_pipe_is_class_q[i];
			// Trace: macro expansion of FFL at design.sv:52228:91
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:52228:188
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:52228:285
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:52228:475
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:52228:572
						out_pipe_tag_q[i + 1] <= out_pipe_tag_q[i];
			// Trace: macro expansion of FFL at design.sv:52229:91
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at design.sv:52229:188
				if (!rst_ni)
					// Trace: macro expansion of FFL at design.sv:52229:285
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at design.sv:52229:475
					if (reg_ena)
						// Trace: macro expansion of FFL at design.sv:52229:572
						out_pipe_aux_q[i + 1] <= out_pipe_aux_q[i];
		end
	endgenerate
	// Trace: design.sv:52232:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: design.sv:52234:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: design.sv:52235:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: design.sv:52236:3
	assign extension_bit_o = out_pipe_extension_bit_q[NUM_OUT_REGS];
	// Trace: design.sv:52237:3
	assign class_mask_o = out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 10+:10];
	// Trace: design.sv:52238:3
	assign is_class_o = out_pipe_is_class_q[NUM_OUT_REGS];
	// Trace: design.sv:52239:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: design.sv:52240:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: design.sv:52241:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: design.sv:52242:3
	assign busy_o = |{inp_pipe_valid_q, out_pipe_valid_q};
	initial _sv2v_0 = 0;
endmodule
module fpnew_opgroup_block_37AAD (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// Trace: design.sv:52260:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: design.sv:52262:13
	parameter [31:0] Width = 32;
	// Trace: design.sv:52263:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: design.sv:52264:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtMask = 1'sb1;
	// Trace: design.sv:52265:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtMask = 1'sb1;
	// Trace: design.sv:52266:13
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	parameter [159:0] FmtPipeRegs = {fpnew_pkg_NUM_FP_FORMATS {32'd0}};
	// Trace: design.sv:52267:13
	// removed localparam type fpnew_pkg_unit_type_t
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	parameter [9:0] FmtUnitTypes = {fpnew_pkg_NUM_FP_FORMATS {2'd1}};
	// Trace: design.sv:52268:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: design.sv:52269:41
	// removed localparam type TagType
	// Trace: design.sv:52271:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: design.sv:52272:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:378:48
		input reg [1:0] grp;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:379:5
		(* full_case, parallel_case *)
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: design.sv:52274:3
	input wire clk_i;
	// Trace: design.sv:52275:3
	input wire rst_ni;
	// Trace: design.sv:52277:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: design.sv:52278:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: design.sv:52279:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:52280:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:52281:3
	input wire op_mod_i;
	// Trace: design.sv:52282:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: design.sv:52283:3
	input wire [2:0] dst_fmt_i;
	// Trace: design.sv:52284:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: design.sv:52285:3
	input wire vectorial_op_i;
	// Trace: design.sv:52286:3
	input wire tag_i;
	// Trace: design.sv:52288:3
	input wire in_valid_i;
	// Trace: design.sv:52289:3
	output wire in_ready_o;
	// Trace: design.sv:52290:3
	input wire flush_i;
	// Trace: design.sv:52292:3
	output wire [Width - 1:0] result_o;
	// Trace: design.sv:52293:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: design.sv:52294:3
	output wire extension_bit_o;
	// Trace: design.sv:52295:3
	output wire tag_o;
	// Trace: design.sv:52297:3
	output wire out_valid_o;
	// Trace: design.sv:52298:3
	input wire out_ready_i;
	// Trace: design.sv:52300:3
	output wire busy_o;
	// Trace: design.sv:52306:3
	// removed localparam type output_t
	// Trace: design.sv:52314:3
	wire [4:0] fmt_in_ready;
	wire [4:0] fmt_out_valid;
	wire [4:0] fmt_out_ready;
	wire [4:0] fmt_busy;
	// Trace: design.sv:52315:3
	wire [((Width + 6) >= 0 ? (5 * (Width + 7)) - 1 : (5 * (1 - (Width + 6))) + (Width + 5)):((Width + 6) >= 0 ? 0 : Width + 6)] fmt_outputs;
	// Trace: design.sv:52320:3
	assign in_ready_o = in_valid_i & fmt_in_ready[dst_fmt_i];
	// Trace: design.sv:52325:3
	genvar _gv_fmt_9;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic fpnew_pkg_any_enabled_multi;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:458:46
		input reg [9:0] types;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:458:70
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:459:5
			begin : sv2v_autoblock_1
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:459:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:459:10
				begin : sv2v_autoblock_2
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_any_enabled_multi = 1'b1;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_any_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	function automatic [2:0] fpnew_pkg_get_first_enabled_multi;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:476:58
		input reg [9:0] types;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:476:82
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:477:5
			begin : sv2v_autoblock_3
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:477:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:477:10
				begin : sv2v_autoblock_4
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_get_first_enabled_multi = sv2v_cast_5D882(i);
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_get_first_enabled_multi = sv2v_cast_5D882(0);
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic fpnew_pkg_is_first_enabled_multi;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:466:51
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:467:51
		input reg [9:0] types;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:468:51
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:469:5
			begin : sv2v_autoblock_5
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:469:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:469:10
				begin : sv2v_autoblock_6
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:470:7
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_is_first_enabled_multi = sv2v_cast_5D882(i) == fmt;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_is_first_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_fmt_9 = 0; _gv_fmt_9 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_9 = _gv_fmt_9 + 1) begin : gen_parallel_slices
			localparam fmt = _gv_fmt_9;
			// Trace: design.sv:52327:5
			localparam [0:0] ANY_MERGED = fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: design.sv:52328:5
			localparam [0:0] IS_FIRST_MERGED = fpnew_pkg_is_first_enabled_multi(sv2v_cast_5D882(fmt), FmtUnitTypes, FpFmtMask);
			if (FpFmtMask[fmt] && (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd1)) begin : active_format
				// Trace: design.sv:52334:7
				wire in_valid;
				// Trace: design.sv:52336:7
				assign in_valid = in_valid_i & (dst_fmt_i == fmt);
				// Trace: design.sv:52338:7
				fpnew_opgroup_fmt_slice_07650 #(
					.OpGroup(OpGroup),
					.FpFormat(sv2v_cast_5D882(fmt)),
					.Width(Width),
					.EnableVectors(EnableVectors),
					.NumPipeRegs(FmtPipeRegs[(4 - fmt) * 32+:32]),
					.PipeConfig(PipeConfig)
				) i_fmt_slice(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.operands_i(operands_i),
					.is_boxed_i(is_boxed_i[fmt * NUM_OPERANDS+:NUM_OPERANDS]),
					.rnd_mode_i(rnd_mode_i),
					.op_i(op_i),
					.op_mod_i(op_mod_i),
					.vectorial_op_i(vectorial_op_i),
					.tag_i(tag_i),
					.in_valid_i(in_valid),
					.in_ready_o(fmt_in_ready[fmt]),
					.flush_i(flush_i),
					.result_o(fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6)) : (((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6))) + ((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))) - 1)-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))]),
					.status_o(fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0) : ((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0)) + 4)-:5]),
					.extension_bit_o(fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 1 : Width + 5)]),
					.tag_o(fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 0 : Width + 6)]),
					.out_valid_o(fmt_out_valid[fmt]),
					.out_ready_i(fmt_out_ready[fmt]),
					.busy_o(fmt_busy[fmt])
				);
			end
			else if ((FpFmtMask[fmt] && ANY_MERGED) && !IS_FIRST_MERGED) begin : merged_unused
				// Trace: design.sv:52370:7
				localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
				// Trace: design.sv:52372:7
				assign fmt_in_ready[fmt] = fmt_in_ready[sv2v_cast_32_signed(FMT)];
				// Trace: design.sv:52374:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: design.sv:52375:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: design.sv:52377:7
				assign fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6)) : (((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6))) + ((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))) - 1)-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: design.sv:52378:7
				assign fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0) : ((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0)) + 4)-:5] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: design.sv:52379:7
				assign fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 1 : Width + 5)] = fpnew_pkg_DONT_CARE;
				// Trace: design.sv:52380:7
				assign fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 0 : Width + 6)] = fpnew_pkg_DONT_CARE;
			end
			else if (!FpFmtMask[fmt] || (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd0)) begin : disable_fmt
				// Trace: design.sv:52384:7
				assign fmt_in_ready[fmt] = 1'b0;
				// Trace: design.sv:52385:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: design.sv:52386:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: design.sv:52388:7
				assign fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6)) : (((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6))) + ((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))) - 1)-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: design.sv:52389:7
				assign fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0) : ((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0)) + 4)-:5] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: design.sv:52390:7
				assign fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 1 : Width + 5)] = fpnew_pkg_DONT_CARE;
				// Trace: design.sv:52391:7
				assign fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 0 : Width + 6)] = fpnew_pkg_DONT_CARE;
			end
		end
	endgenerate
	// Trace: design.sv:52398:3
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:34
		input reg signed [31:0] a;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:41
		input reg signed [31:0] b;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:296:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_get_num_regs_multi;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:484:54
		input reg [159:0] regs;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:485:54
		input reg [9:0] types;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:486:54
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:487:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:488:5
			begin : sv2v_autoblock_7
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:488:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:488:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					begin
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:489:7
						if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2))
							// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:489:41
							res = fpnew_pkg_maximum(res, regs[(4 - i) * 32+:32]);
					end
			end
			fpnew_pkg_get_num_regs_multi = res;
		end
	endfunction
	generate
		if (fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask)) begin : gen_merged_slice
			// Trace: design.sv:52400:5
			localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: design.sv:52401:5
			localparam REG = fpnew_pkg_get_num_regs_multi(FmtPipeRegs, FmtUnitTypes, FpFmtMask);
			// Trace: design.sv:52403:5
			wire in_valid;
			// Trace: design.sv:52405:5
			assign in_valid = in_valid_i & (FmtUnitTypes[(4 - dst_fmt_i) * 2+:2] == 2'd2);
			// Trace: design.sv:52407:5
			fpnew_opgroup_multifmt_slice_23084 #(
				.OpGroup(OpGroup),
				.Width(Width),
				.FpFmtConfig(FpFmtMask),
				.IntFmtConfig(IntFmtMask),
				.EnableVectors(EnableVectors),
				.NumPipeRegs(REG),
				.PipeConfig(PipeConfig)
			) i_multifmt_slice(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i),
				.is_boxed_i(is_boxed_i),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.in_valid_i(in_valid),
				.in_ready_o(fmt_in_ready[FMT]),
				.flush_i(flush_i),
				.result_o(fmt_outputs[((Width + 6) >= 0 ? (FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6)) : (((FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6))) + ((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))) - 1)-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))]),
				.status_o(fmt_outputs[((Width + 6) >= 0 ? (FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0) : ((FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0)) + 4)-:5]),
				.extension_bit_o(fmt_outputs[(FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 1 : Width + 5)]),
				.tag_o(fmt_outputs[(FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 0 : Width + 6)]),
				.out_valid_o(fmt_out_valid[FMT]),
				.out_ready_i(fmt_out_ready[FMT]),
				.busy_o(fmt_busy[FMT])
			);
		end
	endgenerate
	// Trace: design.sv:52446:3
	wire [Width + 6:0] arbiter_output;
	// Trace: design.sv:52449:3
	localparam [31:0] sv2v_uu_i_arbiter_NumIn = NUM_FORMATS;
	localparam [31:0] sv2v_uu_i_arbiter_IdxWidth = $unsigned(3);
	// removed localparam type sv2v_uu_i_arbiter_rr_i
	localparam [sv2v_uu_i_arbiter_IdxWidth - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_3ECCC_46CA0 #(
		.DataType_Width(Width),
		.NumIn(NUM_FORMATS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
		.req_i(fmt_out_valid),
		.gnt_o(fmt_out_ready),
		.data_i(fmt_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: design.sv:52468:3
	assign result_o = arbiter_output[Width + 6-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))];
	// Trace: design.sv:52469:3
	assign status_o = arbiter_output[6-:5];
	// Trace: design.sv:52470:3
	assign extension_bit_o = arbiter_output[1];
	// Trace: design.sv:52471:3
	assign tag_o = arbiter_output[0];
	// Trace: design.sv:52473:3
	assign busy_o = |fmt_busy;
endmodule
module fpnew_opgroup_fmt_slice_07650 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	reg _sv2v_0;
	// Trace: design.sv:52492:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: design.sv:52493:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_5D882(0);
	// Trace: design.sv:52495:13
	parameter [31:0] Width = 32;
	// Trace: design.sv:52496:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: design.sv:52497:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: design.sv:52498:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: design.sv:52499:38
	// removed localparam type TagType
	// Trace: design.sv:52501:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:378:48
		input reg [1:0] grp;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:379:5
		(* full_case, parallel_case *)
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: design.sv:52503:3
	input wire clk_i;
	// Trace: design.sv:52504:3
	input wire rst_ni;
	// Trace: design.sv:52506:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: design.sv:52507:3
	input wire [NUM_OPERANDS - 1:0] is_boxed_i;
	// Trace: design.sv:52508:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:52509:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:52510:3
	input wire op_mod_i;
	// Trace: design.sv:52511:3
	input wire vectorial_op_i;
	// Trace: design.sv:52512:3
	input wire tag_i;
	// Trace: design.sv:52514:3
	input wire in_valid_i;
	// Trace: design.sv:52515:3
	output wire in_ready_o;
	// Trace: design.sv:52516:3
	input wire flush_i;
	// Trace: design.sv:52518:3
	output wire [Width - 1:0] result_o;
	// Trace: design.sv:52519:3
	// removed localparam type fpnew_pkg_status_t
	output reg [4:0] status_o;
	// Trace: design.sv:52520:3
	output wire extension_bit_o;
	// Trace: design.sv:52521:3
	output wire tag_o;
	// Trace: design.sv:52523:3
	output wire out_valid_o;
	// Trace: design.sv:52524:3
	input wire out_ready_i;
	// Trace: design.sv:52526:3
	output wire busy_o;
	// Trace: design.sv:52529:3
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: design.sv:52530:3
	function automatic [31:0] fpnew_pkg_num_lanes;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:389:45
		input reg [31:0] width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:389:65
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:389:82
		input reg vec;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:390:5
		fpnew_pkg_num_lanes = (vec ? width / fpnew_pkg_fp_width(fmt) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_num_lanes(Width, FpFormat, EnableVectors);
	// Trace: design.sv:52533:3
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	// Trace: design.sv:52534:3
	wire vectorial_op;
	// Trace: design.sv:52536:3
	wire [(NUM_LANES * FP_WIDTH) - 1:0] slice_result;
	// Trace: design.sv:52537:3
	wire [Width - 1:0] slice_regular_result;
	wire [Width - 1:0] slice_class_result;
	wire [Width - 1:0] slice_vec_class_result;
	// Trace: design.sv:52539:3
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	// Trace: design.sv:52540:3
	wire [NUM_LANES - 1:0] lane_ext_bit;
	// Trace: design.sv:52541:3
	// removed localparam type fpnew_pkg_classmask_e
	wire [(NUM_LANES * 10) - 1:0] lane_class_mask;
	// Trace: design.sv:52542:3
	wire [NUM_LANES - 1:0] lane_tags;
	// Trace: design.sv:52543:3
	wire [NUM_LANES - 1:0] lane_vectorial;
	wire [NUM_LANES - 1:0] lane_busy;
	wire [NUM_LANES - 1:0] lane_is_class;
	// Trace: design.sv:52545:3
	wire result_is_vector;
	wire result_is_class;
	// Trace: design.sv:52550:3
	assign in_ready_o = lane_in_ready[0];
	// Trace: design.sv:52551:3
	assign vectorial_op = vectorial_op_i & EnableVectors;
	// Trace: design.sv:52556:3
	genvar _gv_lane_1;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_lane_1 = 0; _gv_lane_1 < sv2v_cast_32_signed(NUM_LANES); _gv_lane_1 = _gv_lane_1 + 1) begin : gen_num_lanes
			localparam lane = _gv_lane_1;
			// Trace: design.sv:52557:5
			wire [FP_WIDTH - 1:0] local_result;
			// Trace: design.sv:52558:5
			wire local_sign;
			if ((lane == 0) || EnableVectors) begin : active_lane
				// Trace: design.sv:52562:7
				wire in_valid;
				wire out_valid;
				wire out_ready;
				// Trace: design.sv:52564:7
				reg [(NUM_OPERANDS * FP_WIDTH) - 1:0] local_operands;
				// Trace: design.sv:52565:7
				wire [FP_WIDTH - 1:0] op_result;
				// Trace: design.sv:52566:7
				wire [4:0] op_status;
				// Trace: design.sv:52568:7
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				// Trace: design.sv:52570:7
				always @(*) begin : prepare_input
					if (_sv2v_0)
						;
					// Trace: design.sv:52571:9
					begin : sv2v_autoblock_1
						// Trace: design.sv:52571:14
						reg signed [31:0] i;
						// Trace: design.sv:52571:14
						for (i = 0; i < sv2v_cast_32_signed(NUM_OPERANDS); i = i + 1)
							begin
								// Trace: design.sv:52572:11
								local_operands[i * FP_WIDTH+:FP_WIDTH] = operands_i[(i * Width) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (($unsigned(lane) + 1) * FP_WIDTH) - 1 : (((($unsigned(lane) + 1) * FP_WIDTH) - 1) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:(((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)];
							end
					end
				end
				if (OpGroup == 2'd0) begin : lane_instance
					// Trace: design.sv:52578:9
					fpnew_fma_EA93F #(
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fma(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
					// Trace: design.sv:52606:9
					assign lane_is_class[lane] = 1'b0;
					// Trace: design.sv:52607:9
					assign lane_class_mask[lane * 10+:10] = 10'b0000000001;
				end
				else if (OpGroup == 2'd1) begin
					;
				end
				else if (OpGroup == 2'd2) begin : lane_instance
					// Trace: design.sv:52639:9
					fpnew_noncomp_DE16F #(
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_noncomp(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.class_mask_o(lane_class_mask[lane * 10+:10]),
						.is_class_o(lane_is_class[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				// Trace: design.sv:52672:7
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				// Trace: design.sv:52673:7
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				// Trace: design.sv:52676:7
				assign local_result = (lane_out_valid[lane] ? op_result : {FP_WIDTH {lane_ext_bit[0]}});
				// Trace: design.sv:52677:7
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] ? op_status : {5 {1'sb0}});
			end
			else begin : genblk1
				// Trace: design.sv:52681:7
				assign lane_out_valid[lane] = 1'b0;
				// Trace: design.sv:52682:7
				assign lane_in_ready[lane] = 1'b0;
				// Trace: design.sv:52683:7
				assign local_result = {FP_WIDTH {lane_ext_bit[0]}};
				// Trace: design.sv:52684:7
				assign lane_status[lane * 5+:5] = 1'sb0;
				// Trace: design.sv:52685:7
				assign lane_busy[lane] = 1'b0;
				// Trace: design.sv:52686:7
				assign lane_is_class[lane] = 1'b0;
			end
			// Trace: design.sv:52690:5
			assign slice_result[(($unsigned(lane) + 1) * FP_WIDTH) - 1:$unsigned(lane) * FP_WIDTH] = local_result;
			if (((lane + 1) * 8) <= Width) begin : vectorial_class
				// Trace: design.sv:52694:7
				assign local_sign = (((lane_class_mask[lane * 10+:10] == 10'b0000000001) || (lane_class_mask[lane * 10+:10] == 10'b0000000010)) || (lane_class_mask[lane * 10+:10] == 10'b0000000100)) || (lane_class_mask[lane * 10+:10] == 10'b0000001000);
				// Trace: design.sv:52699:7
				assign slice_vec_class_result[((lane + 1) * 8) - 1:lane * 8] = {local_sign, ~local_sign, lane_class_mask[lane * 10+:10] == 10'b1000000000, lane_class_mask[lane * 10+:10] == 10'b0100000000, (lane_class_mask[lane * 10+:10] == 10'b0000010000) || (lane_class_mask[lane * 10+:10] == 10'b0000001000), (lane_class_mask[lane * 10+:10] == 10'b0000100000) || (lane_class_mask[lane * 10+:10] == 10'b0000000100), (lane_class_mask[lane * 10+:10] == 10'b0001000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000010), (lane_class_mask[lane * 10+:10] == 10'b0010000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000001)};
			end
		end
	endgenerate
	// Trace: design.sv:52719:3
	assign result_is_vector = lane_vectorial[0];
	// Trace: design.sv:52720:3
	assign result_is_class = lane_is_class[0];
	// Trace: design.sv:52722:3
	assign slice_regular_result = $signed({extension_bit_o, slice_result});
	// Trace: design.sv:52724:3
	localparam [31:0] CLASS_VEC_BITS = ((NUM_LANES * 8) > Width ? 8 * (Width / 8) : NUM_LANES * 8);
	// Trace: design.sv:52727:3
	generate
		if (CLASS_VEC_BITS < Width) begin : pad_vectorial_class
			// Trace: design.sv:52728:5
			assign slice_vec_class_result[Width - 1:CLASS_VEC_BITS] = 1'sb0;
		end
	endgenerate
	// Trace: design.sv:52733:3
	assign slice_class_result = (result_is_vector ? slice_vec_class_result : lane_class_mask[0+:10]);
	// Trace: design.sv:52736:3
	assign result_o = (result_is_class ? slice_class_result : slice_regular_result);
	// Trace: design.sv:52738:3
	assign extension_bit_o = lane_ext_bit[0];
	// Trace: design.sv:52739:3
	assign tag_o = lane_tags[0];
	// Trace: design.sv:52740:3
	assign busy_o = |lane_busy;
	// Trace: design.sv:52741:3
	assign out_valid_o = lane_out_valid[0];
	// Trace: design.sv:52745:3
	always @(*) begin : output_processing
		// Trace: design.sv:52747:5
		reg [4:0] temp_status;
		if (_sv2v_0)
			;
		// Trace: design.sv:52748:5
		temp_status = 1'sb0;
		// Trace: design.sv:52749:5
		begin : sv2v_autoblock_2
			// Trace: design.sv:52749:10
			reg signed [31:0] i;
			// Trace: design.sv:52749:10
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				begin
					// Trace: design.sv:52750:7
					temp_status = temp_status | lane_status[i * 5+:5];
				end
		end
		// Trace: design.sv:52751:5
		status_o = temp_status;
	end
	initial _sv2v_0 = 0;
endmodule
module fpnew_opgroup_multifmt_slice_23084 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	reg _sv2v_0;
	// Trace: design.sv:52772:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd3;
	// Trace: design.sv:52773:13
	parameter [31:0] Width = 64;
	// Trace: design.sv:52775:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: design.sv:52776:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtConfig = 1'sb1;
	// Trace: design.sv:52777:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: design.sv:52778:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: design.sv:52779:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: design.sv:52780:38
	// removed localparam type TagType
	// Trace: design.sv:52782:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:378:48
		input reg [1:0] grp;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:379:5
		(* full_case, parallel_case *)
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: design.sv:52783:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: design.sv:52785:3
	input wire clk_i;
	// Trace: design.sv:52786:3
	input wire rst_ni;
	// Trace: design.sv:52788:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: design.sv:52789:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: design.sv:52790:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:52791:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:52792:3
	input wire op_mod_i;
	// Trace: design.sv:52793:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: design.sv:52794:3
	input wire [2:0] dst_fmt_i;
	// Trace: design.sv:52795:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: design.sv:52796:3
	input wire vectorial_op_i;
	// Trace: design.sv:52797:3
	input wire tag_i;
	// Trace: design.sv:52799:3
	input wire in_valid_i;
	// Trace: design.sv:52800:3
	output wire in_ready_o;
	// Trace: design.sv:52801:3
	input wire flush_i;
	// Trace: design.sv:52803:3
	output wire [Width - 1:0] result_o;
	// Trace: design.sv:52804:3
	// removed localparam type fpnew_pkg_status_t
	output reg [4:0] status_o;
	// Trace: design.sv:52805:3
	output wire extension_bit_o;
	// Trace: design.sv:52806:3
	output wire tag_o;
	// Trace: design.sv:52808:3
	output wire out_valid_o;
	// Trace: design.sv:52809:3
	input wire out_ready_i;
	// Trace: design.sv:52811:3
	output wire busy_o;
	// Trace: design.sv:52814:3
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:34
		input reg signed [31:0] a;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:295:41
		input reg signed [31:0] b;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:296:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:308:48
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:309:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:5
			begin : sv2v_autoblock_1
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:310:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:312:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] MAX_FP_WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: design.sv:52815:3
	function automatic [1:0] sv2v_cast_CDB06;
		input reg [1:0] inp;
		sv2v_cast_CDB06 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:88:45
		input reg [1:0] ifmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:89:5
		(* full_case, parallel_case *)
		case (ifmt)
			sv2v_cast_CDB06(0): fpnew_pkg_int_width = 8;
			sv2v_cast_CDB06(1): fpnew_pkg_int_width = 16;
			sv2v_cast_CDB06(2): fpnew_pkg_int_width = 32;
			sv2v_cast_CDB06(3): fpnew_pkg_int_width = 64;
			default: begin
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:96:9
				$fatal(1, "Invalid INT format supplied");
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:100:9
				fpnew_pkg_int_width = sv2v_cast_CDB06(0);
			end
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:355:49
		input reg [0:3] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:356:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:357:5
			begin : sv2v_autoblock_2
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:357:10
				reg signed [31:0] ifmt;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:357:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:358:7
						if (cfg[ifmt])
							// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:358:22
							res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_CDB06(ifmt)));
					end
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	// Trace: design.sv:52816:3
	function automatic signed [31:0] fpnew_pkg_minimum;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:291:34
		input reg signed [31:0] a;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:291:41
		input reg signed [31:0] b;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:292:5
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:317:48
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:318:5
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:319:5
			begin : sv2v_autoblock_3
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:319:10
				reg [31:0] i;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:319:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:321:9
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:394:49
		input reg [31:0] width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:394:69
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:394:86
		input reg vec;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:395:5
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_max_num_lanes(Width, FpFmtConfig, 1'b1);
	// Trace: design.sv:52817:3
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	// Trace: design.sv:52819:3
	localparam [31:0] FMT_BITS = fpnew_pkg_maximum(3, 2);
	// Trace: design.sv:52821:3
	localparam [31:0] AUX_BITS = FMT_BITS + 2;
	// Trace: design.sv:52823:3
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	// Trace: design.sv:52824:3
	wire vectorial_op;
	// Trace: design.sv:52825:3
	wire [FMT_BITS - 1:0] dst_fmt;
	// Trace: design.sv:52826:3
	wire [AUX_BITS - 1:0] aux_data;
	// Trace: design.sv:52829:3
	wire dst_fmt_is_int;
	wire dst_is_cpk;
	// Trace: design.sv:52830:3
	wire [1:0] dst_vec_op;
	// Trace: design.sv:52831:3
	wire [2:0] target_aux_d;
	wire [2:0] target_aux_q;
	// Trace: design.sv:52832:3
	wire is_up_cast;
	wire is_down_cast;
	// Trace: design.sv:52834:3
	wire [(NUM_FORMATS * Width) - 1:0] fmt_slice_result;
	// Trace: design.sv:52835:3
	wire [(NUM_INT_FORMATS * Width) - 1:0] ifmt_slice_result;
	// Trace: design.sv:52836:3
	wire [Width - 1:0] conv_slice_result;
	// Trace: design.sv:52839:3
	wire [Width - 1:0] conv_target_d;
	wire [Width - 1:0] conv_target_q;
	// Trace: design.sv:52841:3
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	// Trace: design.sv:52842:3
	wire [NUM_LANES - 1:0] lane_ext_bit;
	// Trace: design.sv:52843:3
	wire [NUM_LANES - 1:0] lane_tags;
	// Trace: design.sv:52844:3
	wire [(NUM_LANES * AUX_BITS) - 1:0] lane_aux;
	// Trace: design.sv:52845:3
	wire [NUM_LANES - 1:0] lane_busy;
	// Trace: design.sv:52847:3
	wire result_is_vector;
	// Trace: design.sv:52848:3
	wire [FMT_BITS - 1:0] result_fmt;
	// Trace: design.sv:52849:3
	wire result_fmt_is_int;
	wire result_is_cpk;
	// Trace: design.sv:52850:3
	wire [1:0] result_vec_op;
	// Trace: design.sv:52855:3
	assign in_ready_o = lane_in_ready[0];
	// Trace: design.sv:52856:3
	assign vectorial_op = vectorial_op_i & EnableVectors;
	// Trace: design.sv:52859:3
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	assign dst_fmt_is_int = (OpGroup == 2'd3) & (op_i == sv2v_cast_4CD2E(11));
	// Trace: design.sv:52860:3
	assign dst_is_cpk = (OpGroup == 2'd3) & ((op_i == sv2v_cast_4CD2E(13)) || (op_i == sv2v_cast_4CD2E(14)));
	// Trace: design.sv:52862:3
	assign dst_vec_op = (OpGroup == 2'd3) & {op_i == sv2v_cast_4CD2E(14), op_mod_i};
	// Trace: design.sv:52864:3
	assign is_up_cast = fpnew_pkg_fp_width(dst_fmt_i) > fpnew_pkg_fp_width(src_fmt_i);
	// Trace: design.sv:52865:3
	assign is_down_cast = fpnew_pkg_fp_width(dst_fmt_i) < fpnew_pkg_fp_width(src_fmt_i);
	// Trace: design.sv:52868:3
	assign dst_fmt = (dst_fmt_is_int ? int_fmt_i : dst_fmt_i);
	// Trace: design.sv:52871:3
	assign aux_data = {dst_fmt_is_int, vectorial_op, dst_fmt};
	// Trace: design.sv:52872:3
	assign target_aux_d = {dst_vec_op, dst_is_cpk};
	// Trace: design.sv:52875:3
	generate
		if (OpGroup == 2'd3) begin : conv_target
			// Trace: design.sv:52876:5
			assign conv_target_d = (dst_is_cpk ? operands_i[2 * Width+:Width] : operands_i[Width+:Width]);
		end
	endgenerate
	// Trace: design.sv:52880:3
	reg [4:0] is_boxed_1op;
	// Trace: design.sv:52881:3
	reg [9:0] is_boxed_2op;
	// Trace: design.sv:52883:3
	always @(*) begin : boxed_2op
		if (_sv2v_0)
			;
		// Trace: design.sv:52884:5
		begin : sv2v_autoblock_4
			// Trace: design.sv:52884:10
			reg signed [31:0] fmt;
			// Trace: design.sv:52884:10
			for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
				begin
					// Trace: design.sv:52885:7
					is_boxed_1op[fmt] = is_boxed_i[fmt * NUM_OPERANDS];
					// Trace: design.sv:52886:7
					is_boxed_2op[fmt * 2+:2] = is_boxed_i[(fmt * NUM_OPERANDS) + 1-:2];
				end
		end
	end
	// Trace: design.sv:52893:3
	genvar _gv_lane_2;
	localparam [0:4] fpnew_pkg_CPK_FORMATS = 5'b11000;
	function automatic [0:4] fpnew_pkg_get_conv_lane_formats;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:428:56
		input reg [31:0] width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:429:56
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:430:56
		input reg [31:0] lane_no;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:431:5
		reg [0:4] res;
		begin
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:432:5
			begin : sv2v_autoblock_5
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:432:10
				reg [31:0] fmt;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:432:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					begin
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:434:7
						res[fmt] = cfg[fmt] && (((width / fpnew_pkg_fp_width(sv2v_cast_5D882(fmt))) > lane_no) || (fpnew_pkg_CPK_FORMATS[fmt] && (lane_no < 2)));
					end
			end
			fpnew_pkg_get_conv_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_conv_lane_int_formats;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:440:61
		input reg [31:0] width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:441:61
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:442:61
		input reg [0:3] icfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:443:61
		input reg [31:0] lane_no;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:444:5
		reg [0:3] res;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:445:5
		reg [0:4] lanefmts;
		begin
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:446:5
			res = 1'sb0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:447:5
			lanefmts = fpnew_pkg_get_conv_lane_formats(width, cfg, lane_no);
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:449:5
			begin : sv2v_autoblock_6
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:449:10
				reg [31:0] ifmt;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:449:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_7
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:450:12
						reg [31:0] fmt;
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:450:12
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							begin
								// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:452:9
								res[ifmt] = res[ifmt] | ((icfg[ifmt] && lanefmts[fmt]) && (fpnew_pkg_fp_width(sv2v_cast_5D882(fmt)) == fpnew_pkg_int_width(sv2v_cast_CDB06(ifmt))));
							end
					end
			end
			fpnew_pkg_get_conv_lane_int_formats = res;
		end
	endfunction
	function automatic [0:4] fpnew_pkg_get_lane_formats;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:399:51
		input reg [31:0] width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:400:51
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:401:51
		input reg [31:0] lane_no;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:402:5
		reg [0:4] res;
		begin
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:403:5
			begin : sv2v_autoblock_8
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:403:10
				reg [31:0] fmt;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:403:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					begin
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:405:7
						res[fmt] = cfg[fmt] & ((width / fpnew_pkg_fp_width(sv2v_cast_5D882(fmt))) > lane_no);
					end
			end
			fpnew_pkg_get_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_lane_int_formats;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:410:56
		input reg [31:0] width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:411:56
		input reg [0:4] cfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:412:56
		input reg [0:3] icfg;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:413:56
		input reg [31:0] lane_no;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:414:5
		reg [0:3] res;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:415:5
		reg [0:4] lanefmts;
		begin
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:416:5
			res = 1'sb0;
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:417:5
			lanefmts = fpnew_pkg_get_lane_formats(width, cfg, lane_no);
			// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:419:5
			begin : sv2v_autoblock_9
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:419:10
				reg [31:0] ifmt;
				// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:419:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_10
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:420:12
						reg [31:0] fmt;
						// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:420:12
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							if (fpnew_pkg_fp_width(sv2v_cast_5D882(fmt)) == fpnew_pkg_int_width(sv2v_cast_CDB06(ifmt)))
								// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:423:11
								res[ifmt] = res[ifmt] | (icfg[ifmt] && lanefmts[fmt]);
					end
			end
			fpnew_pkg_get_lane_int_formats = res;
		end
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [4:0] sv2v_cast_F930B;
		input reg [4:0] inp;
		sv2v_cast_F930B = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_lane_2 = 0; _gv_lane_2 < sv2v_cast_32_signed(NUM_LANES); _gv_lane_2 = _gv_lane_2 + 1) begin : gen_num_lanes
			localparam lane = _gv_lane_2;
			// Trace: design.sv:52894:5
			localparam [31:0] LANE = $unsigned(lane);
			// Trace: design.sv:52896:5
			localparam [0:4] ACTIVE_FORMATS = fpnew_pkg_get_lane_formats(Width, FpFmtConfig, LANE);
			// Trace: design.sv:52898:5
			localparam [0:3] ACTIVE_INT_FORMATS = fpnew_pkg_get_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			// Trace: design.sv:52900:5
			localparam [31:0] MAX_WIDTH = fpnew_pkg_max_fp_width(ACTIVE_FORMATS);
			// Trace: design.sv:52903:5
			localparam [0:4] CONV_FORMATS = fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, LANE);
			// Trace: design.sv:52905:5
			localparam [0:3] CONV_INT_FORMATS = fpnew_pkg_get_conv_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			// Trace: design.sv:52907:5
			localparam [31:0] CONV_WIDTH = fpnew_pkg_max_fp_width(CONV_FORMATS);
			// Trace: design.sv:52910:5
			localparam [0:4] LANE_FORMATS = (OpGroup == 2'd3 ? CONV_FORMATS : ACTIVE_FORMATS);
			// Trace: design.sv:52912:5
			localparam [31:0] LANE_WIDTH = (OpGroup == 2'd3 ? CONV_WIDTH : MAX_WIDTH);
			// Trace: design.sv:52914:5
			wire [LANE_WIDTH - 1:0] local_result;
			if ((lane == 0) || EnableVectors) begin : active_lane
				// Trace: design.sv:52918:7
				wire in_valid;
				wire out_valid;
				wire out_ready;
				// Trace: design.sv:52920:7
				reg [(NUM_OPERANDS * LANE_WIDTH) - 1:0] local_operands;
				// Trace: design.sv:52921:7
				wire [LANE_WIDTH - 1:0] op_result;
				// Trace: design.sv:52922:7
				wire [4:0] op_status;
				// Trace: design.sv:52924:7
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				// Trace: design.sv:52927:7
				always @(*) begin : prepare_input
					if (_sv2v_0)
						;
					// Trace: design.sv:52928:9
					begin : sv2v_autoblock_11
						// Trace: design.sv:52928:14
						reg [31:0] i;
						// Trace: design.sv:52928:14
						for (i = 0; i < NUM_OPERANDS; i = i + 1)
							begin
								// Trace: design.sv:52929:11
								local_operands[i * (OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))))+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))))] = operands_i[i * Width+:Width] >> (LANE * fpnew_pkg_fp_width(src_fmt_i));
							end
					end
					if (OpGroup == 2'd3) begin
						begin
							// Trace: design.sv:52935:11
							if (op_i == sv2v_cast_4CD2E(12))
								// Trace: design.sv:52936:13
								local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))))] = operands_i[0+:Width] >> (LANE * fpnew_pkg_int_width(int_fmt_i));
							else if (op_i == sv2v_cast_4CD2E(10)) begin
								begin
									// Trace: design.sv:52939:13
									if ((vectorial_op && op_mod_i) && is_up_cast)
										// Trace: design.sv:52940:15
										local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))))] = operands_i[0+:Width] >> ((LANE * fpnew_pkg_fp_width(src_fmt_i)) + (MAX_FP_WIDTH / 2));
								end
							end
							else if (dst_is_cpk) begin
								begin
									// Trace: design.sv:52945:13
									if (lane == 1)
										// Trace: design.sv:52946:15
										local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))))] = operands_i[Width + (LANE_WIDTH - 1)-:LANE_WIDTH];
								end
							end
						end
					end
				end
				if (OpGroup == 2'd0) begin : lane_instance
					// Trace: design.sv:52954:9
					fpnew_fma_multi_B5D6B_A0513 #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_fma_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				else if (OpGroup == 2'd1) begin : lane_instance
					// Trace: design.sv:52986:9
					fpnew_divsqrt_multi_E225A_955F4 #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_divsqrt_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2))))) * 2]),
						.is_boxed_i(is_boxed_2op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				else if (OpGroup == 2'd2) begin
					;
				end
				else if (OpGroup == 2'd3) begin : lane_instance
					// Trace: design.sv:53017:9
					fpnew_cast_multi_2E827_EA7A2 #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.IntFmtConfig(CONV_INT_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_cast_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))))]),
						.is_boxed_i(is_boxed_1op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.int_fmt_i(int_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				// Trace: design.sv:53052:7
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				// Trace: design.sv:53053:7
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				// Trace: design.sv:53056:7
				assign local_result = (lane_out_valid[lane] ? op_result : {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F930B(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2))))) : fpnew_pkg_max_fp_width(sv2v_cast_F930B(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))))) {lane_ext_bit[0]}});
				// Trace: design.sv:53057:7
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] ? op_status : {5 {1'sb0}});
			end
			else begin : inactive_lane
				// Trace: design.sv:53061:7
				assign lane_out_valid[lane] = 1'b0;
				// Trace: design.sv:53062:7
				assign lane_in_ready[lane] = 1'b0;
				// Trace: design.sv:53063:7
				assign local_result = {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F930B(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2))))) : fpnew_pkg_max_fp_width(sv2v_cast_F930B(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_2)))))) {lane_ext_bit[0]}};
				// Trace: design.sv:53064:7
				assign lane_status[lane * 5+:5] = 1'sb0;
				// Trace: design.sv:53065:7
				assign lane_busy[lane] = 1'b0;
			end
			genvar _gv_fmt_10;
			for (_gv_fmt_10 = 0; _gv_fmt_10 < NUM_FORMATS; _gv_fmt_10 = _gv_fmt_10 + 1) begin : pack_fp_result
				localparam fmt = _gv_fmt_10;
				// Trace: design.sv:53071:7
				localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
				if (ACTIVE_FORMATS[fmt]) begin : genblk1
					// Trace: design.sv:53074:9
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = local_result[FP_WIDTH - 1:0];
				end
				else if (((LANE + 1) * FP_WIDTH) <= Width) begin : genblk1
					// Trace: design.sv:53077:9
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = {((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1) {lane_ext_bit[LANE]}};
				end
				else if ((LANE * FP_WIDTH) < Width) begin : genblk1
					// Trace: design.sv:53080:9
					assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (LANE * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[LANE]}};
				end
			end
			if (OpGroup == 2'd3) begin : int_results_enabled
				genvar _gv_ifmt_4;
				for (_gv_ifmt_4 = 0; _gv_ifmt_4 < NUM_INT_FORMATS; _gv_ifmt_4 = _gv_ifmt_4 + 1) begin : pack_int_result
					localparam ifmt = _gv_ifmt_4;
					// Trace: design.sv:53089:9
					localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_CDB06(ifmt));
					if (ACTIVE_INT_FORMATS[ifmt]) begin : genblk1
						// Trace: design.sv:53091:11
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = local_result[INT_WIDTH - 1:0];
					end
					else if (((LANE + 1) * INT_WIDTH) <= Width) begin : genblk1
						// Trace: design.sv:53094:11
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = 1'sb0;
					end
					else if ((LANE * INT_WIDTH) < Width) begin : genblk1
						// Trace: design.sv:53096:11
						assign ifmt_slice_result[(ifmt * Width) + ((Width - 1) >= (LANE * INT_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (LANE * INT_WIDTH) ? ((Width - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (LANE * INT_WIDTH) ? ((Width - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (Width - 1)) + 1)] = 1'sb0;
					end
				end
			end
		end
	endgenerate
	// Trace: design.sv:53103:3
	genvar _gv_fmt_11;
	generate
		for (_gv_fmt_11 = 0; _gv_fmt_11 < NUM_FORMATS; _gv_fmt_11 = _gv_fmt_11 + 1) begin : extend_fp_result
			localparam fmt = _gv_fmt_11;
			// Trace: design.sv:53105:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			if ((NUM_LANES * FP_WIDTH) < Width) begin : genblk1
				// Trace: design.sv:53107:7
				assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[0]}};
			end
		end
	endgenerate
	// Trace: design.sv:53111:3
	genvar _gv_ifmt_5;
	generate
		for (_gv_ifmt_5 = 0; _gv_ifmt_5 < NUM_INT_FORMATS; _gv_ifmt_5 = _gv_ifmt_5 + 1) begin : int_results_disabled
			localparam ifmt = _gv_ifmt_5;
			if (OpGroup != 2'd3) begin : mute_int_result
				// Trace: design.sv:53113:7
				assign ifmt_slice_result[ifmt * Width+:Width] = 1'sb0;
			end
		end
	endgenerate
	// Trace: design.sv:53118:3
	generate
		if (OpGroup == 2'd3) begin : target_regs
			// Trace: design.sv:53120:5
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * Width) + ((NumPipeRegs * Width) - 1) : ((NumPipeRegs + 1) * Width) - 1):(0 >= NumPipeRegs ? NumPipeRegs * Width : 0)] byp_pipe_target_q;
			// Trace: design.sv:53121:5
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * 3) + ((NumPipeRegs * 3) - 1) : ((NumPipeRegs + 1) * 3) - 1):(0 >= NumPipeRegs ? NumPipeRegs * 3 : 0)] byp_pipe_aux_q;
			// Trace: design.sv:53122:5
			reg [0:NumPipeRegs] byp_pipe_valid_q;
			// Trace: design.sv:53124:5
			wire [0:NumPipeRegs] byp_pipe_ready;
			// Trace: design.sv:53127:5
			wire [Width * 1:1] sv2v_tmp_341F5;
			assign sv2v_tmp_341F5 = conv_target_d;
			always @(*) byp_pipe_target_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * Width+:Width] = sv2v_tmp_341F5;
			// Trace: design.sv:53128:5
			wire [3:1] sv2v_tmp_5E9D8;
			assign sv2v_tmp_5E9D8 = target_aux_d;
			always @(*) byp_pipe_aux_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * 3+:3] = sv2v_tmp_5E9D8;
			// Trace: design.sv:53129:5
			wire [1:1] sv2v_tmp_967FD;
			assign sv2v_tmp_967FD = in_valid_i & vectorial_op;
			always @(*) byp_pipe_valid_q[0] = sv2v_tmp_967FD;
			genvar _gv_i_82;
			for (_gv_i_82 = 0; _gv_i_82 < NumPipeRegs; _gv_i_82 = _gv_i_82 + 1) begin : gen_bypass_pipeline
				localparam i = _gv_i_82;
				// Trace: design.sv:53133:7
				wire reg_ena;
				// Trace: design.sv:53137:7
				assign byp_pipe_ready[i] = byp_pipe_ready[i + 1] | ~byp_pipe_valid_q[i + 1];
				// Trace: macro expansion of FFLARNC at design.sv:53139:331
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFLARNC at design.sv:53139:409
					if (!rst_ni)
						// Trace: macro expansion of FFLARNC at design.sv:53139:487
						byp_pipe_valid_q[i + 1] <= 1'b0;
					else
						// Trace: macro expansion of FFLARNC at design.sv:53139:639
						if (flush_i)
							// Trace: macro expansion of FFLARNC at design.sv:53139:717
							byp_pipe_valid_q[i + 1] <= 1'b0;
						else if (byp_pipe_ready[i])
							// Trace: macro expansion of FFLARNC at design.sv:53139:869
							byp_pipe_valid_q[i + 1] <= byp_pipe_valid_q[i];
				// Trace: design.sv:53141:7
				assign reg_ena = byp_pipe_ready[i] & byp_pipe_valid_q[i];
				// Trace: macro expansion of FFL at design.sv:53143:71
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFL at design.sv:53143:168
					if (!rst_ni)
						// Trace: macro expansion of FFL at design.sv:53143:265
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= 1'sb0;
					else
						// Trace: macro expansion of FFL at design.sv:53143:455
						if (reg_ena)
							// Trace: macro expansion of FFL at design.sv:53143:552
							byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= byp_pipe_target_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * Width+:Width];
				// Trace: macro expansion of FFL at design.sv:53144:71
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFL at design.sv:53144:168
					if (!rst_ni)
						// Trace: macro expansion of FFL at design.sv:53144:265
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= 1'sb0;
					else
						// Trace: macro expansion of FFL at design.sv:53144:455
						if (reg_ena)
							// Trace: macro expansion of FFL at design.sv:53144:552
							byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= byp_pipe_aux_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * 3+:3];
			end
			// Trace: design.sv:53147:5
			assign byp_pipe_ready[NumPipeRegs] = out_ready_i & result_is_vector;
			// Trace: design.sv:53149:5
			assign conv_target_q = byp_pipe_target_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * Width+:Width];
			// Trace: design.sv:53152:5
			assign {result_vec_op, result_is_cpk} = byp_pipe_aux_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * 3+:3];
		end
		else begin : no_conv
			// Trace: design.sv:53154:5
			assign {result_vec_op, result_is_cpk} = 1'sb0;
		end
	endgenerate
	// Trace: design.sv:53160:3
	assign {result_fmt_is_int, result_is_vector, result_fmt} = lane_aux[0+:AUX_BITS];
	// Trace: design.sv:53162:3
	assign result_o = (result_fmt_is_int ? ifmt_slice_result[result_fmt * Width+:Width] : fmt_slice_result[result_fmt * Width+:Width]);
	// Trace: design.sv:53166:3
	assign extension_bit_o = lane_ext_bit[0];
	// Trace: design.sv:53167:3
	assign tag_o = lane_tags[0];
	// Trace: design.sv:53168:3
	assign busy_o = |lane_busy;
	// Trace: design.sv:53170:3
	assign out_valid_o = lane_out_valid[0];
	// Trace: design.sv:53173:3
	always @(*) begin : output_processing
		// Trace: design.sv:53175:5
		reg [4:0] temp_status;
		if (_sv2v_0)
			;
		// Trace: design.sv:53176:5
		temp_status = 1'sb0;
		// Trace: design.sv:53177:5
		begin : sv2v_autoblock_12
			// Trace: design.sv:53177:10
			reg signed [31:0] i;
			// Trace: design.sv:53177:10
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				begin
					// Trace: design.sv:53178:7
					temp_status = temp_status | lane_status[i * 5+:5];
				end
		end
		// Trace: design.sv:53179:5
		status_o = temp_status;
	end
	initial _sv2v_0 = 0;
endmodule
module fpnew_rounding (
	abs_value_i,
	sign_i,
	round_sticky_bits_i,
	rnd_mode_i,
	effective_subtraction_i,
	abs_rounded_o,
	sign_o,
	exact_zero_o
);
	reg _sv2v_0;
	// Trace: design.sv:53198:13
	parameter [31:0] AbsWidth = 2;
	// Trace: design.sv:53201:3
	input wire [AbsWidth - 1:0] abs_value_i;
	// Trace: design.sv:53202:3
	input wire sign_i;
	// Trace: design.sv:53204:3
	input wire [1:0] round_sticky_bits_i;
	// Trace: design.sv:53205:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:53206:3
	input wire effective_subtraction_i;
	// Trace: design.sv:53208:3
	output wire [AbsWidth - 1:0] abs_rounded_o;
	// Trace: design.sv:53209:3
	output wire sign_o;
	// Trace: design.sv:53211:3
	output wire exact_zero_o;
	// Trace: design.sv:53214:3
	reg round_up;
	// Trace: design.sv:53225:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	always @(*) begin : rounding_decision
		if (_sv2v_0)
			;
		// Trace: design.sv:53226:5
		(* full_case, parallel_case *)
		case (rnd_mode_i)
			3'b000:
				(* full_case, parallel_case *)
				case (round_sticky_bits_i)
					2'b00, 2'b01:
						// Trace: design.sv:53230:18
						round_up = 1'b0;
					2'b10:
						// Trace: design.sv:53231:18
						round_up = abs_value_i[0];
					2'b11:
						// Trace: design.sv:53232:18
						round_up = 1'b1;
					default:
						// Trace: design.sv:53233:20
						round_up = fpnew_pkg_DONT_CARE;
				endcase
			3'b001:
				// Trace: design.sv:53235:23
				round_up = 1'b0;
			3'b010:
				// Trace: design.sv:53236:23
				round_up = (|round_sticky_bits_i ? sign_i : 1'b0);
			3'b011:
				// Trace: design.sv:53237:23
				round_up = (|round_sticky_bits_i ? ~sign_i : 1'b0);
			3'b100:
				// Trace: design.sv:53238:23
				round_up = round_sticky_bits_i[1];
			default:
				// Trace: design.sv:53239:16
				round_up = fpnew_pkg_DONT_CARE;
		endcase
	end
	// Trace: design.sv:53244:3
	assign abs_rounded_o = abs_value_i + round_up;
	// Trace: design.sv:53247:3
	assign exact_zero_o = (abs_value_i == {AbsWidth {1'sb0}}) && (round_sticky_bits_i == {2 {1'sb0}});
	// Trace: design.sv:53251:3
	assign sign_o = (exact_zero_o && effective_subtraction_i ? rnd_mode_i == 3'b010 : sign_i);
	initial _sv2v_0 = 0;
endmodule
module fpnew_top (
	clk_i,
	rst_ni,
	operands_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	reg _sv2v_0;
	// Trace: design.sv:53273:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	// removed localparam type fpnew_pkg_fpu_features_t
	localparam [42:0] fpnew_pkg_RV64D_Xsflt = 43'h000000207ff;
	parameter [42:0] Features = fpnew_pkg_RV64D_Xsflt;
	// Trace: design.sv:53274:13
	// removed localparam type fpnew_pkg_pipe_config_t
	// removed localparam type fpnew_pkg_unit_type_t
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unit_types_t
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unsigned_t
	// removed localparam type fpnew_pkg_fpu_implementation_t
	function automatic [159:0] sv2v_cast_C3475;
		input reg [159:0] inp;
		sv2v_cast_C3475 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_52F10;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_52F10 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_18D94;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_18D94 = inp;
	endfunction
	localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] fpnew_pkg_DEFAULT_NOREGS = {sv2v_cast_52F10({fpnew_pkg_NUM_OPGROUPS {sv2v_cast_C3475(0)}}), sv2v_cast_18D94({{fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}, {fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}}), 2'd0};
	parameter [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] Implementation = fpnew_pkg_DEFAULT_NOREGS;
	// Trace: design.sv:53275:45
	// removed localparam type TagType
	// Trace: design.sv:53277:14
	localparam [31:0] WIDTH = Features[42-:32];
	// Trace: design.sv:53278:14
	localparam [31:0] NUM_OPERANDS = 3;
	// Trace: design.sv:53280:3
	input wire clk_i;
	// Trace: design.sv:53281:3
	input wire rst_ni;
	// Trace: design.sv:53283:3
	input wire [(NUM_OPERANDS * WIDTH) - 1:0] operands_i;
	// Trace: design.sv:53284:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: design.sv:53285:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: design.sv:53286:3
	input wire op_mod_i;
	// Trace: design.sv:53287:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: design.sv:53288:3
	input wire [2:0] dst_fmt_i;
	// Trace: design.sv:53289:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: design.sv:53290:3
	input wire vectorial_op_i;
	// Trace: design.sv:53291:3
	input wire tag_i;
	// Trace: design.sv:53293:3
	input wire in_valid_i;
	// Trace: design.sv:53294:3
	output wire in_ready_o;
	// Trace: design.sv:53295:3
	input wire flush_i;
	// Trace: design.sv:53297:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: design.sv:53298:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: design.sv:53299:3
	output wire tag_o;
	// Trace: design.sv:53301:3
	output wire out_valid_o;
	// Trace: design.sv:53302:3
	input wire out_ready_i;
	// Trace: design.sv:53304:3
	output wire busy_o;
	// Trace: design.sv:53307:3
	localparam [31:0] NUM_OPGROUPS = fpnew_pkg_NUM_OPGROUPS;
	// Trace: design.sv:53308:3
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: design.sv:53313:3
	// removed localparam type output_t
	// Trace: design.sv:53320:3
	wire [3:0] opgrp_in_ready;
	wire [3:0] opgrp_out_valid;
	wire [3:0] opgrp_out_ready;
	wire [3:0] opgrp_ext;
	wire [3:0] opgrp_busy;
	// Trace: design.sv:53321:3
	wire [((WIDTH + 5) >= 0 ? (4 * (WIDTH + 6)) - 1 : (4 * (1 - (WIDTH + 5))) + (WIDTH + 4)):((WIDTH + 5) >= 0 ? 0 : WIDTH + 5)] opgrp_outputs;
	// Trace: design.sv:53323:3
	wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed;
	// Trace: design.sv:53328:3
	// removed localparam type fpnew_pkg_opgroup_e
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	function automatic [1:0] fpnew_pkg_get_opgroup;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:367:44
		input reg [3:0] op;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:368:5
		(* full_case, parallel_case *)
		case (op)
			sv2v_cast_4CD2E(0), sv2v_cast_4CD2E(1), sv2v_cast_4CD2E(2), sv2v_cast_4CD2E(3): fpnew_pkg_get_opgroup = 2'd0;
			sv2v_cast_4CD2E(4), sv2v_cast_4CD2E(5): fpnew_pkg_get_opgroup = 2'd1;
			sv2v_cast_4CD2E(6), sv2v_cast_4CD2E(7), sv2v_cast_4CD2E(8), sv2v_cast_4CD2E(9): fpnew_pkg_get_opgroup = 2'd2;
			sv2v_cast_4CD2E(10), sv2v_cast_4CD2E(11), sv2v_cast_4CD2E(12), sv2v_cast_4CD2E(13), sv2v_cast_4CD2E(14): fpnew_pkg_get_opgroup = 2'd3;
			default: fpnew_pkg_get_opgroup = 2'd2;
		endcase
	endfunction
	assign in_ready_o = in_valid_i & opgrp_in_ready[fpnew_pkg_get_opgroup(op_i)];
	// Trace: design.sv:53331:3
	genvar _gv_fmt_12;
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:303:44
		input reg [2:0] fmt;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:304:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_fmt_12 = 0; _gv_fmt_12 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_12 = _gv_fmt_12 + 1) begin : gen_nanbox_check
			localparam fmt = _gv_fmt_12;
			// Trace: design.sv:53332:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			if (Features[9] && (FP_WIDTH < WIDTH)) begin : check
				genvar _gv_op_3;
				for (_gv_op_3 = 0; _gv_op_3 < sv2v_cast_32_signed(NUM_OPERANDS); _gv_op_3 = _gv_op_3 + 1) begin : operands
					localparam op = _gv_op_3;
					// Trace: design.sv:53336:9
					assign is_boxed[(fmt * NUM_OPERANDS) + op] = (!vectorial_op_i ? operands_i[(op * WIDTH) + ((WIDTH - 1) >= FP_WIDTH ? WIDTH - 1 : ((WIDTH - 1) + ((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)) - 1)-:((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)] == {((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1) * 1 {1'sb1}} : 1'b1);
				end
			end
			else begin : no_check
				// Trace: design.sv:53341:7
				assign is_boxed[fmt * NUM_OPERANDS+:NUM_OPERANDS] = 1'sb1;
			end
		end
	endgenerate
	// Trace: design.sv:53348:3
	genvar _gv_opgrp_1;
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:378:48
		input reg [1:0] grp;
		// Trace: ../src/pulp-platform.org_ip_fpnew_0/pulp_platform_fpnew/src/fpnew_pkg.sv:379:5
		(* full_case, parallel_case *)
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		for (_gv_opgrp_1 = 0; _gv_opgrp_1 < sv2v_cast_32_signed(NUM_OPGROUPS); _gv_opgrp_1 = _gv_opgrp_1 + 1) begin : gen_operation_groups
			localparam opgrp = _gv_opgrp_1;
			// Trace: design.sv:53349:5
			localparam [31:0] NUM_OPS = fpnew_pkg_num_operands(sv2v_cast_2(opgrp));
			// Trace: design.sv:53351:5
			wire in_valid;
			// Trace: design.sv:53352:5
			reg [(NUM_FORMATS * NUM_OPS) - 1:0] input_boxed;
			// Trace: design.sv:53354:5
			assign in_valid = in_valid_i & (fpnew_pkg_get_opgroup(op_i) == sv2v_cast_2(opgrp));
			// Trace: design.sv:53357:5
			always @(*) begin : slice_inputs
				if (_sv2v_0)
					;
				// Trace: design.sv:53358:7
				begin : sv2v_autoblock_1
					// Trace: design.sv:53358:12
					reg [31:0] fmt;
					// Trace: design.sv:53358:12
					for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
						begin
							// Trace: design.sv:53359:9
							input_boxed[fmt * fpnew_pkg_num_operands(sv2v_cast_2(_gv_opgrp_1))+:fpnew_pkg_num_operands(sv2v_cast_2(_gv_opgrp_1))] = is_boxed[(fmt * NUM_OPERANDS) + (NUM_OPS - 1)-:NUM_OPS];
						end
				end
			end
			// Trace: design.sv:53362:5
			fpnew_opgroup_block_37AAD #(
				.OpGroup(sv2v_cast_2(opgrp)),
				.Width(WIDTH),
				.EnableVectors(Features[10]),
				.FpFmtMask(Features[8-:5]),
				.IntFmtMask(Features[3-:fpnew_pkg_NUM_INT_FORMATS]),
				.FmtPipeRegs(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + (((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1)) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) - 1) - (32 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:160]),
				.FmtUnitTypes(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) - 1) - (2 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:10]),
				.PipeConfig(Implementation[1-:2])
			) i_opgroup_block(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i[WIDTH * ((NUM_OPS - 1) - (NUM_OPS - 1))+:WIDTH * NUM_OPS]),
				.is_boxed_i(input_boxed),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.in_valid_i(in_valid),
				.in_ready_o(opgrp_in_ready[opgrp]),
				.flush_i(flush_i),
				.result_o(opgrp_outputs[((WIDTH + 5) >= 0 ? (opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? WIDTH + 5 : (WIDTH + 5) - (WIDTH + 5)) : (((opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? WIDTH + 5 : (WIDTH + 5) - (WIDTH + 5))) + ((WIDTH + 5) >= 6 ? WIDTH + 0 : 7 - (WIDTH + 5))) - 1)-:((WIDTH + 5) >= 6 ? WIDTH + 0 : 7 - (WIDTH + 5))]),
				.status_o(opgrp_outputs[((WIDTH + 5) >= 0 ? (opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? 5 : WIDTH + 0) : ((opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? 5 : WIDTH + 0)) + 4)-:5]),
				.extension_bit_o(opgrp_ext[opgrp]),
				.tag_o(opgrp_outputs[(opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? 0 : WIDTH + 5)]),
				.out_valid_o(opgrp_out_valid[opgrp]),
				.out_ready_i(opgrp_out_ready[opgrp]),
				.busy_o(opgrp_busy[opgrp])
			);
		end
	endgenerate
	// Trace: design.sv:53401:3
	wire [WIDTH + 5:0] arbiter_output;
	// Trace: design.sv:53404:3
	localparam [31:0] sv2v_uu_i_arbiter_NumIn = NUM_OPGROUPS;
	localparam [31:0] sv2v_uu_i_arbiter_IdxWidth = $unsigned(2);
	// removed localparam type sv2v_uu_i_arbiter_rr_i
	localparam [sv2v_uu_i_arbiter_IdxWidth - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_A5EF3_DDD71 #(
		.DataType_WIDTH(WIDTH),
		.NumIn(NUM_OPGROUPS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
		.req_i(opgrp_out_valid),
		.gnt_o(opgrp_out_ready),
		.data_i(opgrp_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: design.sv:53423:3
	assign result_o = arbiter_output[WIDTH + 5-:((WIDTH + 5) >= 6 ? WIDTH + 0 : 7 - (WIDTH + 5))];
	// Trace: design.sv:53424:3
	assign status_o = arbiter_output[5-:5];
	// Trace: design.sv:53425:3
	assign tag_o = arbiter_output[0];
	// Trace: design.sv:53427:3
	assign busy_o = |opgrp_busy;
	initial _sv2v_0 = 0;
endmodule
// removed package "gpio_reg_pkg"
module gpio_reg_top_04165 (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	reg2hw,
	hw2reg,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:53686:20
	// removed localparam type reg_req_t
	// Trace: design.sv:53687:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:53688:15
	parameter signed [31:0] AW = 11;
	// Trace: design.sv:53690:3
	input clk_i;
	// Trace: design.sv:53691:3
	input rst_ni;
	// Trace: design.sv:53692:3
	input wire [69:0] reg_req_i;
	// Trace: design.sv:53693:3
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:53695:3
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_cfg_reg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_clear_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_mode_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_out_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_set_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_toggle_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_fall_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_fall_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_lvl_high_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_lvl_high_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_lvl_low_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_lvl_low_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_rise_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_rise_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_t
	output wire [642:0] reg2hw;
	// Trace: design.sv:53696:3
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_gpio_in_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_gpio_out_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_info_reg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_fall_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_lvl_high_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_lvl_low_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_rise_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_t
	input wire [403:0] hw2reg;
	// Trace: design.sv:53700:3
	input devmode_i;
	// Trace: design.sv:53703:3
	// removed import gpio_reg_pkg::*;
	// Trace: design.sv:53705:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:53706:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:53709:3
	wire reg_we;
	// Trace: design.sv:53710:3
	wire reg_re;
	// Trace: design.sv:53711:3
	wire [AW - 1:0] reg_addr;
	// Trace: design.sv:53712:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:53713:3
	wire [3:0] reg_be;
	// Trace: design.sv:53714:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:53715:3
	wire reg_error;
	// Trace: design.sv:53717:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:53719:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:53722:3
	wire [69:0] reg_intf_req;
	// Trace: design.sv:53723:3
	wire [33:0] reg_intf_rsp;
	// Trace: design.sv:53726:3
	assign reg_intf_req = reg_req_i;
	// Trace: design.sv:53727:3
	assign reg_rsp_o = reg_intf_rsp;
	// Trace: design.sv:53730:3
	assign reg_we = reg_intf_req[69] & reg_intf_req[68];
	// Trace: design.sv:53731:3
	assign reg_re = reg_intf_req[69] & ~reg_intf_req[68];
	// Trace: design.sv:53732:3
	assign reg_addr = reg_intf_req[63-:32];
	// Trace: design.sv:53733:3
	assign reg_wdata = reg_intf_req[31-:32];
	// Trace: design.sv:53734:3
	assign reg_be = reg_intf_req[67-:4];
	// Trace: design.sv:53735:3
	assign reg_intf_rsp[31-:32] = reg_rdata;
	// Trace: design.sv:53736:3
	assign reg_intf_rsp[33] = reg_error;
	// Trace: design.sv:53737:3
	assign reg_intf_rsp[32] = 1'b1;
	// Trace: design.sv:53739:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:53740:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:53746:3
	wire [9:0] info_gpio_cnt_qs;
	// Trace: design.sv:53747:3
	wire info_gpio_cnt_re;
	// Trace: design.sv:53748:3
	wire [9:0] info_version_qs;
	// Trace: design.sv:53749:3
	wire info_version_re;
	// Trace: design.sv:53750:3
	wire cfg_glbl_intrpt_mode_qs;
	// Trace: design.sv:53751:3
	wire cfg_glbl_intrpt_mode_wd;
	// Trace: design.sv:53752:3
	wire cfg_glbl_intrpt_mode_we;
	// Trace: design.sv:53753:3
	wire cfg_pin_lvl_intrpt_mode_qs;
	// Trace: design.sv:53754:3
	wire cfg_pin_lvl_intrpt_mode_wd;
	// Trace: design.sv:53755:3
	wire cfg_pin_lvl_intrpt_mode_we;
	// Trace: design.sv:53756:3
	wire cfg_reserved_qs;
	// Trace: design.sv:53757:3
	wire cfg_reserved_wd;
	// Trace: design.sv:53758:3
	wire cfg_reserved_we;
	// Trace: design.sv:53759:3
	wire [1:0] gpio_mode_0_mode_0_qs;
	// Trace: design.sv:53760:3
	wire [1:0] gpio_mode_0_mode_0_wd;
	// Trace: design.sv:53761:3
	wire gpio_mode_0_mode_0_we;
	// Trace: design.sv:53762:3
	wire [1:0] gpio_mode_0_mode_1_qs;
	// Trace: design.sv:53763:3
	wire [1:0] gpio_mode_0_mode_1_wd;
	// Trace: design.sv:53764:3
	wire gpio_mode_0_mode_1_we;
	// Trace: design.sv:53765:3
	wire [1:0] gpio_mode_0_mode_2_qs;
	// Trace: design.sv:53766:3
	wire [1:0] gpio_mode_0_mode_2_wd;
	// Trace: design.sv:53767:3
	wire gpio_mode_0_mode_2_we;
	// Trace: design.sv:53768:3
	wire [1:0] gpio_mode_0_mode_3_qs;
	// Trace: design.sv:53769:3
	wire [1:0] gpio_mode_0_mode_3_wd;
	// Trace: design.sv:53770:3
	wire gpio_mode_0_mode_3_we;
	// Trace: design.sv:53771:3
	wire [1:0] gpio_mode_0_mode_4_qs;
	// Trace: design.sv:53772:3
	wire [1:0] gpio_mode_0_mode_4_wd;
	// Trace: design.sv:53773:3
	wire gpio_mode_0_mode_4_we;
	// Trace: design.sv:53774:3
	wire [1:0] gpio_mode_0_mode_5_qs;
	// Trace: design.sv:53775:3
	wire [1:0] gpio_mode_0_mode_5_wd;
	// Trace: design.sv:53776:3
	wire gpio_mode_0_mode_5_we;
	// Trace: design.sv:53777:3
	wire [1:0] gpio_mode_0_mode_6_qs;
	// Trace: design.sv:53778:3
	wire [1:0] gpio_mode_0_mode_6_wd;
	// Trace: design.sv:53779:3
	wire gpio_mode_0_mode_6_we;
	// Trace: design.sv:53780:3
	wire [1:0] gpio_mode_0_mode_7_qs;
	// Trace: design.sv:53781:3
	wire [1:0] gpio_mode_0_mode_7_wd;
	// Trace: design.sv:53782:3
	wire gpio_mode_0_mode_7_we;
	// Trace: design.sv:53783:3
	wire [1:0] gpio_mode_0_mode_8_qs;
	// Trace: design.sv:53784:3
	wire [1:0] gpio_mode_0_mode_8_wd;
	// Trace: design.sv:53785:3
	wire gpio_mode_0_mode_8_we;
	// Trace: design.sv:53786:3
	wire [1:0] gpio_mode_0_mode_9_qs;
	// Trace: design.sv:53787:3
	wire [1:0] gpio_mode_0_mode_9_wd;
	// Trace: design.sv:53788:3
	wire gpio_mode_0_mode_9_we;
	// Trace: design.sv:53789:3
	wire [1:0] gpio_mode_0_mode_10_qs;
	// Trace: design.sv:53790:3
	wire [1:0] gpio_mode_0_mode_10_wd;
	// Trace: design.sv:53791:3
	wire gpio_mode_0_mode_10_we;
	// Trace: design.sv:53792:3
	wire [1:0] gpio_mode_0_mode_11_qs;
	// Trace: design.sv:53793:3
	wire [1:0] gpio_mode_0_mode_11_wd;
	// Trace: design.sv:53794:3
	wire gpio_mode_0_mode_11_we;
	// Trace: design.sv:53795:3
	wire [1:0] gpio_mode_0_mode_12_qs;
	// Trace: design.sv:53796:3
	wire [1:0] gpio_mode_0_mode_12_wd;
	// Trace: design.sv:53797:3
	wire gpio_mode_0_mode_12_we;
	// Trace: design.sv:53798:3
	wire [1:0] gpio_mode_0_mode_13_qs;
	// Trace: design.sv:53799:3
	wire [1:0] gpio_mode_0_mode_13_wd;
	// Trace: design.sv:53800:3
	wire gpio_mode_0_mode_13_we;
	// Trace: design.sv:53801:3
	wire [1:0] gpio_mode_0_mode_14_qs;
	// Trace: design.sv:53802:3
	wire [1:0] gpio_mode_0_mode_14_wd;
	// Trace: design.sv:53803:3
	wire gpio_mode_0_mode_14_we;
	// Trace: design.sv:53804:3
	wire [1:0] gpio_mode_0_mode_15_qs;
	// Trace: design.sv:53805:3
	wire [1:0] gpio_mode_0_mode_15_wd;
	// Trace: design.sv:53806:3
	wire gpio_mode_0_mode_15_we;
	// Trace: design.sv:53807:3
	wire [1:0] gpio_mode_1_mode_16_qs;
	// Trace: design.sv:53808:3
	wire [1:0] gpio_mode_1_mode_16_wd;
	// Trace: design.sv:53809:3
	wire gpio_mode_1_mode_16_we;
	// Trace: design.sv:53810:3
	wire [1:0] gpio_mode_1_mode_17_qs;
	// Trace: design.sv:53811:3
	wire [1:0] gpio_mode_1_mode_17_wd;
	// Trace: design.sv:53812:3
	wire gpio_mode_1_mode_17_we;
	// Trace: design.sv:53813:3
	wire [1:0] gpio_mode_1_mode_18_qs;
	// Trace: design.sv:53814:3
	wire [1:0] gpio_mode_1_mode_18_wd;
	// Trace: design.sv:53815:3
	wire gpio_mode_1_mode_18_we;
	// Trace: design.sv:53816:3
	wire [1:0] gpio_mode_1_mode_19_qs;
	// Trace: design.sv:53817:3
	wire [1:0] gpio_mode_1_mode_19_wd;
	// Trace: design.sv:53818:3
	wire gpio_mode_1_mode_19_we;
	// Trace: design.sv:53819:3
	wire [1:0] gpio_mode_1_mode_20_qs;
	// Trace: design.sv:53820:3
	wire [1:0] gpio_mode_1_mode_20_wd;
	// Trace: design.sv:53821:3
	wire gpio_mode_1_mode_20_we;
	// Trace: design.sv:53822:3
	wire [1:0] gpio_mode_1_mode_21_qs;
	// Trace: design.sv:53823:3
	wire [1:0] gpio_mode_1_mode_21_wd;
	// Trace: design.sv:53824:3
	wire gpio_mode_1_mode_21_we;
	// Trace: design.sv:53825:3
	wire [1:0] gpio_mode_1_mode_22_qs;
	// Trace: design.sv:53826:3
	wire [1:0] gpio_mode_1_mode_22_wd;
	// Trace: design.sv:53827:3
	wire gpio_mode_1_mode_22_we;
	// Trace: design.sv:53828:3
	wire [1:0] gpio_mode_1_mode_23_qs;
	// Trace: design.sv:53829:3
	wire [1:0] gpio_mode_1_mode_23_wd;
	// Trace: design.sv:53830:3
	wire gpio_mode_1_mode_23_we;
	// Trace: design.sv:53831:3
	wire [1:0] gpio_mode_1_mode_24_qs;
	// Trace: design.sv:53832:3
	wire [1:0] gpio_mode_1_mode_24_wd;
	// Trace: design.sv:53833:3
	wire gpio_mode_1_mode_24_we;
	// Trace: design.sv:53834:3
	wire [1:0] gpio_mode_1_mode_25_qs;
	// Trace: design.sv:53835:3
	wire [1:0] gpio_mode_1_mode_25_wd;
	// Trace: design.sv:53836:3
	wire gpio_mode_1_mode_25_we;
	// Trace: design.sv:53837:3
	wire [1:0] gpio_mode_1_mode_26_qs;
	// Trace: design.sv:53838:3
	wire [1:0] gpio_mode_1_mode_26_wd;
	// Trace: design.sv:53839:3
	wire gpio_mode_1_mode_26_we;
	// Trace: design.sv:53840:3
	wire [1:0] gpio_mode_1_mode_27_qs;
	// Trace: design.sv:53841:3
	wire [1:0] gpio_mode_1_mode_27_wd;
	// Trace: design.sv:53842:3
	wire gpio_mode_1_mode_27_we;
	// Trace: design.sv:53843:3
	wire [1:0] gpio_mode_1_mode_28_qs;
	// Trace: design.sv:53844:3
	wire [1:0] gpio_mode_1_mode_28_wd;
	// Trace: design.sv:53845:3
	wire gpio_mode_1_mode_28_we;
	// Trace: design.sv:53846:3
	wire [1:0] gpio_mode_1_mode_29_qs;
	// Trace: design.sv:53847:3
	wire [1:0] gpio_mode_1_mode_29_wd;
	// Trace: design.sv:53848:3
	wire gpio_mode_1_mode_29_we;
	// Trace: design.sv:53849:3
	wire [1:0] gpio_mode_1_mode_30_qs;
	// Trace: design.sv:53850:3
	wire [1:0] gpio_mode_1_mode_30_wd;
	// Trace: design.sv:53851:3
	wire gpio_mode_1_mode_30_we;
	// Trace: design.sv:53852:3
	wire [1:0] gpio_mode_1_mode_31_qs;
	// Trace: design.sv:53853:3
	wire [1:0] gpio_mode_1_mode_31_wd;
	// Trace: design.sv:53854:3
	wire gpio_mode_1_mode_31_we;
	// Trace: design.sv:53855:3
	wire gpio_en_gpio_en_0_qs;
	// Trace: design.sv:53856:3
	wire gpio_en_gpio_en_0_wd;
	// Trace: design.sv:53857:3
	wire gpio_en_gpio_en_0_we;
	// Trace: design.sv:53858:3
	wire gpio_en_gpio_en_1_qs;
	// Trace: design.sv:53859:3
	wire gpio_en_gpio_en_1_wd;
	// Trace: design.sv:53860:3
	wire gpio_en_gpio_en_1_we;
	// Trace: design.sv:53861:3
	wire gpio_en_gpio_en_2_qs;
	// Trace: design.sv:53862:3
	wire gpio_en_gpio_en_2_wd;
	// Trace: design.sv:53863:3
	wire gpio_en_gpio_en_2_we;
	// Trace: design.sv:53864:3
	wire gpio_en_gpio_en_3_qs;
	// Trace: design.sv:53865:3
	wire gpio_en_gpio_en_3_wd;
	// Trace: design.sv:53866:3
	wire gpio_en_gpio_en_3_we;
	// Trace: design.sv:53867:3
	wire gpio_en_gpio_en_4_qs;
	// Trace: design.sv:53868:3
	wire gpio_en_gpio_en_4_wd;
	// Trace: design.sv:53869:3
	wire gpio_en_gpio_en_4_we;
	// Trace: design.sv:53870:3
	wire gpio_en_gpio_en_5_qs;
	// Trace: design.sv:53871:3
	wire gpio_en_gpio_en_5_wd;
	// Trace: design.sv:53872:3
	wire gpio_en_gpio_en_5_we;
	// Trace: design.sv:53873:3
	wire gpio_en_gpio_en_6_qs;
	// Trace: design.sv:53874:3
	wire gpio_en_gpio_en_6_wd;
	// Trace: design.sv:53875:3
	wire gpio_en_gpio_en_6_we;
	// Trace: design.sv:53876:3
	wire gpio_en_gpio_en_7_qs;
	// Trace: design.sv:53877:3
	wire gpio_en_gpio_en_7_wd;
	// Trace: design.sv:53878:3
	wire gpio_en_gpio_en_7_we;
	// Trace: design.sv:53879:3
	wire gpio_en_gpio_en_8_qs;
	// Trace: design.sv:53880:3
	wire gpio_en_gpio_en_8_wd;
	// Trace: design.sv:53881:3
	wire gpio_en_gpio_en_8_we;
	// Trace: design.sv:53882:3
	wire gpio_en_gpio_en_9_qs;
	// Trace: design.sv:53883:3
	wire gpio_en_gpio_en_9_wd;
	// Trace: design.sv:53884:3
	wire gpio_en_gpio_en_9_we;
	// Trace: design.sv:53885:3
	wire gpio_en_gpio_en_10_qs;
	// Trace: design.sv:53886:3
	wire gpio_en_gpio_en_10_wd;
	// Trace: design.sv:53887:3
	wire gpio_en_gpio_en_10_we;
	// Trace: design.sv:53888:3
	wire gpio_en_gpio_en_11_qs;
	// Trace: design.sv:53889:3
	wire gpio_en_gpio_en_11_wd;
	// Trace: design.sv:53890:3
	wire gpio_en_gpio_en_11_we;
	// Trace: design.sv:53891:3
	wire gpio_en_gpio_en_12_qs;
	// Trace: design.sv:53892:3
	wire gpio_en_gpio_en_12_wd;
	// Trace: design.sv:53893:3
	wire gpio_en_gpio_en_12_we;
	// Trace: design.sv:53894:3
	wire gpio_en_gpio_en_13_qs;
	// Trace: design.sv:53895:3
	wire gpio_en_gpio_en_13_wd;
	// Trace: design.sv:53896:3
	wire gpio_en_gpio_en_13_we;
	// Trace: design.sv:53897:3
	wire gpio_en_gpio_en_14_qs;
	// Trace: design.sv:53898:3
	wire gpio_en_gpio_en_14_wd;
	// Trace: design.sv:53899:3
	wire gpio_en_gpio_en_14_we;
	// Trace: design.sv:53900:3
	wire gpio_en_gpio_en_15_qs;
	// Trace: design.sv:53901:3
	wire gpio_en_gpio_en_15_wd;
	// Trace: design.sv:53902:3
	wire gpio_en_gpio_en_15_we;
	// Trace: design.sv:53903:3
	wire gpio_en_gpio_en_16_qs;
	// Trace: design.sv:53904:3
	wire gpio_en_gpio_en_16_wd;
	// Trace: design.sv:53905:3
	wire gpio_en_gpio_en_16_we;
	// Trace: design.sv:53906:3
	wire gpio_en_gpio_en_17_qs;
	// Trace: design.sv:53907:3
	wire gpio_en_gpio_en_17_wd;
	// Trace: design.sv:53908:3
	wire gpio_en_gpio_en_17_we;
	// Trace: design.sv:53909:3
	wire gpio_en_gpio_en_18_qs;
	// Trace: design.sv:53910:3
	wire gpio_en_gpio_en_18_wd;
	// Trace: design.sv:53911:3
	wire gpio_en_gpio_en_18_we;
	// Trace: design.sv:53912:3
	wire gpio_en_gpio_en_19_qs;
	// Trace: design.sv:53913:3
	wire gpio_en_gpio_en_19_wd;
	// Trace: design.sv:53914:3
	wire gpio_en_gpio_en_19_we;
	// Trace: design.sv:53915:3
	wire gpio_en_gpio_en_20_qs;
	// Trace: design.sv:53916:3
	wire gpio_en_gpio_en_20_wd;
	// Trace: design.sv:53917:3
	wire gpio_en_gpio_en_20_we;
	// Trace: design.sv:53918:3
	wire gpio_en_gpio_en_21_qs;
	// Trace: design.sv:53919:3
	wire gpio_en_gpio_en_21_wd;
	// Trace: design.sv:53920:3
	wire gpio_en_gpio_en_21_we;
	// Trace: design.sv:53921:3
	wire gpio_en_gpio_en_22_qs;
	// Trace: design.sv:53922:3
	wire gpio_en_gpio_en_22_wd;
	// Trace: design.sv:53923:3
	wire gpio_en_gpio_en_22_we;
	// Trace: design.sv:53924:3
	wire gpio_en_gpio_en_23_qs;
	// Trace: design.sv:53925:3
	wire gpio_en_gpio_en_23_wd;
	// Trace: design.sv:53926:3
	wire gpio_en_gpio_en_23_we;
	// Trace: design.sv:53927:3
	wire gpio_en_gpio_en_24_qs;
	// Trace: design.sv:53928:3
	wire gpio_en_gpio_en_24_wd;
	// Trace: design.sv:53929:3
	wire gpio_en_gpio_en_24_we;
	// Trace: design.sv:53930:3
	wire gpio_en_gpio_en_25_qs;
	// Trace: design.sv:53931:3
	wire gpio_en_gpio_en_25_wd;
	// Trace: design.sv:53932:3
	wire gpio_en_gpio_en_25_we;
	// Trace: design.sv:53933:3
	wire gpio_en_gpio_en_26_qs;
	// Trace: design.sv:53934:3
	wire gpio_en_gpio_en_26_wd;
	// Trace: design.sv:53935:3
	wire gpio_en_gpio_en_26_we;
	// Trace: design.sv:53936:3
	wire gpio_en_gpio_en_27_qs;
	// Trace: design.sv:53937:3
	wire gpio_en_gpio_en_27_wd;
	// Trace: design.sv:53938:3
	wire gpio_en_gpio_en_27_we;
	// Trace: design.sv:53939:3
	wire gpio_en_gpio_en_28_qs;
	// Trace: design.sv:53940:3
	wire gpio_en_gpio_en_28_wd;
	// Trace: design.sv:53941:3
	wire gpio_en_gpio_en_28_we;
	// Trace: design.sv:53942:3
	wire gpio_en_gpio_en_29_qs;
	// Trace: design.sv:53943:3
	wire gpio_en_gpio_en_29_wd;
	// Trace: design.sv:53944:3
	wire gpio_en_gpio_en_29_we;
	// Trace: design.sv:53945:3
	wire gpio_en_gpio_en_30_qs;
	// Trace: design.sv:53946:3
	wire gpio_en_gpio_en_30_wd;
	// Trace: design.sv:53947:3
	wire gpio_en_gpio_en_30_we;
	// Trace: design.sv:53948:3
	wire gpio_en_gpio_en_31_qs;
	// Trace: design.sv:53949:3
	wire gpio_en_gpio_en_31_wd;
	// Trace: design.sv:53950:3
	wire gpio_en_gpio_en_31_we;
	// Trace: design.sv:53951:3
	wire gpio_in_gpio_in_0_qs;
	// Trace: design.sv:53952:3
	wire gpio_in_gpio_in_0_re;
	// Trace: design.sv:53953:3
	wire gpio_in_gpio_in_1_qs;
	// Trace: design.sv:53954:3
	wire gpio_in_gpio_in_1_re;
	// Trace: design.sv:53955:3
	wire gpio_in_gpio_in_2_qs;
	// Trace: design.sv:53956:3
	wire gpio_in_gpio_in_2_re;
	// Trace: design.sv:53957:3
	wire gpio_in_gpio_in_3_qs;
	// Trace: design.sv:53958:3
	wire gpio_in_gpio_in_3_re;
	// Trace: design.sv:53959:3
	wire gpio_in_gpio_in_4_qs;
	// Trace: design.sv:53960:3
	wire gpio_in_gpio_in_4_re;
	// Trace: design.sv:53961:3
	wire gpio_in_gpio_in_5_qs;
	// Trace: design.sv:53962:3
	wire gpio_in_gpio_in_5_re;
	// Trace: design.sv:53963:3
	wire gpio_in_gpio_in_6_qs;
	// Trace: design.sv:53964:3
	wire gpio_in_gpio_in_6_re;
	// Trace: design.sv:53965:3
	wire gpio_in_gpio_in_7_qs;
	// Trace: design.sv:53966:3
	wire gpio_in_gpio_in_7_re;
	// Trace: design.sv:53967:3
	wire gpio_in_gpio_in_8_qs;
	// Trace: design.sv:53968:3
	wire gpio_in_gpio_in_8_re;
	// Trace: design.sv:53969:3
	wire gpio_in_gpio_in_9_qs;
	// Trace: design.sv:53970:3
	wire gpio_in_gpio_in_9_re;
	// Trace: design.sv:53971:3
	wire gpio_in_gpio_in_10_qs;
	// Trace: design.sv:53972:3
	wire gpio_in_gpio_in_10_re;
	// Trace: design.sv:53973:3
	wire gpio_in_gpio_in_11_qs;
	// Trace: design.sv:53974:3
	wire gpio_in_gpio_in_11_re;
	// Trace: design.sv:53975:3
	wire gpio_in_gpio_in_12_qs;
	// Trace: design.sv:53976:3
	wire gpio_in_gpio_in_12_re;
	// Trace: design.sv:53977:3
	wire gpio_in_gpio_in_13_qs;
	// Trace: design.sv:53978:3
	wire gpio_in_gpio_in_13_re;
	// Trace: design.sv:53979:3
	wire gpio_in_gpio_in_14_qs;
	// Trace: design.sv:53980:3
	wire gpio_in_gpio_in_14_re;
	// Trace: design.sv:53981:3
	wire gpio_in_gpio_in_15_qs;
	// Trace: design.sv:53982:3
	wire gpio_in_gpio_in_15_re;
	// Trace: design.sv:53983:3
	wire gpio_in_gpio_in_16_qs;
	// Trace: design.sv:53984:3
	wire gpio_in_gpio_in_16_re;
	// Trace: design.sv:53985:3
	wire gpio_in_gpio_in_17_qs;
	// Trace: design.sv:53986:3
	wire gpio_in_gpio_in_17_re;
	// Trace: design.sv:53987:3
	wire gpio_in_gpio_in_18_qs;
	// Trace: design.sv:53988:3
	wire gpio_in_gpio_in_18_re;
	// Trace: design.sv:53989:3
	wire gpio_in_gpio_in_19_qs;
	// Trace: design.sv:53990:3
	wire gpio_in_gpio_in_19_re;
	// Trace: design.sv:53991:3
	wire gpio_in_gpio_in_20_qs;
	// Trace: design.sv:53992:3
	wire gpio_in_gpio_in_20_re;
	// Trace: design.sv:53993:3
	wire gpio_in_gpio_in_21_qs;
	// Trace: design.sv:53994:3
	wire gpio_in_gpio_in_21_re;
	// Trace: design.sv:53995:3
	wire gpio_in_gpio_in_22_qs;
	// Trace: design.sv:53996:3
	wire gpio_in_gpio_in_22_re;
	// Trace: design.sv:53997:3
	wire gpio_in_gpio_in_23_qs;
	// Trace: design.sv:53998:3
	wire gpio_in_gpio_in_23_re;
	// Trace: design.sv:53999:3
	wire gpio_in_gpio_in_24_qs;
	// Trace: design.sv:54000:3
	wire gpio_in_gpio_in_24_re;
	// Trace: design.sv:54001:3
	wire gpio_in_gpio_in_25_qs;
	// Trace: design.sv:54002:3
	wire gpio_in_gpio_in_25_re;
	// Trace: design.sv:54003:3
	wire gpio_in_gpio_in_26_qs;
	// Trace: design.sv:54004:3
	wire gpio_in_gpio_in_26_re;
	// Trace: design.sv:54005:3
	wire gpio_in_gpio_in_27_qs;
	// Trace: design.sv:54006:3
	wire gpio_in_gpio_in_27_re;
	// Trace: design.sv:54007:3
	wire gpio_in_gpio_in_28_qs;
	// Trace: design.sv:54008:3
	wire gpio_in_gpio_in_28_re;
	// Trace: design.sv:54009:3
	wire gpio_in_gpio_in_29_qs;
	// Trace: design.sv:54010:3
	wire gpio_in_gpio_in_29_re;
	// Trace: design.sv:54011:3
	wire gpio_in_gpio_in_30_qs;
	// Trace: design.sv:54012:3
	wire gpio_in_gpio_in_30_re;
	// Trace: design.sv:54013:3
	wire gpio_in_gpio_in_31_qs;
	// Trace: design.sv:54014:3
	wire gpio_in_gpio_in_31_re;
	// Trace: design.sv:54015:3
	wire gpio_out_gpio_out_0_qs;
	// Trace: design.sv:54016:3
	wire gpio_out_gpio_out_0_wd;
	// Trace: design.sv:54017:3
	wire gpio_out_gpio_out_0_we;
	// Trace: design.sv:54018:3
	wire gpio_out_gpio_out_1_qs;
	// Trace: design.sv:54019:3
	wire gpio_out_gpio_out_1_wd;
	// Trace: design.sv:54020:3
	wire gpio_out_gpio_out_1_we;
	// Trace: design.sv:54021:3
	wire gpio_out_gpio_out_2_qs;
	// Trace: design.sv:54022:3
	wire gpio_out_gpio_out_2_wd;
	// Trace: design.sv:54023:3
	wire gpio_out_gpio_out_2_we;
	// Trace: design.sv:54024:3
	wire gpio_out_gpio_out_3_qs;
	// Trace: design.sv:54025:3
	wire gpio_out_gpio_out_3_wd;
	// Trace: design.sv:54026:3
	wire gpio_out_gpio_out_3_we;
	// Trace: design.sv:54027:3
	wire gpio_out_gpio_out_4_qs;
	// Trace: design.sv:54028:3
	wire gpio_out_gpio_out_4_wd;
	// Trace: design.sv:54029:3
	wire gpio_out_gpio_out_4_we;
	// Trace: design.sv:54030:3
	wire gpio_out_gpio_out_5_qs;
	// Trace: design.sv:54031:3
	wire gpio_out_gpio_out_5_wd;
	// Trace: design.sv:54032:3
	wire gpio_out_gpio_out_5_we;
	// Trace: design.sv:54033:3
	wire gpio_out_gpio_out_6_qs;
	// Trace: design.sv:54034:3
	wire gpio_out_gpio_out_6_wd;
	// Trace: design.sv:54035:3
	wire gpio_out_gpio_out_6_we;
	// Trace: design.sv:54036:3
	wire gpio_out_gpio_out_7_qs;
	// Trace: design.sv:54037:3
	wire gpio_out_gpio_out_7_wd;
	// Trace: design.sv:54038:3
	wire gpio_out_gpio_out_7_we;
	// Trace: design.sv:54039:3
	wire gpio_out_gpio_out_8_qs;
	// Trace: design.sv:54040:3
	wire gpio_out_gpio_out_8_wd;
	// Trace: design.sv:54041:3
	wire gpio_out_gpio_out_8_we;
	// Trace: design.sv:54042:3
	wire gpio_out_gpio_out_9_qs;
	// Trace: design.sv:54043:3
	wire gpio_out_gpio_out_9_wd;
	// Trace: design.sv:54044:3
	wire gpio_out_gpio_out_9_we;
	// Trace: design.sv:54045:3
	wire gpio_out_gpio_out_10_qs;
	// Trace: design.sv:54046:3
	wire gpio_out_gpio_out_10_wd;
	// Trace: design.sv:54047:3
	wire gpio_out_gpio_out_10_we;
	// Trace: design.sv:54048:3
	wire gpio_out_gpio_out_11_qs;
	// Trace: design.sv:54049:3
	wire gpio_out_gpio_out_11_wd;
	// Trace: design.sv:54050:3
	wire gpio_out_gpio_out_11_we;
	// Trace: design.sv:54051:3
	wire gpio_out_gpio_out_12_qs;
	// Trace: design.sv:54052:3
	wire gpio_out_gpio_out_12_wd;
	// Trace: design.sv:54053:3
	wire gpio_out_gpio_out_12_we;
	// Trace: design.sv:54054:3
	wire gpio_out_gpio_out_13_qs;
	// Trace: design.sv:54055:3
	wire gpio_out_gpio_out_13_wd;
	// Trace: design.sv:54056:3
	wire gpio_out_gpio_out_13_we;
	// Trace: design.sv:54057:3
	wire gpio_out_gpio_out_14_qs;
	// Trace: design.sv:54058:3
	wire gpio_out_gpio_out_14_wd;
	// Trace: design.sv:54059:3
	wire gpio_out_gpio_out_14_we;
	// Trace: design.sv:54060:3
	wire gpio_out_gpio_out_15_qs;
	// Trace: design.sv:54061:3
	wire gpio_out_gpio_out_15_wd;
	// Trace: design.sv:54062:3
	wire gpio_out_gpio_out_15_we;
	// Trace: design.sv:54063:3
	wire gpio_out_gpio_out_16_qs;
	// Trace: design.sv:54064:3
	wire gpio_out_gpio_out_16_wd;
	// Trace: design.sv:54065:3
	wire gpio_out_gpio_out_16_we;
	// Trace: design.sv:54066:3
	wire gpio_out_gpio_out_17_qs;
	// Trace: design.sv:54067:3
	wire gpio_out_gpio_out_17_wd;
	// Trace: design.sv:54068:3
	wire gpio_out_gpio_out_17_we;
	// Trace: design.sv:54069:3
	wire gpio_out_gpio_out_18_qs;
	// Trace: design.sv:54070:3
	wire gpio_out_gpio_out_18_wd;
	// Trace: design.sv:54071:3
	wire gpio_out_gpio_out_18_we;
	// Trace: design.sv:54072:3
	wire gpio_out_gpio_out_19_qs;
	// Trace: design.sv:54073:3
	wire gpio_out_gpio_out_19_wd;
	// Trace: design.sv:54074:3
	wire gpio_out_gpio_out_19_we;
	// Trace: design.sv:54075:3
	wire gpio_out_gpio_out_20_qs;
	// Trace: design.sv:54076:3
	wire gpio_out_gpio_out_20_wd;
	// Trace: design.sv:54077:3
	wire gpio_out_gpio_out_20_we;
	// Trace: design.sv:54078:3
	wire gpio_out_gpio_out_21_qs;
	// Trace: design.sv:54079:3
	wire gpio_out_gpio_out_21_wd;
	// Trace: design.sv:54080:3
	wire gpio_out_gpio_out_21_we;
	// Trace: design.sv:54081:3
	wire gpio_out_gpio_out_22_qs;
	// Trace: design.sv:54082:3
	wire gpio_out_gpio_out_22_wd;
	// Trace: design.sv:54083:3
	wire gpio_out_gpio_out_22_we;
	// Trace: design.sv:54084:3
	wire gpio_out_gpio_out_23_qs;
	// Trace: design.sv:54085:3
	wire gpio_out_gpio_out_23_wd;
	// Trace: design.sv:54086:3
	wire gpio_out_gpio_out_23_we;
	// Trace: design.sv:54087:3
	wire gpio_out_gpio_out_24_qs;
	// Trace: design.sv:54088:3
	wire gpio_out_gpio_out_24_wd;
	// Trace: design.sv:54089:3
	wire gpio_out_gpio_out_24_we;
	// Trace: design.sv:54090:3
	wire gpio_out_gpio_out_25_qs;
	// Trace: design.sv:54091:3
	wire gpio_out_gpio_out_25_wd;
	// Trace: design.sv:54092:3
	wire gpio_out_gpio_out_25_we;
	// Trace: design.sv:54093:3
	wire gpio_out_gpio_out_26_qs;
	// Trace: design.sv:54094:3
	wire gpio_out_gpio_out_26_wd;
	// Trace: design.sv:54095:3
	wire gpio_out_gpio_out_26_we;
	// Trace: design.sv:54096:3
	wire gpio_out_gpio_out_27_qs;
	// Trace: design.sv:54097:3
	wire gpio_out_gpio_out_27_wd;
	// Trace: design.sv:54098:3
	wire gpio_out_gpio_out_27_we;
	// Trace: design.sv:54099:3
	wire gpio_out_gpio_out_28_qs;
	// Trace: design.sv:54100:3
	wire gpio_out_gpio_out_28_wd;
	// Trace: design.sv:54101:3
	wire gpio_out_gpio_out_28_we;
	// Trace: design.sv:54102:3
	wire gpio_out_gpio_out_29_qs;
	// Trace: design.sv:54103:3
	wire gpio_out_gpio_out_29_wd;
	// Trace: design.sv:54104:3
	wire gpio_out_gpio_out_29_we;
	// Trace: design.sv:54105:3
	wire gpio_out_gpio_out_30_qs;
	// Trace: design.sv:54106:3
	wire gpio_out_gpio_out_30_wd;
	// Trace: design.sv:54107:3
	wire gpio_out_gpio_out_30_we;
	// Trace: design.sv:54108:3
	wire gpio_out_gpio_out_31_qs;
	// Trace: design.sv:54109:3
	wire gpio_out_gpio_out_31_wd;
	// Trace: design.sv:54110:3
	wire gpio_out_gpio_out_31_we;
	// Trace: design.sv:54111:3
	wire gpio_set_gpio_set_0_wd;
	// Trace: design.sv:54112:3
	wire gpio_set_gpio_set_0_we;
	// Trace: design.sv:54113:3
	wire gpio_set_gpio_set_1_wd;
	// Trace: design.sv:54114:3
	wire gpio_set_gpio_set_1_we;
	// Trace: design.sv:54115:3
	wire gpio_set_gpio_set_2_wd;
	// Trace: design.sv:54116:3
	wire gpio_set_gpio_set_2_we;
	// Trace: design.sv:54117:3
	wire gpio_set_gpio_set_3_wd;
	// Trace: design.sv:54118:3
	wire gpio_set_gpio_set_3_we;
	// Trace: design.sv:54119:3
	wire gpio_set_gpio_set_4_wd;
	// Trace: design.sv:54120:3
	wire gpio_set_gpio_set_4_we;
	// Trace: design.sv:54121:3
	wire gpio_set_gpio_set_5_wd;
	// Trace: design.sv:54122:3
	wire gpio_set_gpio_set_5_we;
	// Trace: design.sv:54123:3
	wire gpio_set_gpio_set_6_wd;
	// Trace: design.sv:54124:3
	wire gpio_set_gpio_set_6_we;
	// Trace: design.sv:54125:3
	wire gpio_set_gpio_set_7_wd;
	// Trace: design.sv:54126:3
	wire gpio_set_gpio_set_7_we;
	// Trace: design.sv:54127:3
	wire gpio_set_gpio_set_8_wd;
	// Trace: design.sv:54128:3
	wire gpio_set_gpio_set_8_we;
	// Trace: design.sv:54129:3
	wire gpio_set_gpio_set_9_wd;
	// Trace: design.sv:54130:3
	wire gpio_set_gpio_set_9_we;
	// Trace: design.sv:54131:3
	wire gpio_set_gpio_set_10_wd;
	// Trace: design.sv:54132:3
	wire gpio_set_gpio_set_10_we;
	// Trace: design.sv:54133:3
	wire gpio_set_gpio_set_11_wd;
	// Trace: design.sv:54134:3
	wire gpio_set_gpio_set_11_we;
	// Trace: design.sv:54135:3
	wire gpio_set_gpio_set_12_wd;
	// Trace: design.sv:54136:3
	wire gpio_set_gpio_set_12_we;
	// Trace: design.sv:54137:3
	wire gpio_set_gpio_set_13_wd;
	// Trace: design.sv:54138:3
	wire gpio_set_gpio_set_13_we;
	// Trace: design.sv:54139:3
	wire gpio_set_gpio_set_14_wd;
	// Trace: design.sv:54140:3
	wire gpio_set_gpio_set_14_we;
	// Trace: design.sv:54141:3
	wire gpio_set_gpio_set_15_wd;
	// Trace: design.sv:54142:3
	wire gpio_set_gpio_set_15_we;
	// Trace: design.sv:54143:3
	wire gpio_set_gpio_set_16_wd;
	// Trace: design.sv:54144:3
	wire gpio_set_gpio_set_16_we;
	// Trace: design.sv:54145:3
	wire gpio_set_gpio_set_17_wd;
	// Trace: design.sv:54146:3
	wire gpio_set_gpio_set_17_we;
	// Trace: design.sv:54147:3
	wire gpio_set_gpio_set_18_wd;
	// Trace: design.sv:54148:3
	wire gpio_set_gpio_set_18_we;
	// Trace: design.sv:54149:3
	wire gpio_set_gpio_set_19_wd;
	// Trace: design.sv:54150:3
	wire gpio_set_gpio_set_19_we;
	// Trace: design.sv:54151:3
	wire gpio_set_gpio_set_20_wd;
	// Trace: design.sv:54152:3
	wire gpio_set_gpio_set_20_we;
	// Trace: design.sv:54153:3
	wire gpio_set_gpio_set_21_wd;
	// Trace: design.sv:54154:3
	wire gpio_set_gpio_set_21_we;
	// Trace: design.sv:54155:3
	wire gpio_set_gpio_set_22_wd;
	// Trace: design.sv:54156:3
	wire gpio_set_gpio_set_22_we;
	// Trace: design.sv:54157:3
	wire gpio_set_gpio_set_23_wd;
	// Trace: design.sv:54158:3
	wire gpio_set_gpio_set_23_we;
	// Trace: design.sv:54159:3
	wire gpio_set_gpio_set_24_wd;
	// Trace: design.sv:54160:3
	wire gpio_set_gpio_set_24_we;
	// Trace: design.sv:54161:3
	wire gpio_set_gpio_set_25_wd;
	// Trace: design.sv:54162:3
	wire gpio_set_gpio_set_25_we;
	// Trace: design.sv:54163:3
	wire gpio_set_gpio_set_26_wd;
	// Trace: design.sv:54164:3
	wire gpio_set_gpio_set_26_we;
	// Trace: design.sv:54165:3
	wire gpio_set_gpio_set_27_wd;
	// Trace: design.sv:54166:3
	wire gpio_set_gpio_set_27_we;
	// Trace: design.sv:54167:3
	wire gpio_set_gpio_set_28_wd;
	// Trace: design.sv:54168:3
	wire gpio_set_gpio_set_28_we;
	// Trace: design.sv:54169:3
	wire gpio_set_gpio_set_29_wd;
	// Trace: design.sv:54170:3
	wire gpio_set_gpio_set_29_we;
	// Trace: design.sv:54171:3
	wire gpio_set_gpio_set_30_wd;
	// Trace: design.sv:54172:3
	wire gpio_set_gpio_set_30_we;
	// Trace: design.sv:54173:3
	wire gpio_set_gpio_set_31_wd;
	// Trace: design.sv:54174:3
	wire gpio_set_gpio_set_31_we;
	// Trace: design.sv:54175:3
	wire gpio_clear_gpio_clear_0_wd;
	// Trace: design.sv:54176:3
	wire gpio_clear_gpio_clear_0_we;
	// Trace: design.sv:54177:3
	wire gpio_clear_gpio_clear_1_wd;
	// Trace: design.sv:54178:3
	wire gpio_clear_gpio_clear_1_we;
	// Trace: design.sv:54179:3
	wire gpio_clear_gpio_clear_2_wd;
	// Trace: design.sv:54180:3
	wire gpio_clear_gpio_clear_2_we;
	// Trace: design.sv:54181:3
	wire gpio_clear_gpio_clear_3_wd;
	// Trace: design.sv:54182:3
	wire gpio_clear_gpio_clear_3_we;
	// Trace: design.sv:54183:3
	wire gpio_clear_gpio_clear_4_wd;
	// Trace: design.sv:54184:3
	wire gpio_clear_gpio_clear_4_we;
	// Trace: design.sv:54185:3
	wire gpio_clear_gpio_clear_5_wd;
	// Trace: design.sv:54186:3
	wire gpio_clear_gpio_clear_5_we;
	// Trace: design.sv:54187:3
	wire gpio_clear_gpio_clear_6_wd;
	// Trace: design.sv:54188:3
	wire gpio_clear_gpio_clear_6_we;
	// Trace: design.sv:54189:3
	wire gpio_clear_gpio_clear_7_wd;
	// Trace: design.sv:54190:3
	wire gpio_clear_gpio_clear_7_we;
	// Trace: design.sv:54191:3
	wire gpio_clear_gpio_clear_8_wd;
	// Trace: design.sv:54192:3
	wire gpio_clear_gpio_clear_8_we;
	// Trace: design.sv:54193:3
	wire gpio_clear_gpio_clear_9_wd;
	// Trace: design.sv:54194:3
	wire gpio_clear_gpio_clear_9_we;
	// Trace: design.sv:54195:3
	wire gpio_clear_gpio_clear_10_wd;
	// Trace: design.sv:54196:3
	wire gpio_clear_gpio_clear_10_we;
	// Trace: design.sv:54197:3
	wire gpio_clear_gpio_clear_11_wd;
	// Trace: design.sv:54198:3
	wire gpio_clear_gpio_clear_11_we;
	// Trace: design.sv:54199:3
	wire gpio_clear_gpio_clear_12_wd;
	// Trace: design.sv:54200:3
	wire gpio_clear_gpio_clear_12_we;
	// Trace: design.sv:54201:3
	wire gpio_clear_gpio_clear_13_wd;
	// Trace: design.sv:54202:3
	wire gpio_clear_gpio_clear_13_we;
	// Trace: design.sv:54203:3
	wire gpio_clear_gpio_clear_14_wd;
	// Trace: design.sv:54204:3
	wire gpio_clear_gpio_clear_14_we;
	// Trace: design.sv:54205:3
	wire gpio_clear_gpio_clear_15_wd;
	// Trace: design.sv:54206:3
	wire gpio_clear_gpio_clear_15_we;
	// Trace: design.sv:54207:3
	wire gpio_clear_gpio_clear_16_wd;
	// Trace: design.sv:54208:3
	wire gpio_clear_gpio_clear_16_we;
	// Trace: design.sv:54209:3
	wire gpio_clear_gpio_clear_17_wd;
	// Trace: design.sv:54210:3
	wire gpio_clear_gpio_clear_17_we;
	// Trace: design.sv:54211:3
	wire gpio_clear_gpio_clear_18_wd;
	// Trace: design.sv:54212:3
	wire gpio_clear_gpio_clear_18_we;
	// Trace: design.sv:54213:3
	wire gpio_clear_gpio_clear_19_wd;
	// Trace: design.sv:54214:3
	wire gpio_clear_gpio_clear_19_we;
	// Trace: design.sv:54215:3
	wire gpio_clear_gpio_clear_20_wd;
	// Trace: design.sv:54216:3
	wire gpio_clear_gpio_clear_20_we;
	// Trace: design.sv:54217:3
	wire gpio_clear_gpio_clear_21_wd;
	// Trace: design.sv:54218:3
	wire gpio_clear_gpio_clear_21_we;
	// Trace: design.sv:54219:3
	wire gpio_clear_gpio_clear_22_wd;
	// Trace: design.sv:54220:3
	wire gpio_clear_gpio_clear_22_we;
	// Trace: design.sv:54221:3
	wire gpio_clear_gpio_clear_23_wd;
	// Trace: design.sv:54222:3
	wire gpio_clear_gpio_clear_23_we;
	// Trace: design.sv:54223:3
	wire gpio_clear_gpio_clear_24_wd;
	// Trace: design.sv:54224:3
	wire gpio_clear_gpio_clear_24_we;
	// Trace: design.sv:54225:3
	wire gpio_clear_gpio_clear_25_wd;
	// Trace: design.sv:54226:3
	wire gpio_clear_gpio_clear_25_we;
	// Trace: design.sv:54227:3
	wire gpio_clear_gpio_clear_26_wd;
	// Trace: design.sv:54228:3
	wire gpio_clear_gpio_clear_26_we;
	// Trace: design.sv:54229:3
	wire gpio_clear_gpio_clear_27_wd;
	// Trace: design.sv:54230:3
	wire gpio_clear_gpio_clear_27_we;
	// Trace: design.sv:54231:3
	wire gpio_clear_gpio_clear_28_wd;
	// Trace: design.sv:54232:3
	wire gpio_clear_gpio_clear_28_we;
	// Trace: design.sv:54233:3
	wire gpio_clear_gpio_clear_29_wd;
	// Trace: design.sv:54234:3
	wire gpio_clear_gpio_clear_29_we;
	// Trace: design.sv:54235:3
	wire gpio_clear_gpio_clear_30_wd;
	// Trace: design.sv:54236:3
	wire gpio_clear_gpio_clear_30_we;
	// Trace: design.sv:54237:3
	wire gpio_clear_gpio_clear_31_wd;
	// Trace: design.sv:54238:3
	wire gpio_clear_gpio_clear_31_we;
	// Trace: design.sv:54239:3
	wire gpio_toggle_gpio_toggle_0_wd;
	// Trace: design.sv:54240:3
	wire gpio_toggle_gpio_toggle_0_we;
	// Trace: design.sv:54241:3
	wire gpio_toggle_gpio_toggle_1_wd;
	// Trace: design.sv:54242:3
	wire gpio_toggle_gpio_toggle_1_we;
	// Trace: design.sv:54243:3
	wire gpio_toggle_gpio_toggle_2_wd;
	// Trace: design.sv:54244:3
	wire gpio_toggle_gpio_toggle_2_we;
	// Trace: design.sv:54245:3
	wire gpio_toggle_gpio_toggle_3_wd;
	// Trace: design.sv:54246:3
	wire gpio_toggle_gpio_toggle_3_we;
	// Trace: design.sv:54247:3
	wire gpio_toggle_gpio_toggle_4_wd;
	// Trace: design.sv:54248:3
	wire gpio_toggle_gpio_toggle_4_we;
	// Trace: design.sv:54249:3
	wire gpio_toggle_gpio_toggle_5_wd;
	// Trace: design.sv:54250:3
	wire gpio_toggle_gpio_toggle_5_we;
	// Trace: design.sv:54251:3
	wire gpio_toggle_gpio_toggle_6_wd;
	// Trace: design.sv:54252:3
	wire gpio_toggle_gpio_toggle_6_we;
	// Trace: design.sv:54253:3
	wire gpio_toggle_gpio_toggle_7_wd;
	// Trace: design.sv:54254:3
	wire gpio_toggle_gpio_toggle_7_we;
	// Trace: design.sv:54255:3
	wire gpio_toggle_gpio_toggle_8_wd;
	// Trace: design.sv:54256:3
	wire gpio_toggle_gpio_toggle_8_we;
	// Trace: design.sv:54257:3
	wire gpio_toggle_gpio_toggle_9_wd;
	// Trace: design.sv:54258:3
	wire gpio_toggle_gpio_toggle_9_we;
	// Trace: design.sv:54259:3
	wire gpio_toggle_gpio_toggle_10_wd;
	// Trace: design.sv:54260:3
	wire gpio_toggle_gpio_toggle_10_we;
	// Trace: design.sv:54261:3
	wire gpio_toggle_gpio_toggle_11_wd;
	// Trace: design.sv:54262:3
	wire gpio_toggle_gpio_toggle_11_we;
	// Trace: design.sv:54263:3
	wire gpio_toggle_gpio_toggle_12_wd;
	// Trace: design.sv:54264:3
	wire gpio_toggle_gpio_toggle_12_we;
	// Trace: design.sv:54265:3
	wire gpio_toggle_gpio_toggle_13_wd;
	// Trace: design.sv:54266:3
	wire gpio_toggle_gpio_toggle_13_we;
	// Trace: design.sv:54267:3
	wire gpio_toggle_gpio_toggle_14_wd;
	// Trace: design.sv:54268:3
	wire gpio_toggle_gpio_toggle_14_we;
	// Trace: design.sv:54269:3
	wire gpio_toggle_gpio_toggle_15_wd;
	// Trace: design.sv:54270:3
	wire gpio_toggle_gpio_toggle_15_we;
	// Trace: design.sv:54271:3
	wire gpio_toggle_gpio_toggle_16_wd;
	// Trace: design.sv:54272:3
	wire gpio_toggle_gpio_toggle_16_we;
	// Trace: design.sv:54273:3
	wire gpio_toggle_gpio_toggle_17_wd;
	// Trace: design.sv:54274:3
	wire gpio_toggle_gpio_toggle_17_we;
	// Trace: design.sv:54275:3
	wire gpio_toggle_gpio_toggle_18_wd;
	// Trace: design.sv:54276:3
	wire gpio_toggle_gpio_toggle_18_we;
	// Trace: design.sv:54277:3
	wire gpio_toggle_gpio_toggle_19_wd;
	// Trace: design.sv:54278:3
	wire gpio_toggle_gpio_toggle_19_we;
	// Trace: design.sv:54279:3
	wire gpio_toggle_gpio_toggle_20_wd;
	// Trace: design.sv:54280:3
	wire gpio_toggle_gpio_toggle_20_we;
	// Trace: design.sv:54281:3
	wire gpio_toggle_gpio_toggle_21_wd;
	// Trace: design.sv:54282:3
	wire gpio_toggle_gpio_toggle_21_we;
	// Trace: design.sv:54283:3
	wire gpio_toggle_gpio_toggle_22_wd;
	// Trace: design.sv:54284:3
	wire gpio_toggle_gpio_toggle_22_we;
	// Trace: design.sv:54285:3
	wire gpio_toggle_gpio_toggle_23_wd;
	// Trace: design.sv:54286:3
	wire gpio_toggle_gpio_toggle_23_we;
	// Trace: design.sv:54287:3
	wire gpio_toggle_gpio_toggle_24_wd;
	// Trace: design.sv:54288:3
	wire gpio_toggle_gpio_toggle_24_we;
	// Trace: design.sv:54289:3
	wire gpio_toggle_gpio_toggle_25_wd;
	// Trace: design.sv:54290:3
	wire gpio_toggle_gpio_toggle_25_we;
	// Trace: design.sv:54291:3
	wire gpio_toggle_gpio_toggle_26_wd;
	// Trace: design.sv:54292:3
	wire gpio_toggle_gpio_toggle_26_we;
	// Trace: design.sv:54293:3
	wire gpio_toggle_gpio_toggle_27_wd;
	// Trace: design.sv:54294:3
	wire gpio_toggle_gpio_toggle_27_we;
	// Trace: design.sv:54295:3
	wire gpio_toggle_gpio_toggle_28_wd;
	// Trace: design.sv:54296:3
	wire gpio_toggle_gpio_toggle_28_we;
	// Trace: design.sv:54297:3
	wire gpio_toggle_gpio_toggle_29_wd;
	// Trace: design.sv:54298:3
	wire gpio_toggle_gpio_toggle_29_we;
	// Trace: design.sv:54299:3
	wire gpio_toggle_gpio_toggle_30_wd;
	// Trace: design.sv:54300:3
	wire gpio_toggle_gpio_toggle_30_we;
	// Trace: design.sv:54301:3
	wire gpio_toggle_gpio_toggle_31_wd;
	// Trace: design.sv:54302:3
	wire gpio_toggle_gpio_toggle_31_we;
	// Trace: design.sv:54303:3
	wire intrpt_rise_en_intrpt_rise_en_0_qs;
	// Trace: design.sv:54304:3
	wire intrpt_rise_en_intrpt_rise_en_0_wd;
	// Trace: design.sv:54305:3
	wire intrpt_rise_en_intrpt_rise_en_0_we;
	// Trace: design.sv:54306:3
	wire intrpt_rise_en_intrpt_rise_en_1_qs;
	// Trace: design.sv:54307:3
	wire intrpt_rise_en_intrpt_rise_en_1_wd;
	// Trace: design.sv:54308:3
	wire intrpt_rise_en_intrpt_rise_en_1_we;
	// Trace: design.sv:54309:3
	wire intrpt_rise_en_intrpt_rise_en_2_qs;
	// Trace: design.sv:54310:3
	wire intrpt_rise_en_intrpt_rise_en_2_wd;
	// Trace: design.sv:54311:3
	wire intrpt_rise_en_intrpt_rise_en_2_we;
	// Trace: design.sv:54312:3
	wire intrpt_rise_en_intrpt_rise_en_3_qs;
	// Trace: design.sv:54313:3
	wire intrpt_rise_en_intrpt_rise_en_3_wd;
	// Trace: design.sv:54314:3
	wire intrpt_rise_en_intrpt_rise_en_3_we;
	// Trace: design.sv:54315:3
	wire intrpt_rise_en_intrpt_rise_en_4_qs;
	// Trace: design.sv:54316:3
	wire intrpt_rise_en_intrpt_rise_en_4_wd;
	// Trace: design.sv:54317:3
	wire intrpt_rise_en_intrpt_rise_en_4_we;
	// Trace: design.sv:54318:3
	wire intrpt_rise_en_intrpt_rise_en_5_qs;
	// Trace: design.sv:54319:3
	wire intrpt_rise_en_intrpt_rise_en_5_wd;
	// Trace: design.sv:54320:3
	wire intrpt_rise_en_intrpt_rise_en_5_we;
	// Trace: design.sv:54321:3
	wire intrpt_rise_en_intrpt_rise_en_6_qs;
	// Trace: design.sv:54322:3
	wire intrpt_rise_en_intrpt_rise_en_6_wd;
	// Trace: design.sv:54323:3
	wire intrpt_rise_en_intrpt_rise_en_6_we;
	// Trace: design.sv:54324:3
	wire intrpt_rise_en_intrpt_rise_en_7_qs;
	// Trace: design.sv:54325:3
	wire intrpt_rise_en_intrpt_rise_en_7_wd;
	// Trace: design.sv:54326:3
	wire intrpt_rise_en_intrpt_rise_en_7_we;
	// Trace: design.sv:54327:3
	wire intrpt_rise_en_intrpt_rise_en_8_qs;
	// Trace: design.sv:54328:3
	wire intrpt_rise_en_intrpt_rise_en_8_wd;
	// Trace: design.sv:54329:3
	wire intrpt_rise_en_intrpt_rise_en_8_we;
	// Trace: design.sv:54330:3
	wire intrpt_rise_en_intrpt_rise_en_9_qs;
	// Trace: design.sv:54331:3
	wire intrpt_rise_en_intrpt_rise_en_9_wd;
	// Trace: design.sv:54332:3
	wire intrpt_rise_en_intrpt_rise_en_9_we;
	// Trace: design.sv:54333:3
	wire intrpt_rise_en_intrpt_rise_en_10_qs;
	// Trace: design.sv:54334:3
	wire intrpt_rise_en_intrpt_rise_en_10_wd;
	// Trace: design.sv:54335:3
	wire intrpt_rise_en_intrpt_rise_en_10_we;
	// Trace: design.sv:54336:3
	wire intrpt_rise_en_intrpt_rise_en_11_qs;
	// Trace: design.sv:54337:3
	wire intrpt_rise_en_intrpt_rise_en_11_wd;
	// Trace: design.sv:54338:3
	wire intrpt_rise_en_intrpt_rise_en_11_we;
	// Trace: design.sv:54339:3
	wire intrpt_rise_en_intrpt_rise_en_12_qs;
	// Trace: design.sv:54340:3
	wire intrpt_rise_en_intrpt_rise_en_12_wd;
	// Trace: design.sv:54341:3
	wire intrpt_rise_en_intrpt_rise_en_12_we;
	// Trace: design.sv:54342:3
	wire intrpt_rise_en_intrpt_rise_en_13_qs;
	// Trace: design.sv:54343:3
	wire intrpt_rise_en_intrpt_rise_en_13_wd;
	// Trace: design.sv:54344:3
	wire intrpt_rise_en_intrpt_rise_en_13_we;
	// Trace: design.sv:54345:3
	wire intrpt_rise_en_intrpt_rise_en_14_qs;
	// Trace: design.sv:54346:3
	wire intrpt_rise_en_intrpt_rise_en_14_wd;
	// Trace: design.sv:54347:3
	wire intrpt_rise_en_intrpt_rise_en_14_we;
	// Trace: design.sv:54348:3
	wire intrpt_rise_en_intrpt_rise_en_15_qs;
	// Trace: design.sv:54349:3
	wire intrpt_rise_en_intrpt_rise_en_15_wd;
	// Trace: design.sv:54350:3
	wire intrpt_rise_en_intrpt_rise_en_15_we;
	// Trace: design.sv:54351:3
	wire intrpt_rise_en_intrpt_rise_en_16_qs;
	// Trace: design.sv:54352:3
	wire intrpt_rise_en_intrpt_rise_en_16_wd;
	// Trace: design.sv:54353:3
	wire intrpt_rise_en_intrpt_rise_en_16_we;
	// Trace: design.sv:54354:3
	wire intrpt_rise_en_intrpt_rise_en_17_qs;
	// Trace: design.sv:54355:3
	wire intrpt_rise_en_intrpt_rise_en_17_wd;
	// Trace: design.sv:54356:3
	wire intrpt_rise_en_intrpt_rise_en_17_we;
	// Trace: design.sv:54357:3
	wire intrpt_rise_en_intrpt_rise_en_18_qs;
	// Trace: design.sv:54358:3
	wire intrpt_rise_en_intrpt_rise_en_18_wd;
	// Trace: design.sv:54359:3
	wire intrpt_rise_en_intrpt_rise_en_18_we;
	// Trace: design.sv:54360:3
	wire intrpt_rise_en_intrpt_rise_en_19_qs;
	// Trace: design.sv:54361:3
	wire intrpt_rise_en_intrpt_rise_en_19_wd;
	// Trace: design.sv:54362:3
	wire intrpt_rise_en_intrpt_rise_en_19_we;
	// Trace: design.sv:54363:3
	wire intrpt_rise_en_intrpt_rise_en_20_qs;
	// Trace: design.sv:54364:3
	wire intrpt_rise_en_intrpt_rise_en_20_wd;
	// Trace: design.sv:54365:3
	wire intrpt_rise_en_intrpt_rise_en_20_we;
	// Trace: design.sv:54366:3
	wire intrpt_rise_en_intrpt_rise_en_21_qs;
	// Trace: design.sv:54367:3
	wire intrpt_rise_en_intrpt_rise_en_21_wd;
	// Trace: design.sv:54368:3
	wire intrpt_rise_en_intrpt_rise_en_21_we;
	// Trace: design.sv:54369:3
	wire intrpt_rise_en_intrpt_rise_en_22_qs;
	// Trace: design.sv:54370:3
	wire intrpt_rise_en_intrpt_rise_en_22_wd;
	// Trace: design.sv:54371:3
	wire intrpt_rise_en_intrpt_rise_en_22_we;
	// Trace: design.sv:54372:3
	wire intrpt_rise_en_intrpt_rise_en_23_qs;
	// Trace: design.sv:54373:3
	wire intrpt_rise_en_intrpt_rise_en_23_wd;
	// Trace: design.sv:54374:3
	wire intrpt_rise_en_intrpt_rise_en_23_we;
	// Trace: design.sv:54375:3
	wire intrpt_rise_en_intrpt_rise_en_24_qs;
	// Trace: design.sv:54376:3
	wire intrpt_rise_en_intrpt_rise_en_24_wd;
	// Trace: design.sv:54377:3
	wire intrpt_rise_en_intrpt_rise_en_24_we;
	// Trace: design.sv:54378:3
	wire intrpt_rise_en_intrpt_rise_en_25_qs;
	// Trace: design.sv:54379:3
	wire intrpt_rise_en_intrpt_rise_en_25_wd;
	// Trace: design.sv:54380:3
	wire intrpt_rise_en_intrpt_rise_en_25_we;
	// Trace: design.sv:54381:3
	wire intrpt_rise_en_intrpt_rise_en_26_qs;
	// Trace: design.sv:54382:3
	wire intrpt_rise_en_intrpt_rise_en_26_wd;
	// Trace: design.sv:54383:3
	wire intrpt_rise_en_intrpt_rise_en_26_we;
	// Trace: design.sv:54384:3
	wire intrpt_rise_en_intrpt_rise_en_27_qs;
	// Trace: design.sv:54385:3
	wire intrpt_rise_en_intrpt_rise_en_27_wd;
	// Trace: design.sv:54386:3
	wire intrpt_rise_en_intrpt_rise_en_27_we;
	// Trace: design.sv:54387:3
	wire intrpt_rise_en_intrpt_rise_en_28_qs;
	// Trace: design.sv:54388:3
	wire intrpt_rise_en_intrpt_rise_en_28_wd;
	// Trace: design.sv:54389:3
	wire intrpt_rise_en_intrpt_rise_en_28_we;
	// Trace: design.sv:54390:3
	wire intrpt_rise_en_intrpt_rise_en_29_qs;
	// Trace: design.sv:54391:3
	wire intrpt_rise_en_intrpt_rise_en_29_wd;
	// Trace: design.sv:54392:3
	wire intrpt_rise_en_intrpt_rise_en_29_we;
	// Trace: design.sv:54393:3
	wire intrpt_rise_en_intrpt_rise_en_30_qs;
	// Trace: design.sv:54394:3
	wire intrpt_rise_en_intrpt_rise_en_30_wd;
	// Trace: design.sv:54395:3
	wire intrpt_rise_en_intrpt_rise_en_30_we;
	// Trace: design.sv:54396:3
	wire intrpt_rise_en_intrpt_rise_en_31_qs;
	// Trace: design.sv:54397:3
	wire intrpt_rise_en_intrpt_rise_en_31_wd;
	// Trace: design.sv:54398:3
	wire intrpt_rise_en_intrpt_rise_en_31_we;
	// Trace: design.sv:54399:3
	wire intrpt_fall_en_intrpt_fall_en_0_qs;
	// Trace: design.sv:54400:3
	wire intrpt_fall_en_intrpt_fall_en_0_wd;
	// Trace: design.sv:54401:3
	wire intrpt_fall_en_intrpt_fall_en_0_we;
	// Trace: design.sv:54402:3
	wire intrpt_fall_en_intrpt_fall_en_1_qs;
	// Trace: design.sv:54403:3
	wire intrpt_fall_en_intrpt_fall_en_1_wd;
	// Trace: design.sv:54404:3
	wire intrpt_fall_en_intrpt_fall_en_1_we;
	// Trace: design.sv:54405:3
	wire intrpt_fall_en_intrpt_fall_en_2_qs;
	// Trace: design.sv:54406:3
	wire intrpt_fall_en_intrpt_fall_en_2_wd;
	// Trace: design.sv:54407:3
	wire intrpt_fall_en_intrpt_fall_en_2_we;
	// Trace: design.sv:54408:3
	wire intrpt_fall_en_intrpt_fall_en_3_qs;
	// Trace: design.sv:54409:3
	wire intrpt_fall_en_intrpt_fall_en_3_wd;
	// Trace: design.sv:54410:3
	wire intrpt_fall_en_intrpt_fall_en_3_we;
	// Trace: design.sv:54411:3
	wire intrpt_fall_en_intrpt_fall_en_4_qs;
	// Trace: design.sv:54412:3
	wire intrpt_fall_en_intrpt_fall_en_4_wd;
	// Trace: design.sv:54413:3
	wire intrpt_fall_en_intrpt_fall_en_4_we;
	// Trace: design.sv:54414:3
	wire intrpt_fall_en_intrpt_fall_en_5_qs;
	// Trace: design.sv:54415:3
	wire intrpt_fall_en_intrpt_fall_en_5_wd;
	// Trace: design.sv:54416:3
	wire intrpt_fall_en_intrpt_fall_en_5_we;
	// Trace: design.sv:54417:3
	wire intrpt_fall_en_intrpt_fall_en_6_qs;
	// Trace: design.sv:54418:3
	wire intrpt_fall_en_intrpt_fall_en_6_wd;
	// Trace: design.sv:54419:3
	wire intrpt_fall_en_intrpt_fall_en_6_we;
	// Trace: design.sv:54420:3
	wire intrpt_fall_en_intrpt_fall_en_7_qs;
	// Trace: design.sv:54421:3
	wire intrpt_fall_en_intrpt_fall_en_7_wd;
	// Trace: design.sv:54422:3
	wire intrpt_fall_en_intrpt_fall_en_7_we;
	// Trace: design.sv:54423:3
	wire intrpt_fall_en_intrpt_fall_en_8_qs;
	// Trace: design.sv:54424:3
	wire intrpt_fall_en_intrpt_fall_en_8_wd;
	// Trace: design.sv:54425:3
	wire intrpt_fall_en_intrpt_fall_en_8_we;
	// Trace: design.sv:54426:3
	wire intrpt_fall_en_intrpt_fall_en_9_qs;
	// Trace: design.sv:54427:3
	wire intrpt_fall_en_intrpt_fall_en_9_wd;
	// Trace: design.sv:54428:3
	wire intrpt_fall_en_intrpt_fall_en_9_we;
	// Trace: design.sv:54429:3
	wire intrpt_fall_en_intrpt_fall_en_10_qs;
	// Trace: design.sv:54430:3
	wire intrpt_fall_en_intrpt_fall_en_10_wd;
	// Trace: design.sv:54431:3
	wire intrpt_fall_en_intrpt_fall_en_10_we;
	// Trace: design.sv:54432:3
	wire intrpt_fall_en_intrpt_fall_en_11_qs;
	// Trace: design.sv:54433:3
	wire intrpt_fall_en_intrpt_fall_en_11_wd;
	// Trace: design.sv:54434:3
	wire intrpt_fall_en_intrpt_fall_en_11_we;
	// Trace: design.sv:54435:3
	wire intrpt_fall_en_intrpt_fall_en_12_qs;
	// Trace: design.sv:54436:3
	wire intrpt_fall_en_intrpt_fall_en_12_wd;
	// Trace: design.sv:54437:3
	wire intrpt_fall_en_intrpt_fall_en_12_we;
	// Trace: design.sv:54438:3
	wire intrpt_fall_en_intrpt_fall_en_13_qs;
	// Trace: design.sv:54439:3
	wire intrpt_fall_en_intrpt_fall_en_13_wd;
	// Trace: design.sv:54440:3
	wire intrpt_fall_en_intrpt_fall_en_13_we;
	// Trace: design.sv:54441:3
	wire intrpt_fall_en_intrpt_fall_en_14_qs;
	// Trace: design.sv:54442:3
	wire intrpt_fall_en_intrpt_fall_en_14_wd;
	// Trace: design.sv:54443:3
	wire intrpt_fall_en_intrpt_fall_en_14_we;
	// Trace: design.sv:54444:3
	wire intrpt_fall_en_intrpt_fall_en_15_qs;
	// Trace: design.sv:54445:3
	wire intrpt_fall_en_intrpt_fall_en_15_wd;
	// Trace: design.sv:54446:3
	wire intrpt_fall_en_intrpt_fall_en_15_we;
	// Trace: design.sv:54447:3
	wire intrpt_fall_en_intrpt_fall_en_16_qs;
	// Trace: design.sv:54448:3
	wire intrpt_fall_en_intrpt_fall_en_16_wd;
	// Trace: design.sv:54449:3
	wire intrpt_fall_en_intrpt_fall_en_16_we;
	// Trace: design.sv:54450:3
	wire intrpt_fall_en_intrpt_fall_en_17_qs;
	// Trace: design.sv:54451:3
	wire intrpt_fall_en_intrpt_fall_en_17_wd;
	// Trace: design.sv:54452:3
	wire intrpt_fall_en_intrpt_fall_en_17_we;
	// Trace: design.sv:54453:3
	wire intrpt_fall_en_intrpt_fall_en_18_qs;
	// Trace: design.sv:54454:3
	wire intrpt_fall_en_intrpt_fall_en_18_wd;
	// Trace: design.sv:54455:3
	wire intrpt_fall_en_intrpt_fall_en_18_we;
	// Trace: design.sv:54456:3
	wire intrpt_fall_en_intrpt_fall_en_19_qs;
	// Trace: design.sv:54457:3
	wire intrpt_fall_en_intrpt_fall_en_19_wd;
	// Trace: design.sv:54458:3
	wire intrpt_fall_en_intrpt_fall_en_19_we;
	// Trace: design.sv:54459:3
	wire intrpt_fall_en_intrpt_fall_en_20_qs;
	// Trace: design.sv:54460:3
	wire intrpt_fall_en_intrpt_fall_en_20_wd;
	// Trace: design.sv:54461:3
	wire intrpt_fall_en_intrpt_fall_en_20_we;
	// Trace: design.sv:54462:3
	wire intrpt_fall_en_intrpt_fall_en_21_qs;
	// Trace: design.sv:54463:3
	wire intrpt_fall_en_intrpt_fall_en_21_wd;
	// Trace: design.sv:54464:3
	wire intrpt_fall_en_intrpt_fall_en_21_we;
	// Trace: design.sv:54465:3
	wire intrpt_fall_en_intrpt_fall_en_22_qs;
	// Trace: design.sv:54466:3
	wire intrpt_fall_en_intrpt_fall_en_22_wd;
	// Trace: design.sv:54467:3
	wire intrpt_fall_en_intrpt_fall_en_22_we;
	// Trace: design.sv:54468:3
	wire intrpt_fall_en_intrpt_fall_en_23_qs;
	// Trace: design.sv:54469:3
	wire intrpt_fall_en_intrpt_fall_en_23_wd;
	// Trace: design.sv:54470:3
	wire intrpt_fall_en_intrpt_fall_en_23_we;
	// Trace: design.sv:54471:3
	wire intrpt_fall_en_intrpt_fall_en_24_qs;
	// Trace: design.sv:54472:3
	wire intrpt_fall_en_intrpt_fall_en_24_wd;
	// Trace: design.sv:54473:3
	wire intrpt_fall_en_intrpt_fall_en_24_we;
	// Trace: design.sv:54474:3
	wire intrpt_fall_en_intrpt_fall_en_25_qs;
	// Trace: design.sv:54475:3
	wire intrpt_fall_en_intrpt_fall_en_25_wd;
	// Trace: design.sv:54476:3
	wire intrpt_fall_en_intrpt_fall_en_25_we;
	// Trace: design.sv:54477:3
	wire intrpt_fall_en_intrpt_fall_en_26_qs;
	// Trace: design.sv:54478:3
	wire intrpt_fall_en_intrpt_fall_en_26_wd;
	// Trace: design.sv:54479:3
	wire intrpt_fall_en_intrpt_fall_en_26_we;
	// Trace: design.sv:54480:3
	wire intrpt_fall_en_intrpt_fall_en_27_qs;
	// Trace: design.sv:54481:3
	wire intrpt_fall_en_intrpt_fall_en_27_wd;
	// Trace: design.sv:54482:3
	wire intrpt_fall_en_intrpt_fall_en_27_we;
	// Trace: design.sv:54483:3
	wire intrpt_fall_en_intrpt_fall_en_28_qs;
	// Trace: design.sv:54484:3
	wire intrpt_fall_en_intrpt_fall_en_28_wd;
	// Trace: design.sv:54485:3
	wire intrpt_fall_en_intrpt_fall_en_28_we;
	// Trace: design.sv:54486:3
	wire intrpt_fall_en_intrpt_fall_en_29_qs;
	// Trace: design.sv:54487:3
	wire intrpt_fall_en_intrpt_fall_en_29_wd;
	// Trace: design.sv:54488:3
	wire intrpt_fall_en_intrpt_fall_en_29_we;
	// Trace: design.sv:54489:3
	wire intrpt_fall_en_intrpt_fall_en_30_qs;
	// Trace: design.sv:54490:3
	wire intrpt_fall_en_intrpt_fall_en_30_wd;
	// Trace: design.sv:54491:3
	wire intrpt_fall_en_intrpt_fall_en_30_we;
	// Trace: design.sv:54492:3
	wire intrpt_fall_en_intrpt_fall_en_31_qs;
	// Trace: design.sv:54493:3
	wire intrpt_fall_en_intrpt_fall_en_31_wd;
	// Trace: design.sv:54494:3
	wire intrpt_fall_en_intrpt_fall_en_31_we;
	// Trace: design.sv:54495:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_0_qs;
	// Trace: design.sv:54496:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_0_wd;
	// Trace: design.sv:54497:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_0_we;
	// Trace: design.sv:54498:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_1_qs;
	// Trace: design.sv:54499:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_1_wd;
	// Trace: design.sv:54500:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_1_we;
	// Trace: design.sv:54501:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_2_qs;
	// Trace: design.sv:54502:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_2_wd;
	// Trace: design.sv:54503:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_2_we;
	// Trace: design.sv:54504:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_3_qs;
	// Trace: design.sv:54505:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_3_wd;
	// Trace: design.sv:54506:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_3_we;
	// Trace: design.sv:54507:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_4_qs;
	// Trace: design.sv:54508:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_4_wd;
	// Trace: design.sv:54509:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_4_we;
	// Trace: design.sv:54510:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_5_qs;
	// Trace: design.sv:54511:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_5_wd;
	// Trace: design.sv:54512:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_5_we;
	// Trace: design.sv:54513:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_6_qs;
	// Trace: design.sv:54514:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_6_wd;
	// Trace: design.sv:54515:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_6_we;
	// Trace: design.sv:54516:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_7_qs;
	// Trace: design.sv:54517:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_7_wd;
	// Trace: design.sv:54518:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_7_we;
	// Trace: design.sv:54519:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_8_qs;
	// Trace: design.sv:54520:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_8_wd;
	// Trace: design.sv:54521:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_8_we;
	// Trace: design.sv:54522:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_9_qs;
	// Trace: design.sv:54523:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_9_wd;
	// Trace: design.sv:54524:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_9_we;
	// Trace: design.sv:54525:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_10_qs;
	// Trace: design.sv:54526:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_10_wd;
	// Trace: design.sv:54527:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_10_we;
	// Trace: design.sv:54528:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_11_qs;
	// Trace: design.sv:54529:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_11_wd;
	// Trace: design.sv:54530:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_11_we;
	// Trace: design.sv:54531:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_12_qs;
	// Trace: design.sv:54532:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_12_wd;
	// Trace: design.sv:54533:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_12_we;
	// Trace: design.sv:54534:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_13_qs;
	// Trace: design.sv:54535:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_13_wd;
	// Trace: design.sv:54536:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_13_we;
	// Trace: design.sv:54537:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_14_qs;
	// Trace: design.sv:54538:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_14_wd;
	// Trace: design.sv:54539:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_14_we;
	// Trace: design.sv:54540:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_15_qs;
	// Trace: design.sv:54541:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_15_wd;
	// Trace: design.sv:54542:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_15_we;
	// Trace: design.sv:54543:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_16_qs;
	// Trace: design.sv:54544:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_16_wd;
	// Trace: design.sv:54545:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_16_we;
	// Trace: design.sv:54546:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_17_qs;
	// Trace: design.sv:54547:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_17_wd;
	// Trace: design.sv:54548:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_17_we;
	// Trace: design.sv:54549:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_18_qs;
	// Trace: design.sv:54550:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_18_wd;
	// Trace: design.sv:54551:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_18_we;
	// Trace: design.sv:54552:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_19_qs;
	// Trace: design.sv:54553:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_19_wd;
	// Trace: design.sv:54554:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_19_we;
	// Trace: design.sv:54555:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_20_qs;
	// Trace: design.sv:54556:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_20_wd;
	// Trace: design.sv:54557:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_20_we;
	// Trace: design.sv:54558:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_21_qs;
	// Trace: design.sv:54559:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_21_wd;
	// Trace: design.sv:54560:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_21_we;
	// Trace: design.sv:54561:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_22_qs;
	// Trace: design.sv:54562:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_22_wd;
	// Trace: design.sv:54563:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_22_we;
	// Trace: design.sv:54564:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_23_qs;
	// Trace: design.sv:54565:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_23_wd;
	// Trace: design.sv:54566:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_23_we;
	// Trace: design.sv:54567:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_24_qs;
	// Trace: design.sv:54568:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_24_wd;
	// Trace: design.sv:54569:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_24_we;
	// Trace: design.sv:54570:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_25_qs;
	// Trace: design.sv:54571:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_25_wd;
	// Trace: design.sv:54572:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_25_we;
	// Trace: design.sv:54573:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_26_qs;
	// Trace: design.sv:54574:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_26_wd;
	// Trace: design.sv:54575:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_26_we;
	// Trace: design.sv:54576:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_27_qs;
	// Trace: design.sv:54577:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_27_wd;
	// Trace: design.sv:54578:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_27_we;
	// Trace: design.sv:54579:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_28_qs;
	// Trace: design.sv:54580:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_28_wd;
	// Trace: design.sv:54581:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_28_we;
	// Trace: design.sv:54582:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_29_qs;
	// Trace: design.sv:54583:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_29_wd;
	// Trace: design.sv:54584:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_29_we;
	// Trace: design.sv:54585:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_30_qs;
	// Trace: design.sv:54586:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_30_wd;
	// Trace: design.sv:54587:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_30_we;
	// Trace: design.sv:54588:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_31_qs;
	// Trace: design.sv:54589:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_31_wd;
	// Trace: design.sv:54590:3
	wire intrpt_lvl_high_en_intrpt_lvl_high_en_31_we;
	// Trace: design.sv:54591:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_0_qs;
	// Trace: design.sv:54592:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_0_wd;
	// Trace: design.sv:54593:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_0_we;
	// Trace: design.sv:54594:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_1_qs;
	// Trace: design.sv:54595:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_1_wd;
	// Trace: design.sv:54596:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_1_we;
	// Trace: design.sv:54597:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_2_qs;
	// Trace: design.sv:54598:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_2_wd;
	// Trace: design.sv:54599:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_2_we;
	// Trace: design.sv:54600:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_3_qs;
	// Trace: design.sv:54601:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_3_wd;
	// Trace: design.sv:54602:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_3_we;
	// Trace: design.sv:54603:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_4_qs;
	// Trace: design.sv:54604:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_4_wd;
	// Trace: design.sv:54605:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_4_we;
	// Trace: design.sv:54606:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_5_qs;
	// Trace: design.sv:54607:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_5_wd;
	// Trace: design.sv:54608:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_5_we;
	// Trace: design.sv:54609:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_6_qs;
	// Trace: design.sv:54610:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_6_wd;
	// Trace: design.sv:54611:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_6_we;
	// Trace: design.sv:54612:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_7_qs;
	// Trace: design.sv:54613:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_7_wd;
	// Trace: design.sv:54614:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_7_we;
	// Trace: design.sv:54615:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_8_qs;
	// Trace: design.sv:54616:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_8_wd;
	// Trace: design.sv:54617:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_8_we;
	// Trace: design.sv:54618:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_9_qs;
	// Trace: design.sv:54619:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_9_wd;
	// Trace: design.sv:54620:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_9_we;
	// Trace: design.sv:54621:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_10_qs;
	// Trace: design.sv:54622:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_10_wd;
	// Trace: design.sv:54623:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_10_we;
	// Trace: design.sv:54624:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_11_qs;
	// Trace: design.sv:54625:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_11_wd;
	// Trace: design.sv:54626:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_11_we;
	// Trace: design.sv:54627:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_12_qs;
	// Trace: design.sv:54628:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_12_wd;
	// Trace: design.sv:54629:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_12_we;
	// Trace: design.sv:54630:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_13_qs;
	// Trace: design.sv:54631:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_13_wd;
	// Trace: design.sv:54632:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_13_we;
	// Trace: design.sv:54633:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_14_qs;
	// Trace: design.sv:54634:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_14_wd;
	// Trace: design.sv:54635:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_14_we;
	// Trace: design.sv:54636:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_15_qs;
	// Trace: design.sv:54637:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_15_wd;
	// Trace: design.sv:54638:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_15_we;
	// Trace: design.sv:54639:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_16_qs;
	// Trace: design.sv:54640:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_16_wd;
	// Trace: design.sv:54641:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_16_we;
	// Trace: design.sv:54642:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_17_qs;
	// Trace: design.sv:54643:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_17_wd;
	// Trace: design.sv:54644:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_17_we;
	// Trace: design.sv:54645:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_18_qs;
	// Trace: design.sv:54646:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_18_wd;
	// Trace: design.sv:54647:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_18_we;
	// Trace: design.sv:54648:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_19_qs;
	// Trace: design.sv:54649:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_19_wd;
	// Trace: design.sv:54650:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_19_we;
	// Trace: design.sv:54651:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_20_qs;
	// Trace: design.sv:54652:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_20_wd;
	// Trace: design.sv:54653:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_20_we;
	// Trace: design.sv:54654:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_21_qs;
	// Trace: design.sv:54655:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_21_wd;
	// Trace: design.sv:54656:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_21_we;
	// Trace: design.sv:54657:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_22_qs;
	// Trace: design.sv:54658:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_22_wd;
	// Trace: design.sv:54659:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_22_we;
	// Trace: design.sv:54660:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_23_qs;
	// Trace: design.sv:54661:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_23_wd;
	// Trace: design.sv:54662:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_23_we;
	// Trace: design.sv:54663:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_24_qs;
	// Trace: design.sv:54664:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_24_wd;
	// Trace: design.sv:54665:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_24_we;
	// Trace: design.sv:54666:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_25_qs;
	// Trace: design.sv:54667:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_25_wd;
	// Trace: design.sv:54668:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_25_we;
	// Trace: design.sv:54669:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_26_qs;
	// Trace: design.sv:54670:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_26_wd;
	// Trace: design.sv:54671:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_26_we;
	// Trace: design.sv:54672:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_27_qs;
	// Trace: design.sv:54673:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_27_wd;
	// Trace: design.sv:54674:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_27_we;
	// Trace: design.sv:54675:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_28_qs;
	// Trace: design.sv:54676:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_28_wd;
	// Trace: design.sv:54677:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_28_we;
	// Trace: design.sv:54678:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_29_qs;
	// Trace: design.sv:54679:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_29_wd;
	// Trace: design.sv:54680:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_29_we;
	// Trace: design.sv:54681:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_30_qs;
	// Trace: design.sv:54682:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_30_wd;
	// Trace: design.sv:54683:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_30_we;
	// Trace: design.sv:54684:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_31_qs;
	// Trace: design.sv:54685:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_31_wd;
	// Trace: design.sv:54686:3
	wire intrpt_lvl_low_en_intrpt_lvl_low_en_31_we;
	// Trace: design.sv:54687:3
	wire intrpt_status_intrpt_status_0_qs;
	// Trace: design.sv:54688:3
	wire intrpt_status_intrpt_status_0_wd;
	// Trace: design.sv:54689:3
	wire intrpt_status_intrpt_status_0_we;
	// Trace: design.sv:54690:3
	wire intrpt_status_intrpt_status_0_re;
	// Trace: design.sv:54691:3
	wire intrpt_status_intrpt_status_1_qs;
	// Trace: design.sv:54692:3
	wire intrpt_status_intrpt_status_1_wd;
	// Trace: design.sv:54693:3
	wire intrpt_status_intrpt_status_1_we;
	// Trace: design.sv:54694:3
	wire intrpt_status_intrpt_status_1_re;
	// Trace: design.sv:54695:3
	wire intrpt_status_intrpt_status_2_qs;
	// Trace: design.sv:54696:3
	wire intrpt_status_intrpt_status_2_wd;
	// Trace: design.sv:54697:3
	wire intrpt_status_intrpt_status_2_we;
	// Trace: design.sv:54698:3
	wire intrpt_status_intrpt_status_2_re;
	// Trace: design.sv:54699:3
	wire intrpt_status_intrpt_status_3_qs;
	// Trace: design.sv:54700:3
	wire intrpt_status_intrpt_status_3_wd;
	// Trace: design.sv:54701:3
	wire intrpt_status_intrpt_status_3_we;
	// Trace: design.sv:54702:3
	wire intrpt_status_intrpt_status_3_re;
	// Trace: design.sv:54703:3
	wire intrpt_status_intrpt_status_4_qs;
	// Trace: design.sv:54704:3
	wire intrpt_status_intrpt_status_4_wd;
	// Trace: design.sv:54705:3
	wire intrpt_status_intrpt_status_4_we;
	// Trace: design.sv:54706:3
	wire intrpt_status_intrpt_status_4_re;
	// Trace: design.sv:54707:3
	wire intrpt_status_intrpt_status_5_qs;
	// Trace: design.sv:54708:3
	wire intrpt_status_intrpt_status_5_wd;
	// Trace: design.sv:54709:3
	wire intrpt_status_intrpt_status_5_we;
	// Trace: design.sv:54710:3
	wire intrpt_status_intrpt_status_5_re;
	// Trace: design.sv:54711:3
	wire intrpt_status_intrpt_status_6_qs;
	// Trace: design.sv:54712:3
	wire intrpt_status_intrpt_status_6_wd;
	// Trace: design.sv:54713:3
	wire intrpt_status_intrpt_status_6_we;
	// Trace: design.sv:54714:3
	wire intrpt_status_intrpt_status_6_re;
	// Trace: design.sv:54715:3
	wire intrpt_status_intrpt_status_7_qs;
	// Trace: design.sv:54716:3
	wire intrpt_status_intrpt_status_7_wd;
	// Trace: design.sv:54717:3
	wire intrpt_status_intrpt_status_7_we;
	// Trace: design.sv:54718:3
	wire intrpt_status_intrpt_status_7_re;
	// Trace: design.sv:54719:3
	wire intrpt_status_intrpt_status_8_qs;
	// Trace: design.sv:54720:3
	wire intrpt_status_intrpt_status_8_wd;
	// Trace: design.sv:54721:3
	wire intrpt_status_intrpt_status_8_we;
	// Trace: design.sv:54722:3
	wire intrpt_status_intrpt_status_8_re;
	// Trace: design.sv:54723:3
	wire intrpt_status_intrpt_status_9_qs;
	// Trace: design.sv:54724:3
	wire intrpt_status_intrpt_status_9_wd;
	// Trace: design.sv:54725:3
	wire intrpt_status_intrpt_status_9_we;
	// Trace: design.sv:54726:3
	wire intrpt_status_intrpt_status_9_re;
	// Trace: design.sv:54727:3
	wire intrpt_status_intrpt_status_10_qs;
	// Trace: design.sv:54728:3
	wire intrpt_status_intrpt_status_10_wd;
	// Trace: design.sv:54729:3
	wire intrpt_status_intrpt_status_10_we;
	// Trace: design.sv:54730:3
	wire intrpt_status_intrpt_status_10_re;
	// Trace: design.sv:54731:3
	wire intrpt_status_intrpt_status_11_qs;
	// Trace: design.sv:54732:3
	wire intrpt_status_intrpt_status_11_wd;
	// Trace: design.sv:54733:3
	wire intrpt_status_intrpt_status_11_we;
	// Trace: design.sv:54734:3
	wire intrpt_status_intrpt_status_11_re;
	// Trace: design.sv:54735:3
	wire intrpt_status_intrpt_status_12_qs;
	// Trace: design.sv:54736:3
	wire intrpt_status_intrpt_status_12_wd;
	// Trace: design.sv:54737:3
	wire intrpt_status_intrpt_status_12_we;
	// Trace: design.sv:54738:3
	wire intrpt_status_intrpt_status_12_re;
	// Trace: design.sv:54739:3
	wire intrpt_status_intrpt_status_13_qs;
	// Trace: design.sv:54740:3
	wire intrpt_status_intrpt_status_13_wd;
	// Trace: design.sv:54741:3
	wire intrpt_status_intrpt_status_13_we;
	// Trace: design.sv:54742:3
	wire intrpt_status_intrpt_status_13_re;
	// Trace: design.sv:54743:3
	wire intrpt_status_intrpt_status_14_qs;
	// Trace: design.sv:54744:3
	wire intrpt_status_intrpt_status_14_wd;
	// Trace: design.sv:54745:3
	wire intrpt_status_intrpt_status_14_we;
	// Trace: design.sv:54746:3
	wire intrpt_status_intrpt_status_14_re;
	// Trace: design.sv:54747:3
	wire intrpt_status_intrpt_status_15_qs;
	// Trace: design.sv:54748:3
	wire intrpt_status_intrpt_status_15_wd;
	// Trace: design.sv:54749:3
	wire intrpt_status_intrpt_status_15_we;
	// Trace: design.sv:54750:3
	wire intrpt_status_intrpt_status_15_re;
	// Trace: design.sv:54751:3
	wire intrpt_status_intrpt_status_16_qs;
	// Trace: design.sv:54752:3
	wire intrpt_status_intrpt_status_16_wd;
	// Trace: design.sv:54753:3
	wire intrpt_status_intrpt_status_16_we;
	// Trace: design.sv:54754:3
	wire intrpt_status_intrpt_status_16_re;
	// Trace: design.sv:54755:3
	wire intrpt_status_intrpt_status_17_qs;
	// Trace: design.sv:54756:3
	wire intrpt_status_intrpt_status_17_wd;
	// Trace: design.sv:54757:3
	wire intrpt_status_intrpt_status_17_we;
	// Trace: design.sv:54758:3
	wire intrpt_status_intrpt_status_17_re;
	// Trace: design.sv:54759:3
	wire intrpt_status_intrpt_status_18_qs;
	// Trace: design.sv:54760:3
	wire intrpt_status_intrpt_status_18_wd;
	// Trace: design.sv:54761:3
	wire intrpt_status_intrpt_status_18_we;
	// Trace: design.sv:54762:3
	wire intrpt_status_intrpt_status_18_re;
	// Trace: design.sv:54763:3
	wire intrpt_status_intrpt_status_19_qs;
	// Trace: design.sv:54764:3
	wire intrpt_status_intrpt_status_19_wd;
	// Trace: design.sv:54765:3
	wire intrpt_status_intrpt_status_19_we;
	// Trace: design.sv:54766:3
	wire intrpt_status_intrpt_status_19_re;
	// Trace: design.sv:54767:3
	wire intrpt_status_intrpt_status_20_qs;
	// Trace: design.sv:54768:3
	wire intrpt_status_intrpt_status_20_wd;
	// Trace: design.sv:54769:3
	wire intrpt_status_intrpt_status_20_we;
	// Trace: design.sv:54770:3
	wire intrpt_status_intrpt_status_20_re;
	// Trace: design.sv:54771:3
	wire intrpt_status_intrpt_status_21_qs;
	// Trace: design.sv:54772:3
	wire intrpt_status_intrpt_status_21_wd;
	// Trace: design.sv:54773:3
	wire intrpt_status_intrpt_status_21_we;
	// Trace: design.sv:54774:3
	wire intrpt_status_intrpt_status_21_re;
	// Trace: design.sv:54775:3
	wire intrpt_status_intrpt_status_22_qs;
	// Trace: design.sv:54776:3
	wire intrpt_status_intrpt_status_22_wd;
	// Trace: design.sv:54777:3
	wire intrpt_status_intrpt_status_22_we;
	// Trace: design.sv:54778:3
	wire intrpt_status_intrpt_status_22_re;
	// Trace: design.sv:54779:3
	wire intrpt_status_intrpt_status_23_qs;
	// Trace: design.sv:54780:3
	wire intrpt_status_intrpt_status_23_wd;
	// Trace: design.sv:54781:3
	wire intrpt_status_intrpt_status_23_we;
	// Trace: design.sv:54782:3
	wire intrpt_status_intrpt_status_23_re;
	// Trace: design.sv:54783:3
	wire intrpt_status_intrpt_status_24_qs;
	// Trace: design.sv:54784:3
	wire intrpt_status_intrpt_status_24_wd;
	// Trace: design.sv:54785:3
	wire intrpt_status_intrpt_status_24_we;
	// Trace: design.sv:54786:3
	wire intrpt_status_intrpt_status_24_re;
	// Trace: design.sv:54787:3
	wire intrpt_status_intrpt_status_25_qs;
	// Trace: design.sv:54788:3
	wire intrpt_status_intrpt_status_25_wd;
	// Trace: design.sv:54789:3
	wire intrpt_status_intrpt_status_25_we;
	// Trace: design.sv:54790:3
	wire intrpt_status_intrpt_status_25_re;
	// Trace: design.sv:54791:3
	wire intrpt_status_intrpt_status_26_qs;
	// Trace: design.sv:54792:3
	wire intrpt_status_intrpt_status_26_wd;
	// Trace: design.sv:54793:3
	wire intrpt_status_intrpt_status_26_we;
	// Trace: design.sv:54794:3
	wire intrpt_status_intrpt_status_26_re;
	// Trace: design.sv:54795:3
	wire intrpt_status_intrpt_status_27_qs;
	// Trace: design.sv:54796:3
	wire intrpt_status_intrpt_status_27_wd;
	// Trace: design.sv:54797:3
	wire intrpt_status_intrpt_status_27_we;
	// Trace: design.sv:54798:3
	wire intrpt_status_intrpt_status_27_re;
	// Trace: design.sv:54799:3
	wire intrpt_status_intrpt_status_28_qs;
	// Trace: design.sv:54800:3
	wire intrpt_status_intrpt_status_28_wd;
	// Trace: design.sv:54801:3
	wire intrpt_status_intrpt_status_28_we;
	// Trace: design.sv:54802:3
	wire intrpt_status_intrpt_status_28_re;
	// Trace: design.sv:54803:3
	wire intrpt_status_intrpt_status_29_qs;
	// Trace: design.sv:54804:3
	wire intrpt_status_intrpt_status_29_wd;
	// Trace: design.sv:54805:3
	wire intrpt_status_intrpt_status_29_we;
	// Trace: design.sv:54806:3
	wire intrpt_status_intrpt_status_29_re;
	// Trace: design.sv:54807:3
	wire intrpt_status_intrpt_status_30_qs;
	// Trace: design.sv:54808:3
	wire intrpt_status_intrpt_status_30_wd;
	// Trace: design.sv:54809:3
	wire intrpt_status_intrpt_status_30_we;
	// Trace: design.sv:54810:3
	wire intrpt_status_intrpt_status_30_re;
	// Trace: design.sv:54811:3
	wire intrpt_status_intrpt_status_31_qs;
	// Trace: design.sv:54812:3
	wire intrpt_status_intrpt_status_31_wd;
	// Trace: design.sv:54813:3
	wire intrpt_status_intrpt_status_31_we;
	// Trace: design.sv:54814:3
	wire intrpt_status_intrpt_status_31_re;
	// Trace: design.sv:54815:3
	wire intrpt_rise_status_intrpt_rise_status_0_qs;
	// Trace: design.sv:54816:3
	wire intrpt_rise_status_intrpt_rise_status_0_wd;
	// Trace: design.sv:54817:3
	wire intrpt_rise_status_intrpt_rise_status_0_we;
	// Trace: design.sv:54818:3
	wire intrpt_rise_status_intrpt_rise_status_1_qs;
	// Trace: design.sv:54819:3
	wire intrpt_rise_status_intrpt_rise_status_1_wd;
	// Trace: design.sv:54820:3
	wire intrpt_rise_status_intrpt_rise_status_1_we;
	// Trace: design.sv:54821:3
	wire intrpt_rise_status_intrpt_rise_status_2_qs;
	// Trace: design.sv:54822:3
	wire intrpt_rise_status_intrpt_rise_status_2_wd;
	// Trace: design.sv:54823:3
	wire intrpt_rise_status_intrpt_rise_status_2_we;
	// Trace: design.sv:54824:3
	wire intrpt_rise_status_intrpt_rise_status_3_qs;
	// Trace: design.sv:54825:3
	wire intrpt_rise_status_intrpt_rise_status_3_wd;
	// Trace: design.sv:54826:3
	wire intrpt_rise_status_intrpt_rise_status_3_we;
	// Trace: design.sv:54827:3
	wire intrpt_rise_status_intrpt_rise_status_4_qs;
	// Trace: design.sv:54828:3
	wire intrpt_rise_status_intrpt_rise_status_4_wd;
	// Trace: design.sv:54829:3
	wire intrpt_rise_status_intrpt_rise_status_4_we;
	// Trace: design.sv:54830:3
	wire intrpt_rise_status_intrpt_rise_status_5_qs;
	// Trace: design.sv:54831:3
	wire intrpt_rise_status_intrpt_rise_status_5_wd;
	// Trace: design.sv:54832:3
	wire intrpt_rise_status_intrpt_rise_status_5_we;
	// Trace: design.sv:54833:3
	wire intrpt_rise_status_intrpt_rise_status_6_qs;
	// Trace: design.sv:54834:3
	wire intrpt_rise_status_intrpt_rise_status_6_wd;
	// Trace: design.sv:54835:3
	wire intrpt_rise_status_intrpt_rise_status_6_we;
	// Trace: design.sv:54836:3
	wire intrpt_rise_status_intrpt_rise_status_7_qs;
	// Trace: design.sv:54837:3
	wire intrpt_rise_status_intrpt_rise_status_7_wd;
	// Trace: design.sv:54838:3
	wire intrpt_rise_status_intrpt_rise_status_7_we;
	// Trace: design.sv:54839:3
	wire intrpt_rise_status_intrpt_rise_status_8_qs;
	// Trace: design.sv:54840:3
	wire intrpt_rise_status_intrpt_rise_status_8_wd;
	// Trace: design.sv:54841:3
	wire intrpt_rise_status_intrpt_rise_status_8_we;
	// Trace: design.sv:54842:3
	wire intrpt_rise_status_intrpt_rise_status_9_qs;
	// Trace: design.sv:54843:3
	wire intrpt_rise_status_intrpt_rise_status_9_wd;
	// Trace: design.sv:54844:3
	wire intrpt_rise_status_intrpt_rise_status_9_we;
	// Trace: design.sv:54845:3
	wire intrpt_rise_status_intrpt_rise_status_10_qs;
	// Trace: design.sv:54846:3
	wire intrpt_rise_status_intrpt_rise_status_10_wd;
	// Trace: design.sv:54847:3
	wire intrpt_rise_status_intrpt_rise_status_10_we;
	// Trace: design.sv:54848:3
	wire intrpt_rise_status_intrpt_rise_status_11_qs;
	// Trace: design.sv:54849:3
	wire intrpt_rise_status_intrpt_rise_status_11_wd;
	// Trace: design.sv:54850:3
	wire intrpt_rise_status_intrpt_rise_status_11_we;
	// Trace: design.sv:54851:3
	wire intrpt_rise_status_intrpt_rise_status_12_qs;
	// Trace: design.sv:54852:3
	wire intrpt_rise_status_intrpt_rise_status_12_wd;
	// Trace: design.sv:54853:3
	wire intrpt_rise_status_intrpt_rise_status_12_we;
	// Trace: design.sv:54854:3
	wire intrpt_rise_status_intrpt_rise_status_13_qs;
	// Trace: design.sv:54855:3
	wire intrpt_rise_status_intrpt_rise_status_13_wd;
	// Trace: design.sv:54856:3
	wire intrpt_rise_status_intrpt_rise_status_13_we;
	// Trace: design.sv:54857:3
	wire intrpt_rise_status_intrpt_rise_status_14_qs;
	// Trace: design.sv:54858:3
	wire intrpt_rise_status_intrpt_rise_status_14_wd;
	// Trace: design.sv:54859:3
	wire intrpt_rise_status_intrpt_rise_status_14_we;
	// Trace: design.sv:54860:3
	wire intrpt_rise_status_intrpt_rise_status_15_qs;
	// Trace: design.sv:54861:3
	wire intrpt_rise_status_intrpt_rise_status_15_wd;
	// Trace: design.sv:54862:3
	wire intrpt_rise_status_intrpt_rise_status_15_we;
	// Trace: design.sv:54863:3
	wire intrpt_rise_status_intrpt_rise_status_16_qs;
	// Trace: design.sv:54864:3
	wire intrpt_rise_status_intrpt_rise_status_16_wd;
	// Trace: design.sv:54865:3
	wire intrpt_rise_status_intrpt_rise_status_16_we;
	// Trace: design.sv:54866:3
	wire intrpt_rise_status_intrpt_rise_status_17_qs;
	// Trace: design.sv:54867:3
	wire intrpt_rise_status_intrpt_rise_status_17_wd;
	// Trace: design.sv:54868:3
	wire intrpt_rise_status_intrpt_rise_status_17_we;
	// Trace: design.sv:54869:3
	wire intrpt_rise_status_intrpt_rise_status_18_qs;
	// Trace: design.sv:54870:3
	wire intrpt_rise_status_intrpt_rise_status_18_wd;
	// Trace: design.sv:54871:3
	wire intrpt_rise_status_intrpt_rise_status_18_we;
	// Trace: design.sv:54872:3
	wire intrpt_rise_status_intrpt_rise_status_19_qs;
	// Trace: design.sv:54873:3
	wire intrpt_rise_status_intrpt_rise_status_19_wd;
	// Trace: design.sv:54874:3
	wire intrpt_rise_status_intrpt_rise_status_19_we;
	// Trace: design.sv:54875:3
	wire intrpt_rise_status_intrpt_rise_status_20_qs;
	// Trace: design.sv:54876:3
	wire intrpt_rise_status_intrpt_rise_status_20_wd;
	// Trace: design.sv:54877:3
	wire intrpt_rise_status_intrpt_rise_status_20_we;
	// Trace: design.sv:54878:3
	wire intrpt_rise_status_intrpt_rise_status_21_qs;
	// Trace: design.sv:54879:3
	wire intrpt_rise_status_intrpt_rise_status_21_wd;
	// Trace: design.sv:54880:3
	wire intrpt_rise_status_intrpt_rise_status_21_we;
	// Trace: design.sv:54881:3
	wire intrpt_rise_status_intrpt_rise_status_22_qs;
	// Trace: design.sv:54882:3
	wire intrpt_rise_status_intrpt_rise_status_22_wd;
	// Trace: design.sv:54883:3
	wire intrpt_rise_status_intrpt_rise_status_22_we;
	// Trace: design.sv:54884:3
	wire intrpt_rise_status_intrpt_rise_status_23_qs;
	// Trace: design.sv:54885:3
	wire intrpt_rise_status_intrpt_rise_status_23_wd;
	// Trace: design.sv:54886:3
	wire intrpt_rise_status_intrpt_rise_status_23_we;
	// Trace: design.sv:54887:3
	wire intrpt_rise_status_intrpt_rise_status_24_qs;
	// Trace: design.sv:54888:3
	wire intrpt_rise_status_intrpt_rise_status_24_wd;
	// Trace: design.sv:54889:3
	wire intrpt_rise_status_intrpt_rise_status_24_we;
	// Trace: design.sv:54890:3
	wire intrpt_rise_status_intrpt_rise_status_25_qs;
	// Trace: design.sv:54891:3
	wire intrpt_rise_status_intrpt_rise_status_25_wd;
	// Trace: design.sv:54892:3
	wire intrpt_rise_status_intrpt_rise_status_25_we;
	// Trace: design.sv:54893:3
	wire intrpt_rise_status_intrpt_rise_status_26_qs;
	// Trace: design.sv:54894:3
	wire intrpt_rise_status_intrpt_rise_status_26_wd;
	// Trace: design.sv:54895:3
	wire intrpt_rise_status_intrpt_rise_status_26_we;
	// Trace: design.sv:54896:3
	wire intrpt_rise_status_intrpt_rise_status_27_qs;
	// Trace: design.sv:54897:3
	wire intrpt_rise_status_intrpt_rise_status_27_wd;
	// Trace: design.sv:54898:3
	wire intrpt_rise_status_intrpt_rise_status_27_we;
	// Trace: design.sv:54899:3
	wire intrpt_rise_status_intrpt_rise_status_28_qs;
	// Trace: design.sv:54900:3
	wire intrpt_rise_status_intrpt_rise_status_28_wd;
	// Trace: design.sv:54901:3
	wire intrpt_rise_status_intrpt_rise_status_28_we;
	// Trace: design.sv:54902:3
	wire intrpt_rise_status_intrpt_rise_status_29_qs;
	// Trace: design.sv:54903:3
	wire intrpt_rise_status_intrpt_rise_status_29_wd;
	// Trace: design.sv:54904:3
	wire intrpt_rise_status_intrpt_rise_status_29_we;
	// Trace: design.sv:54905:3
	wire intrpt_rise_status_intrpt_rise_status_30_qs;
	// Trace: design.sv:54906:3
	wire intrpt_rise_status_intrpt_rise_status_30_wd;
	// Trace: design.sv:54907:3
	wire intrpt_rise_status_intrpt_rise_status_30_we;
	// Trace: design.sv:54908:3
	wire intrpt_rise_status_intrpt_rise_status_31_qs;
	// Trace: design.sv:54909:3
	wire intrpt_rise_status_intrpt_rise_status_31_wd;
	// Trace: design.sv:54910:3
	wire intrpt_rise_status_intrpt_rise_status_31_we;
	// Trace: design.sv:54911:3
	wire intrpt_fall_status_intrpt_fall_status_0_qs;
	// Trace: design.sv:54912:3
	wire intrpt_fall_status_intrpt_fall_status_0_wd;
	// Trace: design.sv:54913:3
	wire intrpt_fall_status_intrpt_fall_status_0_we;
	// Trace: design.sv:54914:3
	wire intrpt_fall_status_intrpt_fall_status_1_qs;
	// Trace: design.sv:54915:3
	wire intrpt_fall_status_intrpt_fall_status_1_wd;
	// Trace: design.sv:54916:3
	wire intrpt_fall_status_intrpt_fall_status_1_we;
	// Trace: design.sv:54917:3
	wire intrpt_fall_status_intrpt_fall_status_2_qs;
	// Trace: design.sv:54918:3
	wire intrpt_fall_status_intrpt_fall_status_2_wd;
	// Trace: design.sv:54919:3
	wire intrpt_fall_status_intrpt_fall_status_2_we;
	// Trace: design.sv:54920:3
	wire intrpt_fall_status_intrpt_fall_status_3_qs;
	// Trace: design.sv:54921:3
	wire intrpt_fall_status_intrpt_fall_status_3_wd;
	// Trace: design.sv:54922:3
	wire intrpt_fall_status_intrpt_fall_status_3_we;
	// Trace: design.sv:54923:3
	wire intrpt_fall_status_intrpt_fall_status_4_qs;
	// Trace: design.sv:54924:3
	wire intrpt_fall_status_intrpt_fall_status_4_wd;
	// Trace: design.sv:54925:3
	wire intrpt_fall_status_intrpt_fall_status_4_we;
	// Trace: design.sv:54926:3
	wire intrpt_fall_status_intrpt_fall_status_5_qs;
	// Trace: design.sv:54927:3
	wire intrpt_fall_status_intrpt_fall_status_5_wd;
	// Trace: design.sv:54928:3
	wire intrpt_fall_status_intrpt_fall_status_5_we;
	// Trace: design.sv:54929:3
	wire intrpt_fall_status_intrpt_fall_status_6_qs;
	// Trace: design.sv:54930:3
	wire intrpt_fall_status_intrpt_fall_status_6_wd;
	// Trace: design.sv:54931:3
	wire intrpt_fall_status_intrpt_fall_status_6_we;
	// Trace: design.sv:54932:3
	wire intrpt_fall_status_intrpt_fall_status_7_qs;
	// Trace: design.sv:54933:3
	wire intrpt_fall_status_intrpt_fall_status_7_wd;
	// Trace: design.sv:54934:3
	wire intrpt_fall_status_intrpt_fall_status_7_we;
	// Trace: design.sv:54935:3
	wire intrpt_fall_status_intrpt_fall_status_8_qs;
	// Trace: design.sv:54936:3
	wire intrpt_fall_status_intrpt_fall_status_8_wd;
	// Trace: design.sv:54937:3
	wire intrpt_fall_status_intrpt_fall_status_8_we;
	// Trace: design.sv:54938:3
	wire intrpt_fall_status_intrpt_fall_status_9_qs;
	// Trace: design.sv:54939:3
	wire intrpt_fall_status_intrpt_fall_status_9_wd;
	// Trace: design.sv:54940:3
	wire intrpt_fall_status_intrpt_fall_status_9_we;
	// Trace: design.sv:54941:3
	wire intrpt_fall_status_intrpt_fall_status_10_qs;
	// Trace: design.sv:54942:3
	wire intrpt_fall_status_intrpt_fall_status_10_wd;
	// Trace: design.sv:54943:3
	wire intrpt_fall_status_intrpt_fall_status_10_we;
	// Trace: design.sv:54944:3
	wire intrpt_fall_status_intrpt_fall_status_11_qs;
	// Trace: design.sv:54945:3
	wire intrpt_fall_status_intrpt_fall_status_11_wd;
	// Trace: design.sv:54946:3
	wire intrpt_fall_status_intrpt_fall_status_11_we;
	// Trace: design.sv:54947:3
	wire intrpt_fall_status_intrpt_fall_status_12_qs;
	// Trace: design.sv:54948:3
	wire intrpt_fall_status_intrpt_fall_status_12_wd;
	// Trace: design.sv:54949:3
	wire intrpt_fall_status_intrpt_fall_status_12_we;
	// Trace: design.sv:54950:3
	wire intrpt_fall_status_intrpt_fall_status_13_qs;
	// Trace: design.sv:54951:3
	wire intrpt_fall_status_intrpt_fall_status_13_wd;
	// Trace: design.sv:54952:3
	wire intrpt_fall_status_intrpt_fall_status_13_we;
	// Trace: design.sv:54953:3
	wire intrpt_fall_status_intrpt_fall_status_14_qs;
	// Trace: design.sv:54954:3
	wire intrpt_fall_status_intrpt_fall_status_14_wd;
	// Trace: design.sv:54955:3
	wire intrpt_fall_status_intrpt_fall_status_14_we;
	// Trace: design.sv:54956:3
	wire intrpt_fall_status_intrpt_fall_status_15_qs;
	// Trace: design.sv:54957:3
	wire intrpt_fall_status_intrpt_fall_status_15_wd;
	// Trace: design.sv:54958:3
	wire intrpt_fall_status_intrpt_fall_status_15_we;
	// Trace: design.sv:54959:3
	wire intrpt_fall_status_intrpt_fall_status_16_qs;
	// Trace: design.sv:54960:3
	wire intrpt_fall_status_intrpt_fall_status_16_wd;
	// Trace: design.sv:54961:3
	wire intrpt_fall_status_intrpt_fall_status_16_we;
	// Trace: design.sv:54962:3
	wire intrpt_fall_status_intrpt_fall_status_17_qs;
	// Trace: design.sv:54963:3
	wire intrpt_fall_status_intrpt_fall_status_17_wd;
	// Trace: design.sv:54964:3
	wire intrpt_fall_status_intrpt_fall_status_17_we;
	// Trace: design.sv:54965:3
	wire intrpt_fall_status_intrpt_fall_status_18_qs;
	// Trace: design.sv:54966:3
	wire intrpt_fall_status_intrpt_fall_status_18_wd;
	// Trace: design.sv:54967:3
	wire intrpt_fall_status_intrpt_fall_status_18_we;
	// Trace: design.sv:54968:3
	wire intrpt_fall_status_intrpt_fall_status_19_qs;
	// Trace: design.sv:54969:3
	wire intrpt_fall_status_intrpt_fall_status_19_wd;
	// Trace: design.sv:54970:3
	wire intrpt_fall_status_intrpt_fall_status_19_we;
	// Trace: design.sv:54971:3
	wire intrpt_fall_status_intrpt_fall_status_20_qs;
	// Trace: design.sv:54972:3
	wire intrpt_fall_status_intrpt_fall_status_20_wd;
	// Trace: design.sv:54973:3
	wire intrpt_fall_status_intrpt_fall_status_20_we;
	// Trace: design.sv:54974:3
	wire intrpt_fall_status_intrpt_fall_status_21_qs;
	// Trace: design.sv:54975:3
	wire intrpt_fall_status_intrpt_fall_status_21_wd;
	// Trace: design.sv:54976:3
	wire intrpt_fall_status_intrpt_fall_status_21_we;
	// Trace: design.sv:54977:3
	wire intrpt_fall_status_intrpt_fall_status_22_qs;
	// Trace: design.sv:54978:3
	wire intrpt_fall_status_intrpt_fall_status_22_wd;
	// Trace: design.sv:54979:3
	wire intrpt_fall_status_intrpt_fall_status_22_we;
	// Trace: design.sv:54980:3
	wire intrpt_fall_status_intrpt_fall_status_23_qs;
	// Trace: design.sv:54981:3
	wire intrpt_fall_status_intrpt_fall_status_23_wd;
	// Trace: design.sv:54982:3
	wire intrpt_fall_status_intrpt_fall_status_23_we;
	// Trace: design.sv:54983:3
	wire intrpt_fall_status_intrpt_fall_status_24_qs;
	// Trace: design.sv:54984:3
	wire intrpt_fall_status_intrpt_fall_status_24_wd;
	// Trace: design.sv:54985:3
	wire intrpt_fall_status_intrpt_fall_status_24_we;
	// Trace: design.sv:54986:3
	wire intrpt_fall_status_intrpt_fall_status_25_qs;
	// Trace: design.sv:54987:3
	wire intrpt_fall_status_intrpt_fall_status_25_wd;
	// Trace: design.sv:54988:3
	wire intrpt_fall_status_intrpt_fall_status_25_we;
	// Trace: design.sv:54989:3
	wire intrpt_fall_status_intrpt_fall_status_26_qs;
	// Trace: design.sv:54990:3
	wire intrpt_fall_status_intrpt_fall_status_26_wd;
	// Trace: design.sv:54991:3
	wire intrpt_fall_status_intrpt_fall_status_26_we;
	// Trace: design.sv:54992:3
	wire intrpt_fall_status_intrpt_fall_status_27_qs;
	// Trace: design.sv:54993:3
	wire intrpt_fall_status_intrpt_fall_status_27_wd;
	// Trace: design.sv:54994:3
	wire intrpt_fall_status_intrpt_fall_status_27_we;
	// Trace: design.sv:54995:3
	wire intrpt_fall_status_intrpt_fall_status_28_qs;
	// Trace: design.sv:54996:3
	wire intrpt_fall_status_intrpt_fall_status_28_wd;
	// Trace: design.sv:54997:3
	wire intrpt_fall_status_intrpt_fall_status_28_we;
	// Trace: design.sv:54998:3
	wire intrpt_fall_status_intrpt_fall_status_29_qs;
	// Trace: design.sv:54999:3
	wire intrpt_fall_status_intrpt_fall_status_29_wd;
	// Trace: design.sv:55000:3
	wire intrpt_fall_status_intrpt_fall_status_29_we;
	// Trace: design.sv:55001:3
	wire intrpt_fall_status_intrpt_fall_status_30_qs;
	// Trace: design.sv:55002:3
	wire intrpt_fall_status_intrpt_fall_status_30_wd;
	// Trace: design.sv:55003:3
	wire intrpt_fall_status_intrpt_fall_status_30_we;
	// Trace: design.sv:55004:3
	wire intrpt_fall_status_intrpt_fall_status_31_qs;
	// Trace: design.sv:55005:3
	wire intrpt_fall_status_intrpt_fall_status_31_wd;
	// Trace: design.sv:55006:3
	wire intrpt_fall_status_intrpt_fall_status_31_we;
	// Trace: design.sv:55007:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_0_qs;
	// Trace: design.sv:55008:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_0_wd;
	// Trace: design.sv:55009:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_0_we;
	// Trace: design.sv:55010:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_1_qs;
	// Trace: design.sv:55011:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_1_wd;
	// Trace: design.sv:55012:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_1_we;
	// Trace: design.sv:55013:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_2_qs;
	// Trace: design.sv:55014:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_2_wd;
	// Trace: design.sv:55015:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_2_we;
	// Trace: design.sv:55016:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_3_qs;
	// Trace: design.sv:55017:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_3_wd;
	// Trace: design.sv:55018:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_3_we;
	// Trace: design.sv:55019:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_4_qs;
	// Trace: design.sv:55020:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_4_wd;
	// Trace: design.sv:55021:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_4_we;
	// Trace: design.sv:55022:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_5_qs;
	// Trace: design.sv:55023:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_5_wd;
	// Trace: design.sv:55024:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_5_we;
	// Trace: design.sv:55025:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_6_qs;
	// Trace: design.sv:55026:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_6_wd;
	// Trace: design.sv:55027:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_6_we;
	// Trace: design.sv:55028:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_7_qs;
	// Trace: design.sv:55029:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_7_wd;
	// Trace: design.sv:55030:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_7_we;
	// Trace: design.sv:55031:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_8_qs;
	// Trace: design.sv:55032:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_8_wd;
	// Trace: design.sv:55033:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_8_we;
	// Trace: design.sv:55034:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_9_qs;
	// Trace: design.sv:55035:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_9_wd;
	// Trace: design.sv:55036:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_9_we;
	// Trace: design.sv:55037:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_10_qs;
	// Trace: design.sv:55038:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_10_wd;
	// Trace: design.sv:55039:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_10_we;
	// Trace: design.sv:55040:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_11_qs;
	// Trace: design.sv:55041:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_11_wd;
	// Trace: design.sv:55042:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_11_we;
	// Trace: design.sv:55043:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_12_qs;
	// Trace: design.sv:55044:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_12_wd;
	// Trace: design.sv:55045:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_12_we;
	// Trace: design.sv:55046:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_13_qs;
	// Trace: design.sv:55047:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_13_wd;
	// Trace: design.sv:55048:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_13_we;
	// Trace: design.sv:55049:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_14_qs;
	// Trace: design.sv:55050:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_14_wd;
	// Trace: design.sv:55051:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_14_we;
	// Trace: design.sv:55052:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_15_qs;
	// Trace: design.sv:55053:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_15_wd;
	// Trace: design.sv:55054:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_15_we;
	// Trace: design.sv:55055:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_16_qs;
	// Trace: design.sv:55056:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_16_wd;
	// Trace: design.sv:55057:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_16_we;
	// Trace: design.sv:55058:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_17_qs;
	// Trace: design.sv:55059:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_17_wd;
	// Trace: design.sv:55060:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_17_we;
	// Trace: design.sv:55061:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_18_qs;
	// Trace: design.sv:55062:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_18_wd;
	// Trace: design.sv:55063:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_18_we;
	// Trace: design.sv:55064:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_19_qs;
	// Trace: design.sv:55065:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_19_wd;
	// Trace: design.sv:55066:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_19_we;
	// Trace: design.sv:55067:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_20_qs;
	// Trace: design.sv:55068:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_20_wd;
	// Trace: design.sv:55069:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_20_we;
	// Trace: design.sv:55070:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_21_qs;
	// Trace: design.sv:55071:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_21_wd;
	// Trace: design.sv:55072:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_21_we;
	// Trace: design.sv:55073:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_22_qs;
	// Trace: design.sv:55074:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_22_wd;
	// Trace: design.sv:55075:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_22_we;
	// Trace: design.sv:55076:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_23_qs;
	// Trace: design.sv:55077:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_23_wd;
	// Trace: design.sv:55078:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_23_we;
	// Trace: design.sv:55079:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_24_qs;
	// Trace: design.sv:55080:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_24_wd;
	// Trace: design.sv:55081:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_24_we;
	// Trace: design.sv:55082:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_25_qs;
	// Trace: design.sv:55083:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_25_wd;
	// Trace: design.sv:55084:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_25_we;
	// Trace: design.sv:55085:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_26_qs;
	// Trace: design.sv:55086:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_26_wd;
	// Trace: design.sv:55087:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_26_we;
	// Trace: design.sv:55088:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_27_qs;
	// Trace: design.sv:55089:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_27_wd;
	// Trace: design.sv:55090:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_27_we;
	// Trace: design.sv:55091:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_28_qs;
	// Trace: design.sv:55092:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_28_wd;
	// Trace: design.sv:55093:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_28_we;
	// Trace: design.sv:55094:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_29_qs;
	// Trace: design.sv:55095:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_29_wd;
	// Trace: design.sv:55096:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_29_we;
	// Trace: design.sv:55097:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_30_qs;
	// Trace: design.sv:55098:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_30_wd;
	// Trace: design.sv:55099:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_30_we;
	// Trace: design.sv:55100:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_31_qs;
	// Trace: design.sv:55101:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_31_wd;
	// Trace: design.sv:55102:3
	wire intrpt_lvl_high_status_intrpt_lvl_high_status_31_we;
	// Trace: design.sv:55103:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_0_qs;
	// Trace: design.sv:55104:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_0_wd;
	// Trace: design.sv:55105:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_0_we;
	// Trace: design.sv:55106:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_1_qs;
	// Trace: design.sv:55107:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_1_wd;
	// Trace: design.sv:55108:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_1_we;
	// Trace: design.sv:55109:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_2_qs;
	// Trace: design.sv:55110:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_2_wd;
	// Trace: design.sv:55111:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_2_we;
	// Trace: design.sv:55112:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_3_qs;
	// Trace: design.sv:55113:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_3_wd;
	// Trace: design.sv:55114:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_3_we;
	// Trace: design.sv:55115:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_4_qs;
	// Trace: design.sv:55116:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_4_wd;
	// Trace: design.sv:55117:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_4_we;
	// Trace: design.sv:55118:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_5_qs;
	// Trace: design.sv:55119:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_5_wd;
	// Trace: design.sv:55120:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_5_we;
	// Trace: design.sv:55121:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_6_qs;
	// Trace: design.sv:55122:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_6_wd;
	// Trace: design.sv:55123:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_6_we;
	// Trace: design.sv:55124:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_7_qs;
	// Trace: design.sv:55125:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_7_wd;
	// Trace: design.sv:55126:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_7_we;
	// Trace: design.sv:55127:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_8_qs;
	// Trace: design.sv:55128:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_8_wd;
	// Trace: design.sv:55129:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_8_we;
	// Trace: design.sv:55130:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_9_qs;
	// Trace: design.sv:55131:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_9_wd;
	// Trace: design.sv:55132:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_9_we;
	// Trace: design.sv:55133:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_10_qs;
	// Trace: design.sv:55134:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_10_wd;
	// Trace: design.sv:55135:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_10_we;
	// Trace: design.sv:55136:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_11_qs;
	// Trace: design.sv:55137:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_11_wd;
	// Trace: design.sv:55138:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_11_we;
	// Trace: design.sv:55139:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_12_qs;
	// Trace: design.sv:55140:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_12_wd;
	// Trace: design.sv:55141:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_12_we;
	// Trace: design.sv:55142:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_13_qs;
	// Trace: design.sv:55143:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_13_wd;
	// Trace: design.sv:55144:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_13_we;
	// Trace: design.sv:55145:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_14_qs;
	// Trace: design.sv:55146:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_14_wd;
	// Trace: design.sv:55147:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_14_we;
	// Trace: design.sv:55148:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_15_qs;
	// Trace: design.sv:55149:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_15_wd;
	// Trace: design.sv:55150:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_15_we;
	// Trace: design.sv:55151:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_16_qs;
	// Trace: design.sv:55152:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_16_wd;
	// Trace: design.sv:55153:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_16_we;
	// Trace: design.sv:55154:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_17_qs;
	// Trace: design.sv:55155:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_17_wd;
	// Trace: design.sv:55156:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_17_we;
	// Trace: design.sv:55157:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_18_qs;
	// Trace: design.sv:55158:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_18_wd;
	// Trace: design.sv:55159:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_18_we;
	// Trace: design.sv:55160:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_19_qs;
	// Trace: design.sv:55161:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_19_wd;
	// Trace: design.sv:55162:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_19_we;
	// Trace: design.sv:55163:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_20_qs;
	// Trace: design.sv:55164:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_20_wd;
	// Trace: design.sv:55165:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_20_we;
	// Trace: design.sv:55166:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_21_qs;
	// Trace: design.sv:55167:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_21_wd;
	// Trace: design.sv:55168:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_21_we;
	// Trace: design.sv:55169:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_22_qs;
	// Trace: design.sv:55170:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_22_wd;
	// Trace: design.sv:55171:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_22_we;
	// Trace: design.sv:55172:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_23_qs;
	// Trace: design.sv:55173:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_23_wd;
	// Trace: design.sv:55174:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_23_we;
	// Trace: design.sv:55175:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_24_qs;
	// Trace: design.sv:55176:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_24_wd;
	// Trace: design.sv:55177:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_24_we;
	// Trace: design.sv:55178:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_25_qs;
	// Trace: design.sv:55179:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_25_wd;
	// Trace: design.sv:55180:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_25_we;
	// Trace: design.sv:55181:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_26_qs;
	// Trace: design.sv:55182:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_26_wd;
	// Trace: design.sv:55183:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_26_we;
	// Trace: design.sv:55184:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_27_qs;
	// Trace: design.sv:55185:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_27_wd;
	// Trace: design.sv:55186:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_27_we;
	// Trace: design.sv:55187:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_28_qs;
	// Trace: design.sv:55188:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_28_wd;
	// Trace: design.sv:55189:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_28_we;
	// Trace: design.sv:55190:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_29_qs;
	// Trace: design.sv:55191:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_29_wd;
	// Trace: design.sv:55192:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_29_we;
	// Trace: design.sv:55193:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_30_qs;
	// Trace: design.sv:55194:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_30_wd;
	// Trace: design.sv:55195:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_30_we;
	// Trace: design.sv:55196:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_31_qs;
	// Trace: design.sv:55197:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_31_wd;
	// Trace: design.sv:55198:3
	wire intrpt_lvl_low_status_intrpt_lvl_low_status_31_we;
	// Trace: design.sv:55204:3
	localparam [31:0] sv2v_uu_u_info_gpio_cnt_DW = 10;
	// removed localparam type sv2v_uu_u_info_gpio_cnt_wd
	localparam [9:0] sv2v_uu_u_info_gpio_cnt_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(10)) u_info_gpio_cnt(
		.re(info_gpio_cnt_re),
		.we(1'b0),
		.wd(sv2v_uu_u_info_gpio_cnt_ext_wd_0),
		.d(hw2reg[403-:10]),
		.qre(),
		.qe(),
		.q(),
		.qs(info_gpio_cnt_qs)
	);
	// Trace: design.sv:55219:3
	localparam [31:0] sv2v_uu_u_info_version_DW = 10;
	// removed localparam type sv2v_uu_u_info_version_wd
	localparam [9:0] sv2v_uu_u_info_version_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(10)) u_info_version(
		.re(info_version_re),
		.we(1'b0),
		.wd(sv2v_uu_u_info_version_ext_wd_0),
		.d(hw2reg[393-:10]),
		.qre(),
		.qe(),
		.q(),
		.qs(info_version_qs)
	);
	// Trace: design.sv:55236:3
	localparam signed [31:0] sv2v_uu_u_cfg_glbl_intrpt_mode_DW = 1;
	// removed localparam type sv2v_uu_u_cfg_glbl_intrpt_mode_d
	localparam [0:0] sv2v_uu_u_cfg_glbl_intrpt_mode_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cfg_glbl_intrpt_mode(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cfg_glbl_intrpt_mode_we),
		.wd(cfg_glbl_intrpt_mode_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cfg_glbl_intrpt_mode_ext_d_0),
		.qe(),
		.q(reg2hw[642]),
		.qs(cfg_glbl_intrpt_mode_qs)
	);
	// Trace: design.sv:55262:3
	localparam signed [31:0] sv2v_uu_u_cfg_pin_lvl_intrpt_mode_DW = 1;
	// removed localparam type sv2v_uu_u_cfg_pin_lvl_intrpt_mode_d
	localparam [0:0] sv2v_uu_u_cfg_pin_lvl_intrpt_mode_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cfg_pin_lvl_intrpt_mode(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cfg_pin_lvl_intrpt_mode_we),
		.wd(cfg_pin_lvl_intrpt_mode_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cfg_pin_lvl_intrpt_mode_ext_d_0),
		.qe(),
		.q(reg2hw[641]),
		.qs(cfg_pin_lvl_intrpt_mode_qs)
	);
	// Trace: design.sv:55288:3
	localparam signed [31:0] sv2v_uu_u_cfg_reserved_DW = 1;
	// removed localparam type sv2v_uu_u_cfg_reserved_d
	localparam [0:0] sv2v_uu_u_cfg_reserved_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cfg_reserved(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cfg_reserved_we),
		.wd(cfg_reserved_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cfg_reserved_ext_d_0),
		.qe(),
		.q(reg2hw[640]),
		.qs(cfg_reserved_qs)
	);
	// Trace: design.sv:55318:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_0_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_0_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_0_we),
		.wd(gpio_mode_0_mode_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_0_ext_d_0),
		.qe(),
		.q(reg2hw[577-:2]),
		.qs(gpio_mode_0_mode_0_qs)
	);
	// Trace: design.sv:55344:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_1_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_1_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_1_we),
		.wd(gpio_mode_0_mode_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_1_ext_d_0),
		.qe(),
		.q(reg2hw[579-:2]),
		.qs(gpio_mode_0_mode_1_qs)
	);
	// Trace: design.sv:55370:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_2_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_2_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_2_we),
		.wd(gpio_mode_0_mode_2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_2_ext_d_0),
		.qe(),
		.q(reg2hw[581-:2]),
		.qs(gpio_mode_0_mode_2_qs)
	);
	// Trace: design.sv:55396:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_3_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_3_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_3_we),
		.wd(gpio_mode_0_mode_3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_3_ext_d_0),
		.qe(),
		.q(reg2hw[583-:2]),
		.qs(gpio_mode_0_mode_3_qs)
	);
	// Trace: design.sv:55422:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_4_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_4_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_4_we),
		.wd(gpio_mode_0_mode_4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_4_ext_d_0),
		.qe(),
		.q(reg2hw[585-:2]),
		.qs(gpio_mode_0_mode_4_qs)
	);
	// Trace: design.sv:55448:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_5_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_5_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_5_we),
		.wd(gpio_mode_0_mode_5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_5_ext_d_0),
		.qe(),
		.q(reg2hw[587-:2]),
		.qs(gpio_mode_0_mode_5_qs)
	);
	// Trace: design.sv:55474:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_6_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_6_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_6_we),
		.wd(gpio_mode_0_mode_6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_6_ext_d_0),
		.qe(),
		.q(reg2hw[589-:2]),
		.qs(gpio_mode_0_mode_6_qs)
	);
	// Trace: design.sv:55500:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_7_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_7_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_7_we),
		.wd(gpio_mode_0_mode_7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_7_ext_d_0),
		.qe(),
		.q(reg2hw[591-:2]),
		.qs(gpio_mode_0_mode_7_qs)
	);
	// Trace: design.sv:55526:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_8_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_8_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_8_we),
		.wd(gpio_mode_0_mode_8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_8_ext_d_0),
		.qe(),
		.q(reg2hw[593-:2]),
		.qs(gpio_mode_0_mode_8_qs)
	);
	// Trace: design.sv:55552:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_9_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_9_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_9_we),
		.wd(gpio_mode_0_mode_9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_9_ext_d_0),
		.qe(),
		.q(reg2hw[595-:2]),
		.qs(gpio_mode_0_mode_9_qs)
	);
	// Trace: design.sv:55578:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_10_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_10_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_10_we),
		.wd(gpio_mode_0_mode_10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_10_ext_d_0),
		.qe(),
		.q(reg2hw[597-:2]),
		.qs(gpio_mode_0_mode_10_qs)
	);
	// Trace: design.sv:55604:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_11_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_11_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_11_we),
		.wd(gpio_mode_0_mode_11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_11_ext_d_0),
		.qe(),
		.q(reg2hw[599-:2]),
		.qs(gpio_mode_0_mode_11_qs)
	);
	// Trace: design.sv:55630:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_12_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_12_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_12_we),
		.wd(gpio_mode_0_mode_12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_12_ext_d_0),
		.qe(),
		.q(reg2hw[601-:2]),
		.qs(gpio_mode_0_mode_12_qs)
	);
	// Trace: design.sv:55656:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_13_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_13_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_13_we),
		.wd(gpio_mode_0_mode_13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_13_ext_d_0),
		.qe(),
		.q(reg2hw[603-:2]),
		.qs(gpio_mode_0_mode_13_qs)
	);
	// Trace: design.sv:55682:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_14_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_14_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_14_we),
		.wd(gpio_mode_0_mode_14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_14_ext_d_0),
		.qe(),
		.q(reg2hw[605-:2]),
		.qs(gpio_mode_0_mode_14_qs)
	);
	// Trace: design.sv:55708:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_0_mode_15_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_0_mode_15_d
	localparam [1:0] sv2v_uu_u_gpio_mode_0_mode_15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_0_mode_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_0_mode_15_we),
		.wd(gpio_mode_0_mode_15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_0_mode_15_ext_d_0),
		.qe(),
		.q(reg2hw[607-:2]),
		.qs(gpio_mode_0_mode_15_qs)
	);
	// Trace: design.sv:55737:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_16_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_16_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_16_we),
		.wd(gpio_mode_1_mode_16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_16_ext_d_0),
		.qe(),
		.q(reg2hw[609-:2]),
		.qs(gpio_mode_1_mode_16_qs)
	);
	// Trace: design.sv:55763:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_17_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_17_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_17_we),
		.wd(gpio_mode_1_mode_17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_17_ext_d_0),
		.qe(),
		.q(reg2hw[611-:2]),
		.qs(gpio_mode_1_mode_17_qs)
	);
	// Trace: design.sv:55789:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_18_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_18_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_18_we),
		.wd(gpio_mode_1_mode_18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_18_ext_d_0),
		.qe(),
		.q(reg2hw[613-:2]),
		.qs(gpio_mode_1_mode_18_qs)
	);
	// Trace: design.sv:55815:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_19_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_19_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_19_we),
		.wd(gpio_mode_1_mode_19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_19_ext_d_0),
		.qe(),
		.q(reg2hw[615-:2]),
		.qs(gpio_mode_1_mode_19_qs)
	);
	// Trace: design.sv:55841:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_20_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_20_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_20_we),
		.wd(gpio_mode_1_mode_20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_20_ext_d_0),
		.qe(),
		.q(reg2hw[617-:2]),
		.qs(gpio_mode_1_mode_20_qs)
	);
	// Trace: design.sv:55867:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_21_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_21_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_21_we),
		.wd(gpio_mode_1_mode_21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_21_ext_d_0),
		.qe(),
		.q(reg2hw[619-:2]),
		.qs(gpio_mode_1_mode_21_qs)
	);
	// Trace: design.sv:55893:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_22_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_22_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_22_we),
		.wd(gpio_mode_1_mode_22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_22_ext_d_0),
		.qe(),
		.q(reg2hw[621-:2]),
		.qs(gpio_mode_1_mode_22_qs)
	);
	// Trace: design.sv:55919:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_23_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_23_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_23_we),
		.wd(gpio_mode_1_mode_23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_23_ext_d_0),
		.qe(),
		.q(reg2hw[623-:2]),
		.qs(gpio_mode_1_mode_23_qs)
	);
	// Trace: design.sv:55945:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_24_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_24_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_24_we),
		.wd(gpio_mode_1_mode_24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_24_ext_d_0),
		.qe(),
		.q(reg2hw[625-:2]),
		.qs(gpio_mode_1_mode_24_qs)
	);
	// Trace: design.sv:55971:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_25_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_25_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_25_we),
		.wd(gpio_mode_1_mode_25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_25_ext_d_0),
		.qe(),
		.q(reg2hw[627-:2]),
		.qs(gpio_mode_1_mode_25_qs)
	);
	// Trace: design.sv:55997:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_26_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_26_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_26_we),
		.wd(gpio_mode_1_mode_26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_26_ext_d_0),
		.qe(),
		.q(reg2hw[629-:2]),
		.qs(gpio_mode_1_mode_26_qs)
	);
	// Trace: design.sv:56023:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_27_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_27_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_27_we),
		.wd(gpio_mode_1_mode_27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_27_ext_d_0),
		.qe(),
		.q(reg2hw[631-:2]),
		.qs(gpio_mode_1_mode_27_qs)
	);
	// Trace: design.sv:56049:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_28_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_28_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_28_we),
		.wd(gpio_mode_1_mode_28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_28_ext_d_0),
		.qe(),
		.q(reg2hw[633-:2]),
		.qs(gpio_mode_1_mode_28_qs)
	);
	// Trace: design.sv:56075:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_29_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_29_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_29_we),
		.wd(gpio_mode_1_mode_29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_29_ext_d_0),
		.qe(),
		.q(reg2hw[635-:2]),
		.qs(gpio_mode_1_mode_29_qs)
	);
	// Trace: design.sv:56101:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_30_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_30_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_30_we),
		.wd(gpio_mode_1_mode_30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_30_ext_d_0),
		.qe(),
		.q(reg2hw[637-:2]),
		.qs(gpio_mode_1_mode_30_qs)
	);
	// Trace: design.sv:56127:3
	localparam signed [31:0] sv2v_uu_u_gpio_mode_1_mode_31_DW = 2;
	// removed localparam type sv2v_uu_u_gpio_mode_1_mode_31_d
	localparam [1:0] sv2v_uu_u_gpio_mode_1_mode_31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_gpio_mode_1_mode_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_mode_1_mode_31_we),
		.wd(gpio_mode_1_mode_31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_mode_1_mode_31_ext_d_0),
		.qe(),
		.q(reg2hw[639-:2]),
		.qs(gpio_mode_1_mode_31_qs)
	);
	// Trace: design.sv:56158:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_0_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_0_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_0_we),
		.wd(gpio_en_gpio_en_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_0_ext_d_0),
		.qe(),
		.q(reg2hw[544]),
		.qs(gpio_en_gpio_en_0_qs)
	);
	// Trace: design.sv:56184:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_1_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_1_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_1_we),
		.wd(gpio_en_gpio_en_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_1_ext_d_0),
		.qe(),
		.q(reg2hw[545]),
		.qs(gpio_en_gpio_en_1_qs)
	);
	// Trace: design.sv:56210:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_2_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_2_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_2_we),
		.wd(gpio_en_gpio_en_2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_2_ext_d_0),
		.qe(),
		.q(reg2hw[546]),
		.qs(gpio_en_gpio_en_2_qs)
	);
	// Trace: design.sv:56236:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_3_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_3_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_3_we),
		.wd(gpio_en_gpio_en_3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_3_ext_d_0),
		.qe(),
		.q(reg2hw[547]),
		.qs(gpio_en_gpio_en_3_qs)
	);
	// Trace: design.sv:56262:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_4_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_4_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_4_we),
		.wd(gpio_en_gpio_en_4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_4_ext_d_0),
		.qe(),
		.q(reg2hw[548]),
		.qs(gpio_en_gpio_en_4_qs)
	);
	// Trace: design.sv:56288:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_5_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_5_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_5_we),
		.wd(gpio_en_gpio_en_5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_5_ext_d_0),
		.qe(),
		.q(reg2hw[549]),
		.qs(gpio_en_gpio_en_5_qs)
	);
	// Trace: design.sv:56314:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_6_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_6_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_6_we),
		.wd(gpio_en_gpio_en_6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_6_ext_d_0),
		.qe(),
		.q(reg2hw[550]),
		.qs(gpio_en_gpio_en_6_qs)
	);
	// Trace: design.sv:56340:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_7_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_7_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_7_we),
		.wd(gpio_en_gpio_en_7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_7_ext_d_0),
		.qe(),
		.q(reg2hw[551]),
		.qs(gpio_en_gpio_en_7_qs)
	);
	// Trace: design.sv:56366:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_8_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_8_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_8_we),
		.wd(gpio_en_gpio_en_8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_8_ext_d_0),
		.qe(),
		.q(reg2hw[552]),
		.qs(gpio_en_gpio_en_8_qs)
	);
	// Trace: design.sv:56392:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_9_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_9_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_9_we),
		.wd(gpio_en_gpio_en_9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_9_ext_d_0),
		.qe(),
		.q(reg2hw[553]),
		.qs(gpio_en_gpio_en_9_qs)
	);
	// Trace: design.sv:56418:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_10_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_10_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_10_we),
		.wd(gpio_en_gpio_en_10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_10_ext_d_0),
		.qe(),
		.q(reg2hw[554]),
		.qs(gpio_en_gpio_en_10_qs)
	);
	// Trace: design.sv:56444:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_11_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_11_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_11_we),
		.wd(gpio_en_gpio_en_11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_11_ext_d_0),
		.qe(),
		.q(reg2hw[555]),
		.qs(gpio_en_gpio_en_11_qs)
	);
	// Trace: design.sv:56470:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_12_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_12_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_12_we),
		.wd(gpio_en_gpio_en_12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_12_ext_d_0),
		.qe(),
		.q(reg2hw[556]),
		.qs(gpio_en_gpio_en_12_qs)
	);
	// Trace: design.sv:56496:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_13_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_13_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_13_we),
		.wd(gpio_en_gpio_en_13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_13_ext_d_0),
		.qe(),
		.q(reg2hw[557]),
		.qs(gpio_en_gpio_en_13_qs)
	);
	// Trace: design.sv:56522:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_14_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_14_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_14_we),
		.wd(gpio_en_gpio_en_14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_14_ext_d_0),
		.qe(),
		.q(reg2hw[558]),
		.qs(gpio_en_gpio_en_14_qs)
	);
	// Trace: design.sv:56548:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_15_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_15_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_15_we),
		.wd(gpio_en_gpio_en_15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_15_ext_d_0),
		.qe(),
		.q(reg2hw[559]),
		.qs(gpio_en_gpio_en_15_qs)
	);
	// Trace: design.sv:56574:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_16_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_16_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_16_we),
		.wd(gpio_en_gpio_en_16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_16_ext_d_0),
		.qe(),
		.q(reg2hw[560]),
		.qs(gpio_en_gpio_en_16_qs)
	);
	// Trace: design.sv:56600:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_17_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_17_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_17_we),
		.wd(gpio_en_gpio_en_17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_17_ext_d_0),
		.qe(),
		.q(reg2hw[561]),
		.qs(gpio_en_gpio_en_17_qs)
	);
	// Trace: design.sv:56626:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_18_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_18_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_18_we),
		.wd(gpio_en_gpio_en_18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_18_ext_d_0),
		.qe(),
		.q(reg2hw[562]),
		.qs(gpio_en_gpio_en_18_qs)
	);
	// Trace: design.sv:56652:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_19_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_19_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_19_we),
		.wd(gpio_en_gpio_en_19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_19_ext_d_0),
		.qe(),
		.q(reg2hw[563]),
		.qs(gpio_en_gpio_en_19_qs)
	);
	// Trace: design.sv:56678:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_20_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_20_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_20_we),
		.wd(gpio_en_gpio_en_20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_20_ext_d_0),
		.qe(),
		.q(reg2hw[564]),
		.qs(gpio_en_gpio_en_20_qs)
	);
	// Trace: design.sv:56704:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_21_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_21_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_21_we),
		.wd(gpio_en_gpio_en_21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_21_ext_d_0),
		.qe(),
		.q(reg2hw[565]),
		.qs(gpio_en_gpio_en_21_qs)
	);
	// Trace: design.sv:56730:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_22_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_22_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_22_we),
		.wd(gpio_en_gpio_en_22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_22_ext_d_0),
		.qe(),
		.q(reg2hw[566]),
		.qs(gpio_en_gpio_en_22_qs)
	);
	// Trace: design.sv:56756:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_23_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_23_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_23_we),
		.wd(gpio_en_gpio_en_23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_23_ext_d_0),
		.qe(),
		.q(reg2hw[567]),
		.qs(gpio_en_gpio_en_23_qs)
	);
	// Trace: design.sv:56782:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_24_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_24_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_24_we),
		.wd(gpio_en_gpio_en_24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_24_ext_d_0),
		.qe(),
		.q(reg2hw[568]),
		.qs(gpio_en_gpio_en_24_qs)
	);
	// Trace: design.sv:56808:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_25_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_25_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_25_we),
		.wd(gpio_en_gpio_en_25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_25_ext_d_0),
		.qe(),
		.q(reg2hw[569]),
		.qs(gpio_en_gpio_en_25_qs)
	);
	// Trace: design.sv:56834:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_26_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_26_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_26_we),
		.wd(gpio_en_gpio_en_26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_26_ext_d_0),
		.qe(),
		.q(reg2hw[570]),
		.qs(gpio_en_gpio_en_26_qs)
	);
	// Trace: design.sv:56860:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_27_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_27_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_27_we),
		.wd(gpio_en_gpio_en_27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_27_ext_d_0),
		.qe(),
		.q(reg2hw[571]),
		.qs(gpio_en_gpio_en_27_qs)
	);
	// Trace: design.sv:56886:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_28_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_28_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_28_we),
		.wd(gpio_en_gpio_en_28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_28_ext_d_0),
		.qe(),
		.q(reg2hw[572]),
		.qs(gpio_en_gpio_en_28_qs)
	);
	// Trace: design.sv:56912:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_29_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_29_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_29_we),
		.wd(gpio_en_gpio_en_29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_29_ext_d_0),
		.qe(),
		.q(reg2hw[573]),
		.qs(gpio_en_gpio_en_29_qs)
	);
	// Trace: design.sv:56938:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_30_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_30_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_30_we),
		.wd(gpio_en_gpio_en_30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_30_ext_d_0),
		.qe(),
		.q(reg2hw[574]),
		.qs(gpio_en_gpio_en_30_qs)
	);
	// Trace: design.sv:56964:3
	localparam signed [31:0] sv2v_uu_u_gpio_en_gpio_en_31_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_en_gpio_en_31_d
	localparam [0:0] sv2v_uu_u_gpio_en_gpio_en_31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_en_gpio_en_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_en_gpio_en_31_we),
		.wd(gpio_en_gpio_en_31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_gpio_en_gpio_en_31_ext_d_0),
		.qe(),
		.q(reg2hw[575]),
		.qs(gpio_en_gpio_en_31_qs)
	);
	// Trace: design.sv:56995:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_0_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_0_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_0_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_0(
		.re(gpio_in_gpio_in_0_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_0_ext_wd_0),
		.d(hw2reg[352]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_0_qs)
	);
	// Trace: design.sv:57010:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_1_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_1_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_1_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_1(
		.re(gpio_in_gpio_in_1_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_1_ext_wd_0),
		.d(hw2reg[353]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_1_qs)
	);
	// Trace: design.sv:57025:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_2_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_2_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_2_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_2(
		.re(gpio_in_gpio_in_2_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_2_ext_wd_0),
		.d(hw2reg[354]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_2_qs)
	);
	// Trace: design.sv:57040:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_3_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_3_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_3_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_3(
		.re(gpio_in_gpio_in_3_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_3_ext_wd_0),
		.d(hw2reg[355]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_3_qs)
	);
	// Trace: design.sv:57055:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_4_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_4_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_4_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_4(
		.re(gpio_in_gpio_in_4_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_4_ext_wd_0),
		.d(hw2reg[356]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_4_qs)
	);
	// Trace: design.sv:57070:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_5_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_5_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_5_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_5(
		.re(gpio_in_gpio_in_5_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_5_ext_wd_0),
		.d(hw2reg[357]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_5_qs)
	);
	// Trace: design.sv:57085:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_6_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_6_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_6_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_6(
		.re(gpio_in_gpio_in_6_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_6_ext_wd_0),
		.d(hw2reg[358]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_6_qs)
	);
	// Trace: design.sv:57100:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_7_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_7_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_7_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_7(
		.re(gpio_in_gpio_in_7_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_7_ext_wd_0),
		.d(hw2reg[359]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_7_qs)
	);
	// Trace: design.sv:57115:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_8_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_8_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_8_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_8(
		.re(gpio_in_gpio_in_8_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_8_ext_wd_0),
		.d(hw2reg[360]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_8_qs)
	);
	// Trace: design.sv:57130:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_9_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_9_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_9_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_9(
		.re(gpio_in_gpio_in_9_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_9_ext_wd_0),
		.d(hw2reg[361]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_9_qs)
	);
	// Trace: design.sv:57145:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_10_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_10_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_10_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_10(
		.re(gpio_in_gpio_in_10_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_10_ext_wd_0),
		.d(hw2reg[362]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_10_qs)
	);
	// Trace: design.sv:57160:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_11_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_11_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_11_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_11(
		.re(gpio_in_gpio_in_11_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_11_ext_wd_0),
		.d(hw2reg[363]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_11_qs)
	);
	// Trace: design.sv:57175:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_12_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_12_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_12_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_12(
		.re(gpio_in_gpio_in_12_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_12_ext_wd_0),
		.d(hw2reg[364]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_12_qs)
	);
	// Trace: design.sv:57190:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_13_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_13_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_13_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_13(
		.re(gpio_in_gpio_in_13_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_13_ext_wd_0),
		.d(hw2reg[365]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_13_qs)
	);
	// Trace: design.sv:57205:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_14_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_14_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_14_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_14(
		.re(gpio_in_gpio_in_14_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_14_ext_wd_0),
		.d(hw2reg[366]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_14_qs)
	);
	// Trace: design.sv:57220:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_15_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_15_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_15_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_15(
		.re(gpio_in_gpio_in_15_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_15_ext_wd_0),
		.d(hw2reg[367]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_15_qs)
	);
	// Trace: design.sv:57235:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_16_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_16_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_16_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_16(
		.re(gpio_in_gpio_in_16_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_16_ext_wd_0),
		.d(hw2reg[368]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_16_qs)
	);
	// Trace: design.sv:57250:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_17_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_17_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_17_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_17(
		.re(gpio_in_gpio_in_17_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_17_ext_wd_0),
		.d(hw2reg[369]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_17_qs)
	);
	// Trace: design.sv:57265:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_18_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_18_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_18_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_18(
		.re(gpio_in_gpio_in_18_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_18_ext_wd_0),
		.d(hw2reg[370]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_18_qs)
	);
	// Trace: design.sv:57280:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_19_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_19_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_19_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_19(
		.re(gpio_in_gpio_in_19_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_19_ext_wd_0),
		.d(hw2reg[371]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_19_qs)
	);
	// Trace: design.sv:57295:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_20_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_20_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_20_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_20(
		.re(gpio_in_gpio_in_20_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_20_ext_wd_0),
		.d(hw2reg[372]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_20_qs)
	);
	// Trace: design.sv:57310:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_21_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_21_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_21_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_21(
		.re(gpio_in_gpio_in_21_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_21_ext_wd_0),
		.d(hw2reg[373]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_21_qs)
	);
	// Trace: design.sv:57325:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_22_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_22_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_22_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_22(
		.re(gpio_in_gpio_in_22_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_22_ext_wd_0),
		.d(hw2reg[374]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_22_qs)
	);
	// Trace: design.sv:57340:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_23_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_23_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_23_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_23(
		.re(gpio_in_gpio_in_23_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_23_ext_wd_0),
		.d(hw2reg[375]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_23_qs)
	);
	// Trace: design.sv:57355:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_24_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_24_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_24_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_24(
		.re(gpio_in_gpio_in_24_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_24_ext_wd_0),
		.d(hw2reg[376]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_24_qs)
	);
	// Trace: design.sv:57370:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_25_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_25_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_25_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_25(
		.re(gpio_in_gpio_in_25_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_25_ext_wd_0),
		.d(hw2reg[377]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_25_qs)
	);
	// Trace: design.sv:57385:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_26_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_26_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_26_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_26(
		.re(gpio_in_gpio_in_26_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_26_ext_wd_0),
		.d(hw2reg[378]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_26_qs)
	);
	// Trace: design.sv:57400:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_27_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_27_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_27_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_27(
		.re(gpio_in_gpio_in_27_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_27_ext_wd_0),
		.d(hw2reg[379]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_27_qs)
	);
	// Trace: design.sv:57415:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_28_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_28_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_28_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_28(
		.re(gpio_in_gpio_in_28_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_28_ext_wd_0),
		.d(hw2reg[380]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_28_qs)
	);
	// Trace: design.sv:57430:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_29_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_29_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_29_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_29(
		.re(gpio_in_gpio_in_29_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_29_ext_wd_0),
		.d(hw2reg[381]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_29_qs)
	);
	// Trace: design.sv:57445:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_30_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_30_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_30_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_30(
		.re(gpio_in_gpio_in_30_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_30_ext_wd_0),
		.d(hw2reg[382]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_30_qs)
	);
	// Trace: design.sv:57460:3
	localparam [31:0] sv2v_uu_u_gpio_in_gpio_in_31_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_in_gpio_in_31_wd
	localparam [0:0] sv2v_uu_u_gpio_in_gpio_in_31_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_in_gpio_in_31(
		.re(gpio_in_gpio_in_31_re),
		.we(1'b0),
		.wd(sv2v_uu_u_gpio_in_gpio_in_31_ext_wd_0),
		.d(hw2reg[383]),
		.qre(),
		.qe(),
		.q(),
		.qs(gpio_in_gpio_in_31_qs)
	);
	// Trace: design.sv:57480:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_0_we),
		.wd(gpio_out_gpio_out_0_wd),
		.de(hw2reg[288]),
		.d(hw2reg[289]),
		.qe(),
		.q(reg2hw[512]),
		.qs(gpio_out_gpio_out_0_qs)
	);
	// Trace: design.sv:57506:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_1_we),
		.wd(gpio_out_gpio_out_1_wd),
		.de(hw2reg[290]),
		.d(hw2reg[291]),
		.qe(),
		.q(reg2hw[513]),
		.qs(gpio_out_gpio_out_1_qs)
	);
	// Trace: design.sv:57532:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_2_we),
		.wd(gpio_out_gpio_out_2_wd),
		.de(hw2reg[292]),
		.d(hw2reg[293]),
		.qe(),
		.q(reg2hw[514]),
		.qs(gpio_out_gpio_out_2_qs)
	);
	// Trace: design.sv:57558:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_3_we),
		.wd(gpio_out_gpio_out_3_wd),
		.de(hw2reg[294]),
		.d(hw2reg[295]),
		.qe(),
		.q(reg2hw[515]),
		.qs(gpio_out_gpio_out_3_qs)
	);
	// Trace: design.sv:57584:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_4_we),
		.wd(gpio_out_gpio_out_4_wd),
		.de(hw2reg[296]),
		.d(hw2reg[297]),
		.qe(),
		.q(reg2hw[516]),
		.qs(gpio_out_gpio_out_4_qs)
	);
	// Trace: design.sv:57610:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_5_we),
		.wd(gpio_out_gpio_out_5_wd),
		.de(hw2reg[298]),
		.d(hw2reg[299]),
		.qe(),
		.q(reg2hw[517]),
		.qs(gpio_out_gpio_out_5_qs)
	);
	// Trace: design.sv:57636:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_6_we),
		.wd(gpio_out_gpio_out_6_wd),
		.de(hw2reg[300]),
		.d(hw2reg[301]),
		.qe(),
		.q(reg2hw[518]),
		.qs(gpio_out_gpio_out_6_qs)
	);
	// Trace: design.sv:57662:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_7_we),
		.wd(gpio_out_gpio_out_7_wd),
		.de(hw2reg[302]),
		.d(hw2reg[303]),
		.qe(),
		.q(reg2hw[519]),
		.qs(gpio_out_gpio_out_7_qs)
	);
	// Trace: design.sv:57688:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_8_we),
		.wd(gpio_out_gpio_out_8_wd),
		.de(hw2reg[304]),
		.d(hw2reg[305]),
		.qe(),
		.q(reg2hw[520]),
		.qs(gpio_out_gpio_out_8_qs)
	);
	// Trace: design.sv:57714:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_9_we),
		.wd(gpio_out_gpio_out_9_wd),
		.de(hw2reg[306]),
		.d(hw2reg[307]),
		.qe(),
		.q(reg2hw[521]),
		.qs(gpio_out_gpio_out_9_qs)
	);
	// Trace: design.sv:57740:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_10_we),
		.wd(gpio_out_gpio_out_10_wd),
		.de(hw2reg[308]),
		.d(hw2reg[309]),
		.qe(),
		.q(reg2hw[522]),
		.qs(gpio_out_gpio_out_10_qs)
	);
	// Trace: design.sv:57766:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_11_we),
		.wd(gpio_out_gpio_out_11_wd),
		.de(hw2reg[310]),
		.d(hw2reg[311]),
		.qe(),
		.q(reg2hw[523]),
		.qs(gpio_out_gpio_out_11_qs)
	);
	// Trace: design.sv:57792:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_12_we),
		.wd(gpio_out_gpio_out_12_wd),
		.de(hw2reg[312]),
		.d(hw2reg[313]),
		.qe(),
		.q(reg2hw[524]),
		.qs(gpio_out_gpio_out_12_qs)
	);
	// Trace: design.sv:57818:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_13_we),
		.wd(gpio_out_gpio_out_13_wd),
		.de(hw2reg[314]),
		.d(hw2reg[315]),
		.qe(),
		.q(reg2hw[525]),
		.qs(gpio_out_gpio_out_13_qs)
	);
	// Trace: design.sv:57844:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_14_we),
		.wd(gpio_out_gpio_out_14_wd),
		.de(hw2reg[316]),
		.d(hw2reg[317]),
		.qe(),
		.q(reg2hw[526]),
		.qs(gpio_out_gpio_out_14_qs)
	);
	// Trace: design.sv:57870:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_15_we),
		.wd(gpio_out_gpio_out_15_wd),
		.de(hw2reg[318]),
		.d(hw2reg[319]),
		.qe(),
		.q(reg2hw[527]),
		.qs(gpio_out_gpio_out_15_qs)
	);
	// Trace: design.sv:57896:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_16_we),
		.wd(gpio_out_gpio_out_16_wd),
		.de(hw2reg[320]),
		.d(hw2reg[321]),
		.qe(),
		.q(reg2hw[528]),
		.qs(gpio_out_gpio_out_16_qs)
	);
	// Trace: design.sv:57922:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_17_we),
		.wd(gpio_out_gpio_out_17_wd),
		.de(hw2reg[322]),
		.d(hw2reg[323]),
		.qe(),
		.q(reg2hw[529]),
		.qs(gpio_out_gpio_out_17_qs)
	);
	// Trace: design.sv:57948:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_18_we),
		.wd(gpio_out_gpio_out_18_wd),
		.de(hw2reg[324]),
		.d(hw2reg[325]),
		.qe(),
		.q(reg2hw[530]),
		.qs(gpio_out_gpio_out_18_qs)
	);
	// Trace: design.sv:57974:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_19_we),
		.wd(gpio_out_gpio_out_19_wd),
		.de(hw2reg[326]),
		.d(hw2reg[327]),
		.qe(),
		.q(reg2hw[531]),
		.qs(gpio_out_gpio_out_19_qs)
	);
	// Trace: design.sv:58000:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_20_we),
		.wd(gpio_out_gpio_out_20_wd),
		.de(hw2reg[328]),
		.d(hw2reg[329]),
		.qe(),
		.q(reg2hw[532]),
		.qs(gpio_out_gpio_out_20_qs)
	);
	// Trace: design.sv:58026:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_21_we),
		.wd(gpio_out_gpio_out_21_wd),
		.de(hw2reg[330]),
		.d(hw2reg[331]),
		.qe(),
		.q(reg2hw[533]),
		.qs(gpio_out_gpio_out_21_qs)
	);
	// Trace: design.sv:58052:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_22_we),
		.wd(gpio_out_gpio_out_22_wd),
		.de(hw2reg[332]),
		.d(hw2reg[333]),
		.qe(),
		.q(reg2hw[534]),
		.qs(gpio_out_gpio_out_22_qs)
	);
	// Trace: design.sv:58078:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_23_we),
		.wd(gpio_out_gpio_out_23_wd),
		.de(hw2reg[334]),
		.d(hw2reg[335]),
		.qe(),
		.q(reg2hw[535]),
		.qs(gpio_out_gpio_out_23_qs)
	);
	// Trace: design.sv:58104:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_24_we),
		.wd(gpio_out_gpio_out_24_wd),
		.de(hw2reg[336]),
		.d(hw2reg[337]),
		.qe(),
		.q(reg2hw[536]),
		.qs(gpio_out_gpio_out_24_qs)
	);
	// Trace: design.sv:58130:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_25_we),
		.wd(gpio_out_gpio_out_25_wd),
		.de(hw2reg[338]),
		.d(hw2reg[339]),
		.qe(),
		.q(reg2hw[537]),
		.qs(gpio_out_gpio_out_25_qs)
	);
	// Trace: design.sv:58156:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_26_we),
		.wd(gpio_out_gpio_out_26_wd),
		.de(hw2reg[340]),
		.d(hw2reg[341]),
		.qe(),
		.q(reg2hw[538]),
		.qs(gpio_out_gpio_out_26_qs)
	);
	// Trace: design.sv:58182:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_27_we),
		.wd(gpio_out_gpio_out_27_wd),
		.de(hw2reg[342]),
		.d(hw2reg[343]),
		.qe(),
		.q(reg2hw[539]),
		.qs(gpio_out_gpio_out_27_qs)
	);
	// Trace: design.sv:58208:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_28_we),
		.wd(gpio_out_gpio_out_28_wd),
		.de(hw2reg[344]),
		.d(hw2reg[345]),
		.qe(),
		.q(reg2hw[540]),
		.qs(gpio_out_gpio_out_28_qs)
	);
	// Trace: design.sv:58234:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_29_we),
		.wd(gpio_out_gpio_out_29_wd),
		.de(hw2reg[346]),
		.d(hw2reg[347]),
		.qe(),
		.q(reg2hw[541]),
		.qs(gpio_out_gpio_out_29_qs)
	);
	// Trace: design.sv:58260:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_30_we),
		.wd(gpio_out_gpio_out_30_wd),
		.de(hw2reg[348]),
		.d(hw2reg[349]),
		.qe(),
		.q(reg2hw[542]),
		.qs(gpio_out_gpio_out_30_qs)
	);
	// Trace: design.sv:58286:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_gpio_out_gpio_out_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(gpio_out_gpio_out_31_we),
		.wd(gpio_out_gpio_out_31_wd),
		.de(hw2reg[350]),
		.d(hw2reg[351]),
		.qe(),
		.q(reg2hw[543]),
		.qs(gpio_out_gpio_out_31_qs)
	);
	// Trace: design.sv:58317:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_0_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_0_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_0_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_0(
		.re(1'b0),
		.we(gpio_set_gpio_set_0_we),
		.wd(gpio_set_gpio_set_0_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_0_ext_d_0),
		.qre(),
		.qe(reg2hw[448]),
		.q(reg2hw[449]),
		.qs()
	);
	// Trace: design.sv:58332:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_1_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_1_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_1_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_1(
		.re(1'b0),
		.we(gpio_set_gpio_set_1_we),
		.wd(gpio_set_gpio_set_1_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_1_ext_d_0),
		.qre(),
		.qe(reg2hw[450]),
		.q(reg2hw[451]),
		.qs()
	);
	// Trace: design.sv:58347:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_2_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_2_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_2_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_2(
		.re(1'b0),
		.we(gpio_set_gpio_set_2_we),
		.wd(gpio_set_gpio_set_2_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_2_ext_d_0),
		.qre(),
		.qe(reg2hw[452]),
		.q(reg2hw[453]),
		.qs()
	);
	// Trace: design.sv:58362:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_3_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_3_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_3_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_3(
		.re(1'b0),
		.we(gpio_set_gpio_set_3_we),
		.wd(gpio_set_gpio_set_3_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_3_ext_d_0),
		.qre(),
		.qe(reg2hw[454]),
		.q(reg2hw[455]),
		.qs()
	);
	// Trace: design.sv:58377:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_4_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_4_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_4_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_4(
		.re(1'b0),
		.we(gpio_set_gpio_set_4_we),
		.wd(gpio_set_gpio_set_4_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_4_ext_d_0),
		.qre(),
		.qe(reg2hw[456]),
		.q(reg2hw[457]),
		.qs()
	);
	// Trace: design.sv:58392:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_5_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_5_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_5_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_5(
		.re(1'b0),
		.we(gpio_set_gpio_set_5_we),
		.wd(gpio_set_gpio_set_5_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_5_ext_d_0),
		.qre(),
		.qe(reg2hw[458]),
		.q(reg2hw[459]),
		.qs()
	);
	// Trace: design.sv:58407:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_6_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_6_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_6_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_6(
		.re(1'b0),
		.we(gpio_set_gpio_set_6_we),
		.wd(gpio_set_gpio_set_6_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_6_ext_d_0),
		.qre(),
		.qe(reg2hw[460]),
		.q(reg2hw[461]),
		.qs()
	);
	// Trace: design.sv:58422:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_7_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_7_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_7_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_7(
		.re(1'b0),
		.we(gpio_set_gpio_set_7_we),
		.wd(gpio_set_gpio_set_7_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_7_ext_d_0),
		.qre(),
		.qe(reg2hw[462]),
		.q(reg2hw[463]),
		.qs()
	);
	// Trace: design.sv:58437:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_8_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_8_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_8_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_8(
		.re(1'b0),
		.we(gpio_set_gpio_set_8_we),
		.wd(gpio_set_gpio_set_8_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_8_ext_d_0),
		.qre(),
		.qe(reg2hw[464]),
		.q(reg2hw[465]),
		.qs()
	);
	// Trace: design.sv:58452:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_9_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_9_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_9_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_9(
		.re(1'b0),
		.we(gpio_set_gpio_set_9_we),
		.wd(gpio_set_gpio_set_9_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_9_ext_d_0),
		.qre(),
		.qe(reg2hw[466]),
		.q(reg2hw[467]),
		.qs()
	);
	// Trace: design.sv:58467:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_10_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_10_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_10_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_10(
		.re(1'b0),
		.we(gpio_set_gpio_set_10_we),
		.wd(gpio_set_gpio_set_10_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_10_ext_d_0),
		.qre(),
		.qe(reg2hw[468]),
		.q(reg2hw[469]),
		.qs()
	);
	// Trace: design.sv:58482:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_11_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_11_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_11_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_11(
		.re(1'b0),
		.we(gpio_set_gpio_set_11_we),
		.wd(gpio_set_gpio_set_11_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_11_ext_d_0),
		.qre(),
		.qe(reg2hw[470]),
		.q(reg2hw[471]),
		.qs()
	);
	// Trace: design.sv:58497:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_12_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_12_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_12_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_12(
		.re(1'b0),
		.we(gpio_set_gpio_set_12_we),
		.wd(gpio_set_gpio_set_12_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_12_ext_d_0),
		.qre(),
		.qe(reg2hw[472]),
		.q(reg2hw[473]),
		.qs()
	);
	// Trace: design.sv:58512:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_13_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_13_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_13_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_13(
		.re(1'b0),
		.we(gpio_set_gpio_set_13_we),
		.wd(gpio_set_gpio_set_13_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_13_ext_d_0),
		.qre(),
		.qe(reg2hw[474]),
		.q(reg2hw[475]),
		.qs()
	);
	// Trace: design.sv:58527:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_14_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_14_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_14_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_14(
		.re(1'b0),
		.we(gpio_set_gpio_set_14_we),
		.wd(gpio_set_gpio_set_14_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_14_ext_d_0),
		.qre(),
		.qe(reg2hw[476]),
		.q(reg2hw[477]),
		.qs()
	);
	// Trace: design.sv:58542:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_15_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_15_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_15_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_15(
		.re(1'b0),
		.we(gpio_set_gpio_set_15_we),
		.wd(gpio_set_gpio_set_15_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_15_ext_d_0),
		.qre(),
		.qe(reg2hw[478]),
		.q(reg2hw[479]),
		.qs()
	);
	// Trace: design.sv:58557:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_16_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_16_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_16_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_16(
		.re(1'b0),
		.we(gpio_set_gpio_set_16_we),
		.wd(gpio_set_gpio_set_16_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_16_ext_d_0),
		.qre(),
		.qe(reg2hw[480]),
		.q(reg2hw[481]),
		.qs()
	);
	// Trace: design.sv:58572:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_17_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_17_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_17_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_17(
		.re(1'b0),
		.we(gpio_set_gpio_set_17_we),
		.wd(gpio_set_gpio_set_17_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_17_ext_d_0),
		.qre(),
		.qe(reg2hw[482]),
		.q(reg2hw[483]),
		.qs()
	);
	// Trace: design.sv:58587:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_18_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_18_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_18_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_18(
		.re(1'b0),
		.we(gpio_set_gpio_set_18_we),
		.wd(gpio_set_gpio_set_18_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_18_ext_d_0),
		.qre(),
		.qe(reg2hw[484]),
		.q(reg2hw[485]),
		.qs()
	);
	// Trace: design.sv:58602:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_19_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_19_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_19_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_19(
		.re(1'b0),
		.we(gpio_set_gpio_set_19_we),
		.wd(gpio_set_gpio_set_19_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_19_ext_d_0),
		.qre(),
		.qe(reg2hw[486]),
		.q(reg2hw[487]),
		.qs()
	);
	// Trace: design.sv:58617:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_20_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_20_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_20_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_20(
		.re(1'b0),
		.we(gpio_set_gpio_set_20_we),
		.wd(gpio_set_gpio_set_20_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_20_ext_d_0),
		.qre(),
		.qe(reg2hw[488]),
		.q(reg2hw[489]),
		.qs()
	);
	// Trace: design.sv:58632:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_21_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_21_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_21_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_21(
		.re(1'b0),
		.we(gpio_set_gpio_set_21_we),
		.wd(gpio_set_gpio_set_21_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_21_ext_d_0),
		.qre(),
		.qe(reg2hw[490]),
		.q(reg2hw[491]),
		.qs()
	);
	// Trace: design.sv:58647:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_22_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_22_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_22_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_22(
		.re(1'b0),
		.we(gpio_set_gpio_set_22_we),
		.wd(gpio_set_gpio_set_22_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_22_ext_d_0),
		.qre(),
		.qe(reg2hw[492]),
		.q(reg2hw[493]),
		.qs()
	);
	// Trace: design.sv:58662:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_23_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_23_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_23_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_23(
		.re(1'b0),
		.we(gpio_set_gpio_set_23_we),
		.wd(gpio_set_gpio_set_23_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_23_ext_d_0),
		.qre(),
		.qe(reg2hw[494]),
		.q(reg2hw[495]),
		.qs()
	);
	// Trace: design.sv:58677:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_24_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_24_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_24_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_24(
		.re(1'b0),
		.we(gpio_set_gpio_set_24_we),
		.wd(gpio_set_gpio_set_24_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_24_ext_d_0),
		.qre(),
		.qe(reg2hw[496]),
		.q(reg2hw[497]),
		.qs()
	);
	// Trace: design.sv:58692:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_25_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_25_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_25_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_25(
		.re(1'b0),
		.we(gpio_set_gpio_set_25_we),
		.wd(gpio_set_gpio_set_25_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_25_ext_d_0),
		.qre(),
		.qe(reg2hw[498]),
		.q(reg2hw[499]),
		.qs()
	);
	// Trace: design.sv:58707:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_26_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_26_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_26_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_26(
		.re(1'b0),
		.we(gpio_set_gpio_set_26_we),
		.wd(gpio_set_gpio_set_26_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_26_ext_d_0),
		.qre(),
		.qe(reg2hw[500]),
		.q(reg2hw[501]),
		.qs()
	);
	// Trace: design.sv:58722:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_27_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_27_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_27_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_27(
		.re(1'b0),
		.we(gpio_set_gpio_set_27_we),
		.wd(gpio_set_gpio_set_27_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_27_ext_d_0),
		.qre(),
		.qe(reg2hw[502]),
		.q(reg2hw[503]),
		.qs()
	);
	// Trace: design.sv:58737:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_28_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_28_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_28_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_28(
		.re(1'b0),
		.we(gpio_set_gpio_set_28_we),
		.wd(gpio_set_gpio_set_28_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_28_ext_d_0),
		.qre(),
		.qe(reg2hw[504]),
		.q(reg2hw[505]),
		.qs()
	);
	// Trace: design.sv:58752:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_29_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_29_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_29_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_29(
		.re(1'b0),
		.we(gpio_set_gpio_set_29_we),
		.wd(gpio_set_gpio_set_29_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_29_ext_d_0),
		.qre(),
		.qe(reg2hw[506]),
		.q(reg2hw[507]),
		.qs()
	);
	// Trace: design.sv:58767:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_30_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_30_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_30_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_30(
		.re(1'b0),
		.we(gpio_set_gpio_set_30_we),
		.wd(gpio_set_gpio_set_30_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_30_ext_d_0),
		.qre(),
		.qe(reg2hw[508]),
		.q(reg2hw[509]),
		.qs()
	);
	// Trace: design.sv:58782:3
	localparam [31:0] sv2v_uu_u_gpio_set_gpio_set_31_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_set_gpio_set_31_d
	localparam [0:0] sv2v_uu_u_gpio_set_gpio_set_31_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_set_gpio_set_31(
		.re(1'b0),
		.we(gpio_set_gpio_set_31_we),
		.wd(gpio_set_gpio_set_31_wd),
		.d(sv2v_uu_u_gpio_set_gpio_set_31_ext_d_0),
		.qre(),
		.qe(reg2hw[510]),
		.q(reg2hw[511]),
		.qs()
	);
	// Trace: design.sv:58802:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_0_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_0_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_0_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_0(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_0_we),
		.wd(gpio_clear_gpio_clear_0_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_0_ext_d_0),
		.qre(),
		.qe(reg2hw[384]),
		.q(reg2hw[385]),
		.qs()
	);
	// Trace: design.sv:58817:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_1_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_1_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_1_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_1(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_1_we),
		.wd(gpio_clear_gpio_clear_1_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_1_ext_d_0),
		.qre(),
		.qe(reg2hw[386]),
		.q(reg2hw[387]),
		.qs()
	);
	// Trace: design.sv:58832:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_2_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_2_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_2_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_2(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_2_we),
		.wd(gpio_clear_gpio_clear_2_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_2_ext_d_0),
		.qre(),
		.qe(reg2hw[388]),
		.q(reg2hw[389]),
		.qs()
	);
	// Trace: design.sv:58847:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_3_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_3_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_3_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_3(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_3_we),
		.wd(gpio_clear_gpio_clear_3_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_3_ext_d_0),
		.qre(),
		.qe(reg2hw[390]),
		.q(reg2hw[391]),
		.qs()
	);
	// Trace: design.sv:58862:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_4_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_4_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_4_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_4(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_4_we),
		.wd(gpio_clear_gpio_clear_4_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_4_ext_d_0),
		.qre(),
		.qe(reg2hw[392]),
		.q(reg2hw[393]),
		.qs()
	);
	// Trace: design.sv:58877:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_5_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_5_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_5_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_5(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_5_we),
		.wd(gpio_clear_gpio_clear_5_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_5_ext_d_0),
		.qre(),
		.qe(reg2hw[394]),
		.q(reg2hw[395]),
		.qs()
	);
	// Trace: design.sv:58892:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_6_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_6_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_6_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_6(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_6_we),
		.wd(gpio_clear_gpio_clear_6_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_6_ext_d_0),
		.qre(),
		.qe(reg2hw[396]),
		.q(reg2hw[397]),
		.qs()
	);
	// Trace: design.sv:58907:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_7_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_7_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_7_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_7(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_7_we),
		.wd(gpio_clear_gpio_clear_7_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_7_ext_d_0),
		.qre(),
		.qe(reg2hw[398]),
		.q(reg2hw[399]),
		.qs()
	);
	// Trace: design.sv:58922:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_8_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_8_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_8_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_8(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_8_we),
		.wd(gpio_clear_gpio_clear_8_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_8_ext_d_0),
		.qre(),
		.qe(reg2hw[400]),
		.q(reg2hw[401]),
		.qs()
	);
	// Trace: design.sv:58937:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_9_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_9_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_9_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_9(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_9_we),
		.wd(gpio_clear_gpio_clear_9_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_9_ext_d_0),
		.qre(),
		.qe(reg2hw[402]),
		.q(reg2hw[403]),
		.qs()
	);
	// Trace: design.sv:58952:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_10_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_10_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_10_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_10(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_10_we),
		.wd(gpio_clear_gpio_clear_10_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_10_ext_d_0),
		.qre(),
		.qe(reg2hw[404]),
		.q(reg2hw[405]),
		.qs()
	);
	// Trace: design.sv:58967:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_11_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_11_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_11_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_11(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_11_we),
		.wd(gpio_clear_gpio_clear_11_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_11_ext_d_0),
		.qre(),
		.qe(reg2hw[406]),
		.q(reg2hw[407]),
		.qs()
	);
	// Trace: design.sv:58982:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_12_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_12_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_12_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_12(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_12_we),
		.wd(gpio_clear_gpio_clear_12_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_12_ext_d_0),
		.qre(),
		.qe(reg2hw[408]),
		.q(reg2hw[409]),
		.qs()
	);
	// Trace: design.sv:58997:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_13_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_13_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_13_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_13(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_13_we),
		.wd(gpio_clear_gpio_clear_13_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_13_ext_d_0),
		.qre(),
		.qe(reg2hw[410]),
		.q(reg2hw[411]),
		.qs()
	);
	// Trace: design.sv:59012:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_14_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_14_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_14_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_14(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_14_we),
		.wd(gpio_clear_gpio_clear_14_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_14_ext_d_0),
		.qre(),
		.qe(reg2hw[412]),
		.q(reg2hw[413]),
		.qs()
	);
	// Trace: design.sv:59027:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_15_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_15_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_15_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_15(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_15_we),
		.wd(gpio_clear_gpio_clear_15_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_15_ext_d_0),
		.qre(),
		.qe(reg2hw[414]),
		.q(reg2hw[415]),
		.qs()
	);
	// Trace: design.sv:59042:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_16_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_16_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_16_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_16(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_16_we),
		.wd(gpio_clear_gpio_clear_16_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_16_ext_d_0),
		.qre(),
		.qe(reg2hw[416]),
		.q(reg2hw[417]),
		.qs()
	);
	// Trace: design.sv:59057:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_17_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_17_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_17_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_17(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_17_we),
		.wd(gpio_clear_gpio_clear_17_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_17_ext_d_0),
		.qre(),
		.qe(reg2hw[418]),
		.q(reg2hw[419]),
		.qs()
	);
	// Trace: design.sv:59072:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_18_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_18_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_18_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_18(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_18_we),
		.wd(gpio_clear_gpio_clear_18_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_18_ext_d_0),
		.qre(),
		.qe(reg2hw[420]),
		.q(reg2hw[421]),
		.qs()
	);
	// Trace: design.sv:59087:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_19_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_19_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_19_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_19(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_19_we),
		.wd(gpio_clear_gpio_clear_19_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_19_ext_d_0),
		.qre(),
		.qe(reg2hw[422]),
		.q(reg2hw[423]),
		.qs()
	);
	// Trace: design.sv:59102:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_20_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_20_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_20_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_20(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_20_we),
		.wd(gpio_clear_gpio_clear_20_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_20_ext_d_0),
		.qre(),
		.qe(reg2hw[424]),
		.q(reg2hw[425]),
		.qs()
	);
	// Trace: design.sv:59117:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_21_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_21_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_21_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_21(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_21_we),
		.wd(gpio_clear_gpio_clear_21_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_21_ext_d_0),
		.qre(),
		.qe(reg2hw[426]),
		.q(reg2hw[427]),
		.qs()
	);
	// Trace: design.sv:59132:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_22_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_22_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_22_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_22(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_22_we),
		.wd(gpio_clear_gpio_clear_22_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_22_ext_d_0),
		.qre(),
		.qe(reg2hw[428]),
		.q(reg2hw[429]),
		.qs()
	);
	// Trace: design.sv:59147:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_23_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_23_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_23_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_23(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_23_we),
		.wd(gpio_clear_gpio_clear_23_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_23_ext_d_0),
		.qre(),
		.qe(reg2hw[430]),
		.q(reg2hw[431]),
		.qs()
	);
	// Trace: design.sv:59162:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_24_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_24_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_24_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_24(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_24_we),
		.wd(gpio_clear_gpio_clear_24_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_24_ext_d_0),
		.qre(),
		.qe(reg2hw[432]),
		.q(reg2hw[433]),
		.qs()
	);
	// Trace: design.sv:59177:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_25_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_25_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_25_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_25(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_25_we),
		.wd(gpio_clear_gpio_clear_25_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_25_ext_d_0),
		.qre(),
		.qe(reg2hw[434]),
		.q(reg2hw[435]),
		.qs()
	);
	// Trace: design.sv:59192:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_26_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_26_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_26_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_26(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_26_we),
		.wd(gpio_clear_gpio_clear_26_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_26_ext_d_0),
		.qre(),
		.qe(reg2hw[436]),
		.q(reg2hw[437]),
		.qs()
	);
	// Trace: design.sv:59207:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_27_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_27_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_27_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_27(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_27_we),
		.wd(gpio_clear_gpio_clear_27_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_27_ext_d_0),
		.qre(),
		.qe(reg2hw[438]),
		.q(reg2hw[439]),
		.qs()
	);
	// Trace: design.sv:59222:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_28_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_28_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_28_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_28(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_28_we),
		.wd(gpio_clear_gpio_clear_28_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_28_ext_d_0),
		.qre(),
		.qe(reg2hw[440]),
		.q(reg2hw[441]),
		.qs()
	);
	// Trace: design.sv:59237:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_29_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_29_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_29_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_29(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_29_we),
		.wd(gpio_clear_gpio_clear_29_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_29_ext_d_0),
		.qre(),
		.qe(reg2hw[442]),
		.q(reg2hw[443]),
		.qs()
	);
	// Trace: design.sv:59252:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_30_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_30_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_30_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_30(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_30_we),
		.wd(gpio_clear_gpio_clear_30_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_30_ext_d_0),
		.qre(),
		.qe(reg2hw[444]),
		.q(reg2hw[445]),
		.qs()
	);
	// Trace: design.sv:59267:3
	localparam [31:0] sv2v_uu_u_gpio_clear_gpio_clear_31_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_clear_gpio_clear_31_d
	localparam [0:0] sv2v_uu_u_gpio_clear_gpio_clear_31_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_clear_gpio_clear_31(
		.re(1'b0),
		.we(gpio_clear_gpio_clear_31_we),
		.wd(gpio_clear_gpio_clear_31_wd),
		.d(sv2v_uu_u_gpio_clear_gpio_clear_31_ext_d_0),
		.qre(),
		.qe(reg2hw[446]),
		.q(reg2hw[447]),
		.qs()
	);
	// Trace: design.sv:59287:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_0_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_0_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_0_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_0(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_0_we),
		.wd(gpio_toggle_gpio_toggle_0_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_0_ext_d_0),
		.qre(),
		.qe(reg2hw[320]),
		.q(reg2hw[321]),
		.qs()
	);
	// Trace: design.sv:59302:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_1_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_1_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_1_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_1(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_1_we),
		.wd(gpio_toggle_gpio_toggle_1_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_1_ext_d_0),
		.qre(),
		.qe(reg2hw[322]),
		.q(reg2hw[323]),
		.qs()
	);
	// Trace: design.sv:59317:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_2_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_2_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_2_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_2(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_2_we),
		.wd(gpio_toggle_gpio_toggle_2_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_2_ext_d_0),
		.qre(),
		.qe(reg2hw[324]),
		.q(reg2hw[325]),
		.qs()
	);
	// Trace: design.sv:59332:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_3_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_3_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_3_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_3(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_3_we),
		.wd(gpio_toggle_gpio_toggle_3_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_3_ext_d_0),
		.qre(),
		.qe(reg2hw[326]),
		.q(reg2hw[327]),
		.qs()
	);
	// Trace: design.sv:59347:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_4_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_4_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_4_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_4(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_4_we),
		.wd(gpio_toggle_gpio_toggle_4_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_4_ext_d_0),
		.qre(),
		.qe(reg2hw[328]),
		.q(reg2hw[329]),
		.qs()
	);
	// Trace: design.sv:59362:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_5_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_5_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_5_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_5(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_5_we),
		.wd(gpio_toggle_gpio_toggle_5_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_5_ext_d_0),
		.qre(),
		.qe(reg2hw[330]),
		.q(reg2hw[331]),
		.qs()
	);
	// Trace: design.sv:59377:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_6_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_6_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_6_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_6(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_6_we),
		.wd(gpio_toggle_gpio_toggle_6_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_6_ext_d_0),
		.qre(),
		.qe(reg2hw[332]),
		.q(reg2hw[333]),
		.qs()
	);
	// Trace: design.sv:59392:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_7_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_7_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_7_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_7(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_7_we),
		.wd(gpio_toggle_gpio_toggle_7_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_7_ext_d_0),
		.qre(),
		.qe(reg2hw[334]),
		.q(reg2hw[335]),
		.qs()
	);
	// Trace: design.sv:59407:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_8_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_8_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_8_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_8(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_8_we),
		.wd(gpio_toggle_gpio_toggle_8_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_8_ext_d_0),
		.qre(),
		.qe(reg2hw[336]),
		.q(reg2hw[337]),
		.qs()
	);
	// Trace: design.sv:59422:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_9_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_9_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_9_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_9(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_9_we),
		.wd(gpio_toggle_gpio_toggle_9_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_9_ext_d_0),
		.qre(),
		.qe(reg2hw[338]),
		.q(reg2hw[339]),
		.qs()
	);
	// Trace: design.sv:59437:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_10_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_10_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_10_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_10(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_10_we),
		.wd(gpio_toggle_gpio_toggle_10_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_10_ext_d_0),
		.qre(),
		.qe(reg2hw[340]),
		.q(reg2hw[341]),
		.qs()
	);
	// Trace: design.sv:59452:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_11_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_11_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_11_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_11(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_11_we),
		.wd(gpio_toggle_gpio_toggle_11_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_11_ext_d_0),
		.qre(),
		.qe(reg2hw[342]),
		.q(reg2hw[343]),
		.qs()
	);
	// Trace: design.sv:59467:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_12_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_12_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_12_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_12(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_12_we),
		.wd(gpio_toggle_gpio_toggle_12_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_12_ext_d_0),
		.qre(),
		.qe(reg2hw[344]),
		.q(reg2hw[345]),
		.qs()
	);
	// Trace: design.sv:59482:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_13_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_13_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_13_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_13(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_13_we),
		.wd(gpio_toggle_gpio_toggle_13_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_13_ext_d_0),
		.qre(),
		.qe(reg2hw[346]),
		.q(reg2hw[347]),
		.qs()
	);
	// Trace: design.sv:59497:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_14_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_14_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_14_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_14(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_14_we),
		.wd(gpio_toggle_gpio_toggle_14_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_14_ext_d_0),
		.qre(),
		.qe(reg2hw[348]),
		.q(reg2hw[349]),
		.qs()
	);
	// Trace: design.sv:59512:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_15_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_15_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_15_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_15(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_15_we),
		.wd(gpio_toggle_gpio_toggle_15_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_15_ext_d_0),
		.qre(),
		.qe(reg2hw[350]),
		.q(reg2hw[351]),
		.qs()
	);
	// Trace: design.sv:59527:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_16_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_16_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_16_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_16(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_16_we),
		.wd(gpio_toggle_gpio_toggle_16_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_16_ext_d_0),
		.qre(),
		.qe(reg2hw[352]),
		.q(reg2hw[353]),
		.qs()
	);
	// Trace: design.sv:59542:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_17_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_17_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_17_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_17(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_17_we),
		.wd(gpio_toggle_gpio_toggle_17_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_17_ext_d_0),
		.qre(),
		.qe(reg2hw[354]),
		.q(reg2hw[355]),
		.qs()
	);
	// Trace: design.sv:59557:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_18_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_18_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_18_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_18(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_18_we),
		.wd(gpio_toggle_gpio_toggle_18_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_18_ext_d_0),
		.qre(),
		.qe(reg2hw[356]),
		.q(reg2hw[357]),
		.qs()
	);
	// Trace: design.sv:59572:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_19_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_19_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_19_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_19(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_19_we),
		.wd(gpio_toggle_gpio_toggle_19_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_19_ext_d_0),
		.qre(),
		.qe(reg2hw[358]),
		.q(reg2hw[359]),
		.qs()
	);
	// Trace: design.sv:59587:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_20_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_20_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_20_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_20(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_20_we),
		.wd(gpio_toggle_gpio_toggle_20_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_20_ext_d_0),
		.qre(),
		.qe(reg2hw[360]),
		.q(reg2hw[361]),
		.qs()
	);
	// Trace: design.sv:59602:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_21_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_21_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_21_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_21(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_21_we),
		.wd(gpio_toggle_gpio_toggle_21_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_21_ext_d_0),
		.qre(),
		.qe(reg2hw[362]),
		.q(reg2hw[363]),
		.qs()
	);
	// Trace: design.sv:59617:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_22_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_22_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_22_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_22(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_22_we),
		.wd(gpio_toggle_gpio_toggle_22_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_22_ext_d_0),
		.qre(),
		.qe(reg2hw[364]),
		.q(reg2hw[365]),
		.qs()
	);
	// Trace: design.sv:59632:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_23_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_23_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_23_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_23(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_23_we),
		.wd(gpio_toggle_gpio_toggle_23_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_23_ext_d_0),
		.qre(),
		.qe(reg2hw[366]),
		.q(reg2hw[367]),
		.qs()
	);
	// Trace: design.sv:59647:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_24_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_24_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_24_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_24(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_24_we),
		.wd(gpio_toggle_gpio_toggle_24_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_24_ext_d_0),
		.qre(),
		.qe(reg2hw[368]),
		.q(reg2hw[369]),
		.qs()
	);
	// Trace: design.sv:59662:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_25_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_25_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_25_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_25(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_25_we),
		.wd(gpio_toggle_gpio_toggle_25_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_25_ext_d_0),
		.qre(),
		.qe(reg2hw[370]),
		.q(reg2hw[371]),
		.qs()
	);
	// Trace: design.sv:59677:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_26_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_26_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_26_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_26(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_26_we),
		.wd(gpio_toggle_gpio_toggle_26_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_26_ext_d_0),
		.qre(),
		.qe(reg2hw[372]),
		.q(reg2hw[373]),
		.qs()
	);
	// Trace: design.sv:59692:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_27_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_27_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_27_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_27(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_27_we),
		.wd(gpio_toggle_gpio_toggle_27_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_27_ext_d_0),
		.qre(),
		.qe(reg2hw[374]),
		.q(reg2hw[375]),
		.qs()
	);
	// Trace: design.sv:59707:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_28_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_28_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_28_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_28(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_28_we),
		.wd(gpio_toggle_gpio_toggle_28_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_28_ext_d_0),
		.qre(),
		.qe(reg2hw[376]),
		.q(reg2hw[377]),
		.qs()
	);
	// Trace: design.sv:59722:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_29_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_29_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_29_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_29(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_29_we),
		.wd(gpio_toggle_gpio_toggle_29_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_29_ext_d_0),
		.qre(),
		.qe(reg2hw[378]),
		.q(reg2hw[379]),
		.qs()
	);
	// Trace: design.sv:59737:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_30_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_30_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_30_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_30(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_30_we),
		.wd(gpio_toggle_gpio_toggle_30_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_30_ext_d_0),
		.qre(),
		.qe(reg2hw[380]),
		.q(reg2hw[381]),
		.qs()
	);
	// Trace: design.sv:59752:3
	localparam [31:0] sv2v_uu_u_gpio_toggle_gpio_toggle_31_DW = 1;
	// removed localparam type sv2v_uu_u_gpio_toggle_gpio_toggle_31_d
	localparam [0:0] sv2v_uu_u_gpio_toggle_gpio_toggle_31_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_gpio_toggle_gpio_toggle_31(
		.re(1'b0),
		.we(gpio_toggle_gpio_toggle_31_we),
		.wd(gpio_toggle_gpio_toggle_31_wd),
		.d(sv2v_uu_u_gpio_toggle_gpio_toggle_31_ext_d_0),
		.qre(),
		.qe(reg2hw[382]),
		.q(reg2hw[383]),
		.qs()
	);
	// Trace: design.sv:59772:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_0_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_0_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_0_we),
		.wd(intrpt_rise_en_intrpt_rise_en_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_0_ext_d_0),
		.qe(),
		.q(reg2hw[288]),
		.qs(intrpt_rise_en_intrpt_rise_en_0_qs)
	);
	// Trace: design.sv:59798:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_1_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_1_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_1_we),
		.wd(intrpt_rise_en_intrpt_rise_en_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_1_ext_d_0),
		.qe(),
		.q(reg2hw[289]),
		.qs(intrpt_rise_en_intrpt_rise_en_1_qs)
	);
	// Trace: design.sv:59824:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_2_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_2_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_2_we),
		.wd(intrpt_rise_en_intrpt_rise_en_2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_2_ext_d_0),
		.qe(),
		.q(reg2hw[290]),
		.qs(intrpt_rise_en_intrpt_rise_en_2_qs)
	);
	// Trace: design.sv:59850:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_3_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_3_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_3_we),
		.wd(intrpt_rise_en_intrpt_rise_en_3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_3_ext_d_0),
		.qe(),
		.q(reg2hw[291]),
		.qs(intrpt_rise_en_intrpt_rise_en_3_qs)
	);
	// Trace: design.sv:59876:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_4_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_4_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_4_we),
		.wd(intrpt_rise_en_intrpt_rise_en_4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_4_ext_d_0),
		.qe(),
		.q(reg2hw[292]),
		.qs(intrpt_rise_en_intrpt_rise_en_4_qs)
	);
	// Trace: design.sv:59902:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_5_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_5_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_5_we),
		.wd(intrpt_rise_en_intrpt_rise_en_5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_5_ext_d_0),
		.qe(),
		.q(reg2hw[293]),
		.qs(intrpt_rise_en_intrpt_rise_en_5_qs)
	);
	// Trace: design.sv:59928:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_6_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_6_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_6_we),
		.wd(intrpt_rise_en_intrpt_rise_en_6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_6_ext_d_0),
		.qe(),
		.q(reg2hw[294]),
		.qs(intrpt_rise_en_intrpt_rise_en_6_qs)
	);
	// Trace: design.sv:59954:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_7_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_7_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_7_we),
		.wd(intrpt_rise_en_intrpt_rise_en_7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_7_ext_d_0),
		.qe(),
		.q(reg2hw[295]),
		.qs(intrpt_rise_en_intrpt_rise_en_7_qs)
	);
	// Trace: design.sv:59980:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_8_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_8_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_8_we),
		.wd(intrpt_rise_en_intrpt_rise_en_8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_8_ext_d_0),
		.qe(),
		.q(reg2hw[296]),
		.qs(intrpt_rise_en_intrpt_rise_en_8_qs)
	);
	// Trace: design.sv:60006:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_9_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_9_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_9_we),
		.wd(intrpt_rise_en_intrpt_rise_en_9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_9_ext_d_0),
		.qe(),
		.q(reg2hw[297]),
		.qs(intrpt_rise_en_intrpt_rise_en_9_qs)
	);
	// Trace: design.sv:60032:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_10_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_10_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_10_we),
		.wd(intrpt_rise_en_intrpt_rise_en_10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_10_ext_d_0),
		.qe(),
		.q(reg2hw[298]),
		.qs(intrpt_rise_en_intrpt_rise_en_10_qs)
	);
	// Trace: design.sv:60058:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_11_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_11_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_11_we),
		.wd(intrpt_rise_en_intrpt_rise_en_11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_11_ext_d_0),
		.qe(),
		.q(reg2hw[299]),
		.qs(intrpt_rise_en_intrpt_rise_en_11_qs)
	);
	// Trace: design.sv:60084:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_12_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_12_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_12_we),
		.wd(intrpt_rise_en_intrpt_rise_en_12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_12_ext_d_0),
		.qe(),
		.q(reg2hw[300]),
		.qs(intrpt_rise_en_intrpt_rise_en_12_qs)
	);
	// Trace: design.sv:60110:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_13_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_13_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_13_we),
		.wd(intrpt_rise_en_intrpt_rise_en_13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_13_ext_d_0),
		.qe(),
		.q(reg2hw[301]),
		.qs(intrpt_rise_en_intrpt_rise_en_13_qs)
	);
	// Trace: design.sv:60136:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_14_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_14_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_14_we),
		.wd(intrpt_rise_en_intrpt_rise_en_14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_14_ext_d_0),
		.qe(),
		.q(reg2hw[302]),
		.qs(intrpt_rise_en_intrpt_rise_en_14_qs)
	);
	// Trace: design.sv:60162:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_15_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_15_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_15_we),
		.wd(intrpt_rise_en_intrpt_rise_en_15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_15_ext_d_0),
		.qe(),
		.q(reg2hw[303]),
		.qs(intrpt_rise_en_intrpt_rise_en_15_qs)
	);
	// Trace: design.sv:60188:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_16_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_16_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_16_we),
		.wd(intrpt_rise_en_intrpt_rise_en_16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_16_ext_d_0),
		.qe(),
		.q(reg2hw[304]),
		.qs(intrpt_rise_en_intrpt_rise_en_16_qs)
	);
	// Trace: design.sv:60214:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_17_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_17_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_17_we),
		.wd(intrpt_rise_en_intrpt_rise_en_17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_17_ext_d_0),
		.qe(),
		.q(reg2hw[305]),
		.qs(intrpt_rise_en_intrpt_rise_en_17_qs)
	);
	// Trace: design.sv:60240:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_18_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_18_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_18_we),
		.wd(intrpt_rise_en_intrpt_rise_en_18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_18_ext_d_0),
		.qe(),
		.q(reg2hw[306]),
		.qs(intrpt_rise_en_intrpt_rise_en_18_qs)
	);
	// Trace: design.sv:60266:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_19_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_19_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_19_we),
		.wd(intrpt_rise_en_intrpt_rise_en_19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_19_ext_d_0),
		.qe(),
		.q(reg2hw[307]),
		.qs(intrpt_rise_en_intrpt_rise_en_19_qs)
	);
	// Trace: design.sv:60292:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_20_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_20_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_20_we),
		.wd(intrpt_rise_en_intrpt_rise_en_20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_20_ext_d_0),
		.qe(),
		.q(reg2hw[308]),
		.qs(intrpt_rise_en_intrpt_rise_en_20_qs)
	);
	// Trace: design.sv:60318:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_21_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_21_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_21_we),
		.wd(intrpt_rise_en_intrpt_rise_en_21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_21_ext_d_0),
		.qe(),
		.q(reg2hw[309]),
		.qs(intrpt_rise_en_intrpt_rise_en_21_qs)
	);
	// Trace: design.sv:60344:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_22_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_22_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_22_we),
		.wd(intrpt_rise_en_intrpt_rise_en_22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_22_ext_d_0),
		.qe(),
		.q(reg2hw[310]),
		.qs(intrpt_rise_en_intrpt_rise_en_22_qs)
	);
	// Trace: design.sv:60370:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_23_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_23_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_23_we),
		.wd(intrpt_rise_en_intrpt_rise_en_23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_23_ext_d_0),
		.qe(),
		.q(reg2hw[311]),
		.qs(intrpt_rise_en_intrpt_rise_en_23_qs)
	);
	// Trace: design.sv:60396:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_24_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_24_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_24_we),
		.wd(intrpt_rise_en_intrpt_rise_en_24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_24_ext_d_0),
		.qe(),
		.q(reg2hw[312]),
		.qs(intrpt_rise_en_intrpt_rise_en_24_qs)
	);
	// Trace: design.sv:60422:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_25_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_25_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_25_we),
		.wd(intrpt_rise_en_intrpt_rise_en_25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_25_ext_d_0),
		.qe(),
		.q(reg2hw[313]),
		.qs(intrpt_rise_en_intrpt_rise_en_25_qs)
	);
	// Trace: design.sv:60448:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_26_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_26_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_26_we),
		.wd(intrpt_rise_en_intrpt_rise_en_26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_26_ext_d_0),
		.qe(),
		.q(reg2hw[314]),
		.qs(intrpt_rise_en_intrpt_rise_en_26_qs)
	);
	// Trace: design.sv:60474:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_27_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_27_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_27_we),
		.wd(intrpt_rise_en_intrpt_rise_en_27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_27_ext_d_0),
		.qe(),
		.q(reg2hw[315]),
		.qs(intrpt_rise_en_intrpt_rise_en_27_qs)
	);
	// Trace: design.sv:60500:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_28_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_28_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_28_we),
		.wd(intrpt_rise_en_intrpt_rise_en_28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_28_ext_d_0),
		.qe(),
		.q(reg2hw[316]),
		.qs(intrpt_rise_en_intrpt_rise_en_28_qs)
	);
	// Trace: design.sv:60526:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_29_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_29_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_29_we),
		.wd(intrpt_rise_en_intrpt_rise_en_29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_29_ext_d_0),
		.qe(),
		.q(reg2hw[317]),
		.qs(intrpt_rise_en_intrpt_rise_en_29_qs)
	);
	// Trace: design.sv:60552:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_30_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_30_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_30_we),
		.wd(intrpt_rise_en_intrpt_rise_en_30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_30_ext_d_0),
		.qe(),
		.q(reg2hw[318]),
		.qs(intrpt_rise_en_intrpt_rise_en_30_qs)
	);
	// Trace: design.sv:60578:3
	localparam signed [31:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_31_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_31_d
	localparam [0:0] sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_rise_en_intrpt_rise_en_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_en_intrpt_rise_en_31_we),
		.wd(intrpt_rise_en_intrpt_rise_en_31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_rise_en_intrpt_rise_en_31_ext_d_0),
		.qe(),
		.q(reg2hw[319]),
		.qs(intrpt_rise_en_intrpt_rise_en_31_qs)
	);
	// Trace: design.sv:60609:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_0_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_0_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_0_we),
		.wd(intrpt_fall_en_intrpt_fall_en_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_0_ext_d_0),
		.qe(),
		.q(reg2hw[256]),
		.qs(intrpt_fall_en_intrpt_fall_en_0_qs)
	);
	// Trace: design.sv:60635:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_1_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_1_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_1_we),
		.wd(intrpt_fall_en_intrpt_fall_en_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_1_ext_d_0),
		.qe(),
		.q(reg2hw[257]),
		.qs(intrpt_fall_en_intrpt_fall_en_1_qs)
	);
	// Trace: design.sv:60661:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_2_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_2_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_2_we),
		.wd(intrpt_fall_en_intrpt_fall_en_2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_2_ext_d_0),
		.qe(),
		.q(reg2hw[258]),
		.qs(intrpt_fall_en_intrpt_fall_en_2_qs)
	);
	// Trace: design.sv:60687:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_3_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_3_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_3_we),
		.wd(intrpt_fall_en_intrpt_fall_en_3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_3_ext_d_0),
		.qe(),
		.q(reg2hw[259]),
		.qs(intrpt_fall_en_intrpt_fall_en_3_qs)
	);
	// Trace: design.sv:60713:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_4_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_4_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_4_we),
		.wd(intrpt_fall_en_intrpt_fall_en_4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_4_ext_d_0),
		.qe(),
		.q(reg2hw[260]),
		.qs(intrpt_fall_en_intrpt_fall_en_4_qs)
	);
	// Trace: design.sv:60739:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_5_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_5_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_5_we),
		.wd(intrpt_fall_en_intrpt_fall_en_5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_5_ext_d_0),
		.qe(),
		.q(reg2hw[261]),
		.qs(intrpt_fall_en_intrpt_fall_en_5_qs)
	);
	// Trace: design.sv:60765:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_6_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_6_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_6_we),
		.wd(intrpt_fall_en_intrpt_fall_en_6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_6_ext_d_0),
		.qe(),
		.q(reg2hw[262]),
		.qs(intrpt_fall_en_intrpt_fall_en_6_qs)
	);
	// Trace: design.sv:60791:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_7_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_7_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_7_we),
		.wd(intrpt_fall_en_intrpt_fall_en_7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_7_ext_d_0),
		.qe(),
		.q(reg2hw[263]),
		.qs(intrpt_fall_en_intrpt_fall_en_7_qs)
	);
	// Trace: design.sv:60817:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_8_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_8_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_8_we),
		.wd(intrpt_fall_en_intrpt_fall_en_8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_8_ext_d_0),
		.qe(),
		.q(reg2hw[264]),
		.qs(intrpt_fall_en_intrpt_fall_en_8_qs)
	);
	// Trace: design.sv:60843:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_9_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_9_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_9_we),
		.wd(intrpt_fall_en_intrpt_fall_en_9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_9_ext_d_0),
		.qe(),
		.q(reg2hw[265]),
		.qs(intrpt_fall_en_intrpt_fall_en_9_qs)
	);
	// Trace: design.sv:60869:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_10_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_10_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_10_we),
		.wd(intrpt_fall_en_intrpt_fall_en_10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_10_ext_d_0),
		.qe(),
		.q(reg2hw[266]),
		.qs(intrpt_fall_en_intrpt_fall_en_10_qs)
	);
	// Trace: design.sv:60895:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_11_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_11_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_11_we),
		.wd(intrpt_fall_en_intrpt_fall_en_11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_11_ext_d_0),
		.qe(),
		.q(reg2hw[267]),
		.qs(intrpt_fall_en_intrpt_fall_en_11_qs)
	);
	// Trace: design.sv:60921:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_12_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_12_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_12_we),
		.wd(intrpt_fall_en_intrpt_fall_en_12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_12_ext_d_0),
		.qe(),
		.q(reg2hw[268]),
		.qs(intrpt_fall_en_intrpt_fall_en_12_qs)
	);
	// Trace: design.sv:60947:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_13_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_13_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_13_we),
		.wd(intrpt_fall_en_intrpt_fall_en_13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_13_ext_d_0),
		.qe(),
		.q(reg2hw[269]),
		.qs(intrpt_fall_en_intrpt_fall_en_13_qs)
	);
	// Trace: design.sv:60973:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_14_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_14_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_14_we),
		.wd(intrpt_fall_en_intrpt_fall_en_14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_14_ext_d_0),
		.qe(),
		.q(reg2hw[270]),
		.qs(intrpt_fall_en_intrpt_fall_en_14_qs)
	);
	// Trace: design.sv:60999:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_15_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_15_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_15_we),
		.wd(intrpt_fall_en_intrpt_fall_en_15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_15_ext_d_0),
		.qe(),
		.q(reg2hw[271]),
		.qs(intrpt_fall_en_intrpt_fall_en_15_qs)
	);
	// Trace: design.sv:61025:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_16_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_16_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_16_we),
		.wd(intrpt_fall_en_intrpt_fall_en_16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_16_ext_d_0),
		.qe(),
		.q(reg2hw[272]),
		.qs(intrpt_fall_en_intrpt_fall_en_16_qs)
	);
	// Trace: design.sv:61051:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_17_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_17_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_17_we),
		.wd(intrpt_fall_en_intrpt_fall_en_17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_17_ext_d_0),
		.qe(),
		.q(reg2hw[273]),
		.qs(intrpt_fall_en_intrpt_fall_en_17_qs)
	);
	// Trace: design.sv:61077:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_18_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_18_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_18_we),
		.wd(intrpt_fall_en_intrpt_fall_en_18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_18_ext_d_0),
		.qe(),
		.q(reg2hw[274]),
		.qs(intrpt_fall_en_intrpt_fall_en_18_qs)
	);
	// Trace: design.sv:61103:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_19_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_19_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_19_we),
		.wd(intrpt_fall_en_intrpt_fall_en_19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_19_ext_d_0),
		.qe(),
		.q(reg2hw[275]),
		.qs(intrpt_fall_en_intrpt_fall_en_19_qs)
	);
	// Trace: design.sv:61129:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_20_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_20_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_20_we),
		.wd(intrpt_fall_en_intrpt_fall_en_20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_20_ext_d_0),
		.qe(),
		.q(reg2hw[276]),
		.qs(intrpt_fall_en_intrpt_fall_en_20_qs)
	);
	// Trace: design.sv:61155:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_21_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_21_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_21_we),
		.wd(intrpt_fall_en_intrpt_fall_en_21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_21_ext_d_0),
		.qe(),
		.q(reg2hw[277]),
		.qs(intrpt_fall_en_intrpt_fall_en_21_qs)
	);
	// Trace: design.sv:61181:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_22_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_22_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_22_we),
		.wd(intrpt_fall_en_intrpt_fall_en_22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_22_ext_d_0),
		.qe(),
		.q(reg2hw[278]),
		.qs(intrpt_fall_en_intrpt_fall_en_22_qs)
	);
	// Trace: design.sv:61207:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_23_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_23_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_23_we),
		.wd(intrpt_fall_en_intrpt_fall_en_23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_23_ext_d_0),
		.qe(),
		.q(reg2hw[279]),
		.qs(intrpt_fall_en_intrpt_fall_en_23_qs)
	);
	// Trace: design.sv:61233:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_24_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_24_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_24_we),
		.wd(intrpt_fall_en_intrpt_fall_en_24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_24_ext_d_0),
		.qe(),
		.q(reg2hw[280]),
		.qs(intrpt_fall_en_intrpt_fall_en_24_qs)
	);
	// Trace: design.sv:61259:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_25_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_25_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_25_we),
		.wd(intrpt_fall_en_intrpt_fall_en_25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_25_ext_d_0),
		.qe(),
		.q(reg2hw[281]),
		.qs(intrpt_fall_en_intrpt_fall_en_25_qs)
	);
	// Trace: design.sv:61285:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_26_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_26_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_26_we),
		.wd(intrpt_fall_en_intrpt_fall_en_26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_26_ext_d_0),
		.qe(),
		.q(reg2hw[282]),
		.qs(intrpt_fall_en_intrpt_fall_en_26_qs)
	);
	// Trace: design.sv:61311:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_27_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_27_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_27_we),
		.wd(intrpt_fall_en_intrpt_fall_en_27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_27_ext_d_0),
		.qe(),
		.q(reg2hw[283]),
		.qs(intrpt_fall_en_intrpt_fall_en_27_qs)
	);
	// Trace: design.sv:61337:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_28_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_28_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_28_we),
		.wd(intrpt_fall_en_intrpt_fall_en_28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_28_ext_d_0),
		.qe(),
		.q(reg2hw[284]),
		.qs(intrpt_fall_en_intrpt_fall_en_28_qs)
	);
	// Trace: design.sv:61363:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_29_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_29_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_29_we),
		.wd(intrpt_fall_en_intrpt_fall_en_29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_29_ext_d_0),
		.qe(),
		.q(reg2hw[285]),
		.qs(intrpt_fall_en_intrpt_fall_en_29_qs)
	);
	// Trace: design.sv:61389:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_30_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_30_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_30_we),
		.wd(intrpt_fall_en_intrpt_fall_en_30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_30_ext_d_0),
		.qe(),
		.q(reg2hw[286]),
		.qs(intrpt_fall_en_intrpt_fall_en_30_qs)
	);
	// Trace: design.sv:61415:3
	localparam signed [31:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_31_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_31_d
	localparam [0:0] sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_fall_en_intrpt_fall_en_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_en_intrpt_fall_en_31_we),
		.wd(intrpt_fall_en_intrpt_fall_en_31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_fall_en_intrpt_fall_en_31_ext_d_0),
		.qe(),
		.q(reg2hw[287]),
		.qs(intrpt_fall_en_intrpt_fall_en_31_qs)
	);
	// Trace: design.sv:61446:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_0_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_0_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_0_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_0_ext_d_0),
		.qe(),
		.q(reg2hw[224]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_0_qs)
	);
	// Trace: design.sv:61472:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_1_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_1_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_1_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_1_ext_d_0),
		.qe(),
		.q(reg2hw[225]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_1_qs)
	);
	// Trace: design.sv:61498:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_2_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_2_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_2_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_2_ext_d_0),
		.qe(),
		.q(reg2hw[226]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_2_qs)
	);
	// Trace: design.sv:61524:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_3_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_3_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_3_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_3_ext_d_0),
		.qe(),
		.q(reg2hw[227]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_3_qs)
	);
	// Trace: design.sv:61550:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_4_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_4_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_4_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_4_ext_d_0),
		.qe(),
		.q(reg2hw[228]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_4_qs)
	);
	// Trace: design.sv:61576:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_5_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_5_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_5_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_5_ext_d_0),
		.qe(),
		.q(reg2hw[229]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_5_qs)
	);
	// Trace: design.sv:61602:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_6_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_6_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_6_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_6_ext_d_0),
		.qe(),
		.q(reg2hw[230]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_6_qs)
	);
	// Trace: design.sv:61628:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_7_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_7_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_7_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_7_ext_d_0),
		.qe(),
		.q(reg2hw[231]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_7_qs)
	);
	// Trace: design.sv:61654:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_8_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_8_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_8_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_8_ext_d_0),
		.qe(),
		.q(reg2hw[232]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_8_qs)
	);
	// Trace: design.sv:61680:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_9_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_9_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_9_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_9_ext_d_0),
		.qe(),
		.q(reg2hw[233]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_9_qs)
	);
	// Trace: design.sv:61706:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_10_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_10_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_10_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_10_ext_d_0),
		.qe(),
		.q(reg2hw[234]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_10_qs)
	);
	// Trace: design.sv:61732:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_11_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_11_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_11_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_11_ext_d_0),
		.qe(),
		.q(reg2hw[235]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_11_qs)
	);
	// Trace: design.sv:61758:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_12_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_12_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_12_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_12_ext_d_0),
		.qe(),
		.q(reg2hw[236]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_12_qs)
	);
	// Trace: design.sv:61784:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_13_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_13_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_13_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_13_ext_d_0),
		.qe(),
		.q(reg2hw[237]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_13_qs)
	);
	// Trace: design.sv:61810:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_14_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_14_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_14_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_14_ext_d_0),
		.qe(),
		.q(reg2hw[238]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_14_qs)
	);
	// Trace: design.sv:61836:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_15_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_15_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_15_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_15_ext_d_0),
		.qe(),
		.q(reg2hw[239]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_15_qs)
	);
	// Trace: design.sv:61862:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_16_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_16_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_16_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_16_ext_d_0),
		.qe(),
		.q(reg2hw[240]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_16_qs)
	);
	// Trace: design.sv:61888:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_17_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_17_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_17_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_17_ext_d_0),
		.qe(),
		.q(reg2hw[241]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_17_qs)
	);
	// Trace: design.sv:61914:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_18_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_18_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_18_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_18_ext_d_0),
		.qe(),
		.q(reg2hw[242]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_18_qs)
	);
	// Trace: design.sv:61940:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_19_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_19_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_19_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_19_ext_d_0),
		.qe(),
		.q(reg2hw[243]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_19_qs)
	);
	// Trace: design.sv:61966:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_20_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_20_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_20_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_20_ext_d_0),
		.qe(),
		.q(reg2hw[244]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_20_qs)
	);
	// Trace: design.sv:61992:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_21_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_21_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_21_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_21_ext_d_0),
		.qe(),
		.q(reg2hw[245]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_21_qs)
	);
	// Trace: design.sv:62018:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_22_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_22_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_22_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_22_ext_d_0),
		.qe(),
		.q(reg2hw[246]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_22_qs)
	);
	// Trace: design.sv:62044:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_23_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_23_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_23_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_23_ext_d_0),
		.qe(),
		.q(reg2hw[247]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_23_qs)
	);
	// Trace: design.sv:62070:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_24_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_24_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_24_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_24_ext_d_0),
		.qe(),
		.q(reg2hw[248]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_24_qs)
	);
	// Trace: design.sv:62096:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_25_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_25_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_25_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_25_ext_d_0),
		.qe(),
		.q(reg2hw[249]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_25_qs)
	);
	// Trace: design.sv:62122:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_26_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_26_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_26_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_26_ext_d_0),
		.qe(),
		.q(reg2hw[250]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_26_qs)
	);
	// Trace: design.sv:62148:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_27_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_27_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_27_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_27_ext_d_0),
		.qe(),
		.q(reg2hw[251]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_27_qs)
	);
	// Trace: design.sv:62174:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_28_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_28_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_28_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_28_ext_d_0),
		.qe(),
		.q(reg2hw[252]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_28_qs)
	);
	// Trace: design.sv:62200:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_29_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_29_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_29_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_29_ext_d_0),
		.qe(),
		.q(reg2hw[253]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_29_qs)
	);
	// Trace: design.sv:62226:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_30_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_30_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_30_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_30_ext_d_0),
		.qe(),
		.q(reg2hw[254]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_30_qs)
	);
	// Trace: design.sv:62252:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_31_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_31_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_en_intrpt_lvl_high_en_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_en_intrpt_lvl_high_en_31_we),
		.wd(intrpt_lvl_high_en_intrpt_lvl_high_en_31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_high_en_intrpt_lvl_high_en_31_ext_d_0),
		.qe(),
		.q(reg2hw[255]),
		.qs(intrpt_lvl_high_en_intrpt_lvl_high_en_31_qs)
	);
	// Trace: design.sv:62283:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_0_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_0_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_0_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_0_ext_d_0),
		.qe(),
		.q(reg2hw[192]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_0_qs)
	);
	// Trace: design.sv:62309:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_1_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_1_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_1_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_1_ext_d_0),
		.qe(),
		.q(reg2hw[193]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_1_qs)
	);
	// Trace: design.sv:62335:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_2_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_2_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_2_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_2_ext_d_0),
		.qe(),
		.q(reg2hw[194]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_2_qs)
	);
	// Trace: design.sv:62361:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_3_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_3_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_3_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_3_ext_d_0),
		.qe(),
		.q(reg2hw[195]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_3_qs)
	);
	// Trace: design.sv:62387:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_4_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_4_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_4_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_4_ext_d_0),
		.qe(),
		.q(reg2hw[196]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_4_qs)
	);
	// Trace: design.sv:62413:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_5_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_5_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_5_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_5_ext_d_0),
		.qe(),
		.q(reg2hw[197]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_5_qs)
	);
	// Trace: design.sv:62439:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_6_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_6_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_6_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_6_ext_d_0),
		.qe(),
		.q(reg2hw[198]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_6_qs)
	);
	// Trace: design.sv:62465:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_7_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_7_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_7_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_7_ext_d_0),
		.qe(),
		.q(reg2hw[199]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_7_qs)
	);
	// Trace: design.sv:62491:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_8_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_8_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_8_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_8_ext_d_0),
		.qe(),
		.q(reg2hw[200]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_8_qs)
	);
	// Trace: design.sv:62517:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_9_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_9_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_9_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_9_ext_d_0),
		.qe(),
		.q(reg2hw[201]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_9_qs)
	);
	// Trace: design.sv:62543:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_10_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_10_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_10_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_10_ext_d_0),
		.qe(),
		.q(reg2hw[202]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_10_qs)
	);
	// Trace: design.sv:62569:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_11_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_11_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_11_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_11_ext_d_0),
		.qe(),
		.q(reg2hw[203]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_11_qs)
	);
	// Trace: design.sv:62595:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_12_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_12_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_12_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_12_ext_d_0),
		.qe(),
		.q(reg2hw[204]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_12_qs)
	);
	// Trace: design.sv:62621:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_13_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_13_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_13_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_13_ext_d_0),
		.qe(),
		.q(reg2hw[205]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_13_qs)
	);
	// Trace: design.sv:62647:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_14_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_14_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_14_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_14_ext_d_0),
		.qe(),
		.q(reg2hw[206]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_14_qs)
	);
	// Trace: design.sv:62673:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_15_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_15_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_15_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_15_ext_d_0),
		.qe(),
		.q(reg2hw[207]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_15_qs)
	);
	// Trace: design.sv:62699:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_16_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_16_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_16_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_16_ext_d_0),
		.qe(),
		.q(reg2hw[208]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_16_qs)
	);
	// Trace: design.sv:62725:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_17_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_17_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_17_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_17_ext_d_0),
		.qe(),
		.q(reg2hw[209]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_17_qs)
	);
	// Trace: design.sv:62751:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_18_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_18_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_18_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_18_ext_d_0),
		.qe(),
		.q(reg2hw[210]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_18_qs)
	);
	// Trace: design.sv:62777:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_19_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_19_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_19_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_19_ext_d_0),
		.qe(),
		.q(reg2hw[211]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_19_qs)
	);
	// Trace: design.sv:62803:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_20_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_20_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_20_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_20_ext_d_0),
		.qe(),
		.q(reg2hw[212]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_20_qs)
	);
	// Trace: design.sv:62829:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_21_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_21_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_21_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_21_ext_d_0),
		.qe(),
		.q(reg2hw[213]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_21_qs)
	);
	// Trace: design.sv:62855:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_22_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_22_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_22_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_22_ext_d_0),
		.qe(),
		.q(reg2hw[214]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_22_qs)
	);
	// Trace: design.sv:62881:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_23_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_23_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_23_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_23_ext_d_0),
		.qe(),
		.q(reg2hw[215]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_23_qs)
	);
	// Trace: design.sv:62907:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_24_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_24_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_24_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_24_ext_d_0),
		.qe(),
		.q(reg2hw[216]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_24_qs)
	);
	// Trace: design.sv:62933:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_25_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_25_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_25_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_25_ext_d_0),
		.qe(),
		.q(reg2hw[217]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_25_qs)
	);
	// Trace: design.sv:62959:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_26_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_26_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_26_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_26_ext_d_0),
		.qe(),
		.q(reg2hw[218]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_26_qs)
	);
	// Trace: design.sv:62985:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_27_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_27_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_27_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_27_ext_d_0),
		.qe(),
		.q(reg2hw[219]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_27_qs)
	);
	// Trace: design.sv:63011:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_28_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_28_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_28_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_28_ext_d_0),
		.qe(),
		.q(reg2hw[220]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_28_qs)
	);
	// Trace: design.sv:63037:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_29_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_29_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_29_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_29_ext_d_0),
		.qe(),
		.q(reg2hw[221]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_29_qs)
	);
	// Trace: design.sv:63063:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_30_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_30_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_30_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_30_ext_d_0),
		.qe(),
		.q(reg2hw[222]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_30_qs)
	);
	// Trace: design.sv:63089:3
	localparam signed [31:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_31_DW = 1;
	// removed localparam type sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_31_d
	localparam [0:0] sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_en_intrpt_lvl_low_en_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_en_intrpt_lvl_low_en_31_we),
		.wd(intrpt_lvl_low_en_intrpt_lvl_low_en_31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intrpt_lvl_low_en_intrpt_lvl_low_en_31_ext_d_0),
		.qe(),
		.q(reg2hw[223]),
		.qs(intrpt_lvl_low_en_intrpt_lvl_low_en_31_qs)
	);
	// Trace: design.sv:63120:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_0(
		.re(intrpt_status_intrpt_status_0_re),
		.we(intrpt_status_intrpt_status_0_we),
		.wd(intrpt_status_intrpt_status_0_wd),
		.d(hw2reg[256]),
		.qre(),
		.qe(reg2hw[128]),
		.q(reg2hw[129]),
		.qs(intrpt_status_intrpt_status_0_qs)
	);
	// Trace: design.sv:63135:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_1(
		.re(intrpt_status_intrpt_status_1_re),
		.we(intrpt_status_intrpt_status_1_we),
		.wd(intrpt_status_intrpt_status_1_wd),
		.d(hw2reg[257]),
		.qre(),
		.qe(reg2hw[130]),
		.q(reg2hw[131]),
		.qs(intrpt_status_intrpt_status_1_qs)
	);
	// Trace: design.sv:63150:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_2(
		.re(intrpt_status_intrpt_status_2_re),
		.we(intrpt_status_intrpt_status_2_we),
		.wd(intrpt_status_intrpt_status_2_wd),
		.d(hw2reg[258]),
		.qre(),
		.qe(reg2hw[132]),
		.q(reg2hw[133]),
		.qs(intrpt_status_intrpt_status_2_qs)
	);
	// Trace: design.sv:63165:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_3(
		.re(intrpt_status_intrpt_status_3_re),
		.we(intrpt_status_intrpt_status_3_we),
		.wd(intrpt_status_intrpt_status_3_wd),
		.d(hw2reg[259]),
		.qre(),
		.qe(reg2hw[134]),
		.q(reg2hw[135]),
		.qs(intrpt_status_intrpt_status_3_qs)
	);
	// Trace: design.sv:63180:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_4(
		.re(intrpt_status_intrpt_status_4_re),
		.we(intrpt_status_intrpt_status_4_we),
		.wd(intrpt_status_intrpt_status_4_wd),
		.d(hw2reg[260]),
		.qre(),
		.qe(reg2hw[136]),
		.q(reg2hw[137]),
		.qs(intrpt_status_intrpt_status_4_qs)
	);
	// Trace: design.sv:63195:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_5(
		.re(intrpt_status_intrpt_status_5_re),
		.we(intrpt_status_intrpt_status_5_we),
		.wd(intrpt_status_intrpt_status_5_wd),
		.d(hw2reg[261]),
		.qre(),
		.qe(reg2hw[138]),
		.q(reg2hw[139]),
		.qs(intrpt_status_intrpt_status_5_qs)
	);
	// Trace: design.sv:63210:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_6(
		.re(intrpt_status_intrpt_status_6_re),
		.we(intrpt_status_intrpt_status_6_we),
		.wd(intrpt_status_intrpt_status_6_wd),
		.d(hw2reg[262]),
		.qre(),
		.qe(reg2hw[140]),
		.q(reg2hw[141]),
		.qs(intrpt_status_intrpt_status_6_qs)
	);
	// Trace: design.sv:63225:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_7(
		.re(intrpt_status_intrpt_status_7_re),
		.we(intrpt_status_intrpt_status_7_we),
		.wd(intrpt_status_intrpt_status_7_wd),
		.d(hw2reg[263]),
		.qre(),
		.qe(reg2hw[142]),
		.q(reg2hw[143]),
		.qs(intrpt_status_intrpt_status_7_qs)
	);
	// Trace: design.sv:63240:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_8(
		.re(intrpt_status_intrpt_status_8_re),
		.we(intrpt_status_intrpt_status_8_we),
		.wd(intrpt_status_intrpt_status_8_wd),
		.d(hw2reg[264]),
		.qre(),
		.qe(reg2hw[144]),
		.q(reg2hw[145]),
		.qs(intrpt_status_intrpt_status_8_qs)
	);
	// Trace: design.sv:63255:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_9(
		.re(intrpt_status_intrpt_status_9_re),
		.we(intrpt_status_intrpt_status_9_we),
		.wd(intrpt_status_intrpt_status_9_wd),
		.d(hw2reg[265]),
		.qre(),
		.qe(reg2hw[146]),
		.q(reg2hw[147]),
		.qs(intrpt_status_intrpt_status_9_qs)
	);
	// Trace: design.sv:63270:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_10(
		.re(intrpt_status_intrpt_status_10_re),
		.we(intrpt_status_intrpt_status_10_we),
		.wd(intrpt_status_intrpt_status_10_wd),
		.d(hw2reg[266]),
		.qre(),
		.qe(reg2hw[148]),
		.q(reg2hw[149]),
		.qs(intrpt_status_intrpt_status_10_qs)
	);
	// Trace: design.sv:63285:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_11(
		.re(intrpt_status_intrpt_status_11_re),
		.we(intrpt_status_intrpt_status_11_we),
		.wd(intrpt_status_intrpt_status_11_wd),
		.d(hw2reg[267]),
		.qre(),
		.qe(reg2hw[150]),
		.q(reg2hw[151]),
		.qs(intrpt_status_intrpt_status_11_qs)
	);
	// Trace: design.sv:63300:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_12(
		.re(intrpt_status_intrpt_status_12_re),
		.we(intrpt_status_intrpt_status_12_we),
		.wd(intrpt_status_intrpt_status_12_wd),
		.d(hw2reg[268]),
		.qre(),
		.qe(reg2hw[152]),
		.q(reg2hw[153]),
		.qs(intrpt_status_intrpt_status_12_qs)
	);
	// Trace: design.sv:63315:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_13(
		.re(intrpt_status_intrpt_status_13_re),
		.we(intrpt_status_intrpt_status_13_we),
		.wd(intrpt_status_intrpt_status_13_wd),
		.d(hw2reg[269]),
		.qre(),
		.qe(reg2hw[154]),
		.q(reg2hw[155]),
		.qs(intrpt_status_intrpt_status_13_qs)
	);
	// Trace: design.sv:63330:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_14(
		.re(intrpt_status_intrpt_status_14_re),
		.we(intrpt_status_intrpt_status_14_we),
		.wd(intrpt_status_intrpt_status_14_wd),
		.d(hw2reg[270]),
		.qre(),
		.qe(reg2hw[156]),
		.q(reg2hw[157]),
		.qs(intrpt_status_intrpt_status_14_qs)
	);
	// Trace: design.sv:63345:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_15(
		.re(intrpt_status_intrpt_status_15_re),
		.we(intrpt_status_intrpt_status_15_we),
		.wd(intrpt_status_intrpt_status_15_wd),
		.d(hw2reg[271]),
		.qre(),
		.qe(reg2hw[158]),
		.q(reg2hw[159]),
		.qs(intrpt_status_intrpt_status_15_qs)
	);
	// Trace: design.sv:63360:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_16(
		.re(intrpt_status_intrpt_status_16_re),
		.we(intrpt_status_intrpt_status_16_we),
		.wd(intrpt_status_intrpt_status_16_wd),
		.d(hw2reg[272]),
		.qre(),
		.qe(reg2hw[160]),
		.q(reg2hw[161]),
		.qs(intrpt_status_intrpt_status_16_qs)
	);
	// Trace: design.sv:63375:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_17(
		.re(intrpt_status_intrpt_status_17_re),
		.we(intrpt_status_intrpt_status_17_we),
		.wd(intrpt_status_intrpt_status_17_wd),
		.d(hw2reg[273]),
		.qre(),
		.qe(reg2hw[162]),
		.q(reg2hw[163]),
		.qs(intrpt_status_intrpt_status_17_qs)
	);
	// Trace: design.sv:63390:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_18(
		.re(intrpt_status_intrpt_status_18_re),
		.we(intrpt_status_intrpt_status_18_we),
		.wd(intrpt_status_intrpt_status_18_wd),
		.d(hw2reg[274]),
		.qre(),
		.qe(reg2hw[164]),
		.q(reg2hw[165]),
		.qs(intrpt_status_intrpt_status_18_qs)
	);
	// Trace: design.sv:63405:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_19(
		.re(intrpt_status_intrpt_status_19_re),
		.we(intrpt_status_intrpt_status_19_we),
		.wd(intrpt_status_intrpt_status_19_wd),
		.d(hw2reg[275]),
		.qre(),
		.qe(reg2hw[166]),
		.q(reg2hw[167]),
		.qs(intrpt_status_intrpt_status_19_qs)
	);
	// Trace: design.sv:63420:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_20(
		.re(intrpt_status_intrpt_status_20_re),
		.we(intrpt_status_intrpt_status_20_we),
		.wd(intrpt_status_intrpt_status_20_wd),
		.d(hw2reg[276]),
		.qre(),
		.qe(reg2hw[168]),
		.q(reg2hw[169]),
		.qs(intrpt_status_intrpt_status_20_qs)
	);
	// Trace: design.sv:63435:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_21(
		.re(intrpt_status_intrpt_status_21_re),
		.we(intrpt_status_intrpt_status_21_we),
		.wd(intrpt_status_intrpt_status_21_wd),
		.d(hw2reg[277]),
		.qre(),
		.qe(reg2hw[170]),
		.q(reg2hw[171]),
		.qs(intrpt_status_intrpt_status_21_qs)
	);
	// Trace: design.sv:63450:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_22(
		.re(intrpt_status_intrpt_status_22_re),
		.we(intrpt_status_intrpt_status_22_we),
		.wd(intrpt_status_intrpt_status_22_wd),
		.d(hw2reg[278]),
		.qre(),
		.qe(reg2hw[172]),
		.q(reg2hw[173]),
		.qs(intrpt_status_intrpt_status_22_qs)
	);
	// Trace: design.sv:63465:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_23(
		.re(intrpt_status_intrpt_status_23_re),
		.we(intrpt_status_intrpt_status_23_we),
		.wd(intrpt_status_intrpt_status_23_wd),
		.d(hw2reg[279]),
		.qre(),
		.qe(reg2hw[174]),
		.q(reg2hw[175]),
		.qs(intrpt_status_intrpt_status_23_qs)
	);
	// Trace: design.sv:63480:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_24(
		.re(intrpt_status_intrpt_status_24_re),
		.we(intrpt_status_intrpt_status_24_we),
		.wd(intrpt_status_intrpt_status_24_wd),
		.d(hw2reg[280]),
		.qre(),
		.qe(reg2hw[176]),
		.q(reg2hw[177]),
		.qs(intrpt_status_intrpt_status_24_qs)
	);
	// Trace: design.sv:63495:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_25(
		.re(intrpt_status_intrpt_status_25_re),
		.we(intrpt_status_intrpt_status_25_we),
		.wd(intrpt_status_intrpt_status_25_wd),
		.d(hw2reg[281]),
		.qre(),
		.qe(reg2hw[178]),
		.q(reg2hw[179]),
		.qs(intrpt_status_intrpt_status_25_qs)
	);
	// Trace: design.sv:63510:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_26(
		.re(intrpt_status_intrpt_status_26_re),
		.we(intrpt_status_intrpt_status_26_we),
		.wd(intrpt_status_intrpt_status_26_wd),
		.d(hw2reg[282]),
		.qre(),
		.qe(reg2hw[180]),
		.q(reg2hw[181]),
		.qs(intrpt_status_intrpt_status_26_qs)
	);
	// Trace: design.sv:63525:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_27(
		.re(intrpt_status_intrpt_status_27_re),
		.we(intrpt_status_intrpt_status_27_we),
		.wd(intrpt_status_intrpt_status_27_wd),
		.d(hw2reg[283]),
		.qre(),
		.qe(reg2hw[182]),
		.q(reg2hw[183]),
		.qs(intrpt_status_intrpt_status_27_qs)
	);
	// Trace: design.sv:63540:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_28(
		.re(intrpt_status_intrpt_status_28_re),
		.we(intrpt_status_intrpt_status_28_we),
		.wd(intrpt_status_intrpt_status_28_wd),
		.d(hw2reg[284]),
		.qre(),
		.qe(reg2hw[184]),
		.q(reg2hw[185]),
		.qs(intrpt_status_intrpt_status_28_qs)
	);
	// Trace: design.sv:63555:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_29(
		.re(intrpt_status_intrpt_status_29_re),
		.we(intrpt_status_intrpt_status_29_we),
		.wd(intrpt_status_intrpt_status_29_wd),
		.d(hw2reg[285]),
		.qre(),
		.qe(reg2hw[186]),
		.q(reg2hw[187]),
		.qs(intrpt_status_intrpt_status_29_qs)
	);
	// Trace: design.sv:63570:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_30(
		.re(intrpt_status_intrpt_status_30_re),
		.we(intrpt_status_intrpt_status_30_we),
		.wd(intrpt_status_intrpt_status_30_wd),
		.d(hw2reg[286]),
		.qre(),
		.qe(reg2hw[188]),
		.q(reg2hw[189]),
		.qs(intrpt_status_intrpt_status_30_qs)
	);
	// Trace: design.sv:63585:3
	prim_subreg_ext #(.DW(1)) u_intrpt_status_intrpt_status_31(
		.re(intrpt_status_intrpt_status_31_re),
		.we(intrpt_status_intrpt_status_31_we),
		.wd(intrpt_status_intrpt_status_31_wd),
		.d(hw2reg[287]),
		.qre(),
		.qe(reg2hw[190]),
		.q(reg2hw[191]),
		.qs(intrpt_status_intrpt_status_31_qs)
	);
	// Trace: design.sv:63605:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_0_we),
		.wd(intrpt_rise_status_intrpt_rise_status_0_wd),
		.de(hw2reg[192]),
		.d(hw2reg[193]),
		.qe(),
		.q(reg2hw[96]),
		.qs(intrpt_rise_status_intrpt_rise_status_0_qs)
	);
	// Trace: design.sv:63631:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_1_we),
		.wd(intrpt_rise_status_intrpt_rise_status_1_wd),
		.de(hw2reg[194]),
		.d(hw2reg[195]),
		.qe(),
		.q(reg2hw[97]),
		.qs(intrpt_rise_status_intrpt_rise_status_1_qs)
	);
	// Trace: design.sv:63657:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_2_we),
		.wd(intrpt_rise_status_intrpt_rise_status_2_wd),
		.de(hw2reg[196]),
		.d(hw2reg[197]),
		.qe(),
		.q(reg2hw[98]),
		.qs(intrpt_rise_status_intrpt_rise_status_2_qs)
	);
	// Trace: design.sv:63683:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_3_we),
		.wd(intrpt_rise_status_intrpt_rise_status_3_wd),
		.de(hw2reg[198]),
		.d(hw2reg[199]),
		.qe(),
		.q(reg2hw[99]),
		.qs(intrpt_rise_status_intrpt_rise_status_3_qs)
	);
	// Trace: design.sv:63709:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_4_we),
		.wd(intrpt_rise_status_intrpt_rise_status_4_wd),
		.de(hw2reg[200]),
		.d(hw2reg[201]),
		.qe(),
		.q(reg2hw[100]),
		.qs(intrpt_rise_status_intrpt_rise_status_4_qs)
	);
	// Trace: design.sv:63735:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_5_we),
		.wd(intrpt_rise_status_intrpt_rise_status_5_wd),
		.de(hw2reg[202]),
		.d(hw2reg[203]),
		.qe(),
		.q(reg2hw[101]),
		.qs(intrpt_rise_status_intrpt_rise_status_5_qs)
	);
	// Trace: design.sv:63761:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_6_we),
		.wd(intrpt_rise_status_intrpt_rise_status_6_wd),
		.de(hw2reg[204]),
		.d(hw2reg[205]),
		.qe(),
		.q(reg2hw[102]),
		.qs(intrpt_rise_status_intrpt_rise_status_6_qs)
	);
	// Trace: design.sv:63787:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_7_we),
		.wd(intrpt_rise_status_intrpt_rise_status_7_wd),
		.de(hw2reg[206]),
		.d(hw2reg[207]),
		.qe(),
		.q(reg2hw[103]),
		.qs(intrpt_rise_status_intrpt_rise_status_7_qs)
	);
	// Trace: design.sv:63813:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_8_we),
		.wd(intrpt_rise_status_intrpt_rise_status_8_wd),
		.de(hw2reg[208]),
		.d(hw2reg[209]),
		.qe(),
		.q(reg2hw[104]),
		.qs(intrpt_rise_status_intrpt_rise_status_8_qs)
	);
	// Trace: design.sv:63839:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_9_we),
		.wd(intrpt_rise_status_intrpt_rise_status_9_wd),
		.de(hw2reg[210]),
		.d(hw2reg[211]),
		.qe(),
		.q(reg2hw[105]),
		.qs(intrpt_rise_status_intrpt_rise_status_9_qs)
	);
	// Trace: design.sv:63865:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_10_we),
		.wd(intrpt_rise_status_intrpt_rise_status_10_wd),
		.de(hw2reg[212]),
		.d(hw2reg[213]),
		.qe(),
		.q(reg2hw[106]),
		.qs(intrpt_rise_status_intrpt_rise_status_10_qs)
	);
	// Trace: design.sv:63891:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_11_we),
		.wd(intrpt_rise_status_intrpt_rise_status_11_wd),
		.de(hw2reg[214]),
		.d(hw2reg[215]),
		.qe(),
		.q(reg2hw[107]),
		.qs(intrpt_rise_status_intrpt_rise_status_11_qs)
	);
	// Trace: design.sv:63917:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_12_we),
		.wd(intrpt_rise_status_intrpt_rise_status_12_wd),
		.de(hw2reg[216]),
		.d(hw2reg[217]),
		.qe(),
		.q(reg2hw[108]),
		.qs(intrpt_rise_status_intrpt_rise_status_12_qs)
	);
	// Trace: design.sv:63943:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_13_we),
		.wd(intrpt_rise_status_intrpt_rise_status_13_wd),
		.de(hw2reg[218]),
		.d(hw2reg[219]),
		.qe(),
		.q(reg2hw[109]),
		.qs(intrpt_rise_status_intrpt_rise_status_13_qs)
	);
	// Trace: design.sv:63969:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_14_we),
		.wd(intrpt_rise_status_intrpt_rise_status_14_wd),
		.de(hw2reg[220]),
		.d(hw2reg[221]),
		.qe(),
		.q(reg2hw[110]),
		.qs(intrpt_rise_status_intrpt_rise_status_14_qs)
	);
	// Trace: design.sv:63995:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_15_we),
		.wd(intrpt_rise_status_intrpt_rise_status_15_wd),
		.de(hw2reg[222]),
		.d(hw2reg[223]),
		.qe(),
		.q(reg2hw[111]),
		.qs(intrpt_rise_status_intrpt_rise_status_15_qs)
	);
	// Trace: design.sv:64021:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_16_we),
		.wd(intrpt_rise_status_intrpt_rise_status_16_wd),
		.de(hw2reg[224]),
		.d(hw2reg[225]),
		.qe(),
		.q(reg2hw[112]),
		.qs(intrpt_rise_status_intrpt_rise_status_16_qs)
	);
	// Trace: design.sv:64047:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_17_we),
		.wd(intrpt_rise_status_intrpt_rise_status_17_wd),
		.de(hw2reg[226]),
		.d(hw2reg[227]),
		.qe(),
		.q(reg2hw[113]),
		.qs(intrpt_rise_status_intrpt_rise_status_17_qs)
	);
	// Trace: design.sv:64073:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_18_we),
		.wd(intrpt_rise_status_intrpt_rise_status_18_wd),
		.de(hw2reg[228]),
		.d(hw2reg[229]),
		.qe(),
		.q(reg2hw[114]),
		.qs(intrpt_rise_status_intrpt_rise_status_18_qs)
	);
	// Trace: design.sv:64099:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_19_we),
		.wd(intrpt_rise_status_intrpt_rise_status_19_wd),
		.de(hw2reg[230]),
		.d(hw2reg[231]),
		.qe(),
		.q(reg2hw[115]),
		.qs(intrpt_rise_status_intrpt_rise_status_19_qs)
	);
	// Trace: design.sv:64125:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_20_we),
		.wd(intrpt_rise_status_intrpt_rise_status_20_wd),
		.de(hw2reg[232]),
		.d(hw2reg[233]),
		.qe(),
		.q(reg2hw[116]),
		.qs(intrpt_rise_status_intrpt_rise_status_20_qs)
	);
	// Trace: design.sv:64151:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_21_we),
		.wd(intrpt_rise_status_intrpt_rise_status_21_wd),
		.de(hw2reg[234]),
		.d(hw2reg[235]),
		.qe(),
		.q(reg2hw[117]),
		.qs(intrpt_rise_status_intrpt_rise_status_21_qs)
	);
	// Trace: design.sv:64177:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_22_we),
		.wd(intrpt_rise_status_intrpt_rise_status_22_wd),
		.de(hw2reg[236]),
		.d(hw2reg[237]),
		.qe(),
		.q(reg2hw[118]),
		.qs(intrpt_rise_status_intrpt_rise_status_22_qs)
	);
	// Trace: design.sv:64203:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_23_we),
		.wd(intrpt_rise_status_intrpt_rise_status_23_wd),
		.de(hw2reg[238]),
		.d(hw2reg[239]),
		.qe(),
		.q(reg2hw[119]),
		.qs(intrpt_rise_status_intrpt_rise_status_23_qs)
	);
	// Trace: design.sv:64229:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_24_we),
		.wd(intrpt_rise_status_intrpt_rise_status_24_wd),
		.de(hw2reg[240]),
		.d(hw2reg[241]),
		.qe(),
		.q(reg2hw[120]),
		.qs(intrpt_rise_status_intrpt_rise_status_24_qs)
	);
	// Trace: design.sv:64255:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_25_we),
		.wd(intrpt_rise_status_intrpt_rise_status_25_wd),
		.de(hw2reg[242]),
		.d(hw2reg[243]),
		.qe(),
		.q(reg2hw[121]),
		.qs(intrpt_rise_status_intrpt_rise_status_25_qs)
	);
	// Trace: design.sv:64281:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_26_we),
		.wd(intrpt_rise_status_intrpt_rise_status_26_wd),
		.de(hw2reg[244]),
		.d(hw2reg[245]),
		.qe(),
		.q(reg2hw[122]),
		.qs(intrpt_rise_status_intrpt_rise_status_26_qs)
	);
	// Trace: design.sv:64307:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_27_we),
		.wd(intrpt_rise_status_intrpt_rise_status_27_wd),
		.de(hw2reg[246]),
		.d(hw2reg[247]),
		.qe(),
		.q(reg2hw[123]),
		.qs(intrpt_rise_status_intrpt_rise_status_27_qs)
	);
	// Trace: design.sv:64333:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_28_we),
		.wd(intrpt_rise_status_intrpt_rise_status_28_wd),
		.de(hw2reg[248]),
		.d(hw2reg[249]),
		.qe(),
		.q(reg2hw[124]),
		.qs(intrpt_rise_status_intrpt_rise_status_28_qs)
	);
	// Trace: design.sv:64359:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_29_we),
		.wd(intrpt_rise_status_intrpt_rise_status_29_wd),
		.de(hw2reg[250]),
		.d(hw2reg[251]),
		.qe(),
		.q(reg2hw[125]),
		.qs(intrpt_rise_status_intrpt_rise_status_29_qs)
	);
	// Trace: design.sv:64385:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_30_we),
		.wd(intrpt_rise_status_intrpt_rise_status_30_wd),
		.de(hw2reg[252]),
		.d(hw2reg[253]),
		.qe(),
		.q(reg2hw[126]),
		.qs(intrpt_rise_status_intrpt_rise_status_30_qs)
	);
	// Trace: design.sv:64411:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_rise_status_intrpt_rise_status_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_rise_status_intrpt_rise_status_31_we),
		.wd(intrpt_rise_status_intrpt_rise_status_31_wd),
		.de(hw2reg[254]),
		.d(hw2reg[255]),
		.qe(),
		.q(reg2hw[127]),
		.qs(intrpt_rise_status_intrpt_rise_status_31_qs)
	);
	// Trace: design.sv:64442:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_0_we),
		.wd(intrpt_fall_status_intrpt_fall_status_0_wd),
		.de(hw2reg[128]),
		.d(hw2reg[129]),
		.qe(),
		.q(reg2hw[64]),
		.qs(intrpt_fall_status_intrpt_fall_status_0_qs)
	);
	// Trace: design.sv:64468:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_1_we),
		.wd(intrpt_fall_status_intrpt_fall_status_1_wd),
		.de(hw2reg[130]),
		.d(hw2reg[131]),
		.qe(),
		.q(reg2hw[65]),
		.qs(intrpt_fall_status_intrpt_fall_status_1_qs)
	);
	// Trace: design.sv:64494:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_2_we),
		.wd(intrpt_fall_status_intrpt_fall_status_2_wd),
		.de(hw2reg[132]),
		.d(hw2reg[133]),
		.qe(),
		.q(reg2hw[66]),
		.qs(intrpt_fall_status_intrpt_fall_status_2_qs)
	);
	// Trace: design.sv:64520:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_3_we),
		.wd(intrpt_fall_status_intrpt_fall_status_3_wd),
		.de(hw2reg[134]),
		.d(hw2reg[135]),
		.qe(),
		.q(reg2hw[67]),
		.qs(intrpt_fall_status_intrpt_fall_status_3_qs)
	);
	// Trace: design.sv:64546:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_4_we),
		.wd(intrpt_fall_status_intrpt_fall_status_4_wd),
		.de(hw2reg[136]),
		.d(hw2reg[137]),
		.qe(),
		.q(reg2hw[68]),
		.qs(intrpt_fall_status_intrpt_fall_status_4_qs)
	);
	// Trace: design.sv:64572:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_5_we),
		.wd(intrpt_fall_status_intrpt_fall_status_5_wd),
		.de(hw2reg[138]),
		.d(hw2reg[139]),
		.qe(),
		.q(reg2hw[69]),
		.qs(intrpt_fall_status_intrpt_fall_status_5_qs)
	);
	// Trace: design.sv:64598:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_6_we),
		.wd(intrpt_fall_status_intrpt_fall_status_6_wd),
		.de(hw2reg[140]),
		.d(hw2reg[141]),
		.qe(),
		.q(reg2hw[70]),
		.qs(intrpt_fall_status_intrpt_fall_status_6_qs)
	);
	// Trace: design.sv:64624:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_7_we),
		.wd(intrpt_fall_status_intrpt_fall_status_7_wd),
		.de(hw2reg[142]),
		.d(hw2reg[143]),
		.qe(),
		.q(reg2hw[71]),
		.qs(intrpt_fall_status_intrpt_fall_status_7_qs)
	);
	// Trace: design.sv:64650:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_8_we),
		.wd(intrpt_fall_status_intrpt_fall_status_8_wd),
		.de(hw2reg[144]),
		.d(hw2reg[145]),
		.qe(),
		.q(reg2hw[72]),
		.qs(intrpt_fall_status_intrpt_fall_status_8_qs)
	);
	// Trace: design.sv:64676:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_9_we),
		.wd(intrpt_fall_status_intrpt_fall_status_9_wd),
		.de(hw2reg[146]),
		.d(hw2reg[147]),
		.qe(),
		.q(reg2hw[73]),
		.qs(intrpt_fall_status_intrpt_fall_status_9_qs)
	);
	// Trace: design.sv:64702:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_10_we),
		.wd(intrpt_fall_status_intrpt_fall_status_10_wd),
		.de(hw2reg[148]),
		.d(hw2reg[149]),
		.qe(),
		.q(reg2hw[74]),
		.qs(intrpt_fall_status_intrpt_fall_status_10_qs)
	);
	// Trace: design.sv:64728:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_11_we),
		.wd(intrpt_fall_status_intrpt_fall_status_11_wd),
		.de(hw2reg[150]),
		.d(hw2reg[151]),
		.qe(),
		.q(reg2hw[75]),
		.qs(intrpt_fall_status_intrpt_fall_status_11_qs)
	);
	// Trace: design.sv:64754:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_12_we),
		.wd(intrpt_fall_status_intrpt_fall_status_12_wd),
		.de(hw2reg[152]),
		.d(hw2reg[153]),
		.qe(),
		.q(reg2hw[76]),
		.qs(intrpt_fall_status_intrpt_fall_status_12_qs)
	);
	// Trace: design.sv:64780:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_13_we),
		.wd(intrpt_fall_status_intrpt_fall_status_13_wd),
		.de(hw2reg[154]),
		.d(hw2reg[155]),
		.qe(),
		.q(reg2hw[77]),
		.qs(intrpt_fall_status_intrpt_fall_status_13_qs)
	);
	// Trace: design.sv:64806:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_14_we),
		.wd(intrpt_fall_status_intrpt_fall_status_14_wd),
		.de(hw2reg[156]),
		.d(hw2reg[157]),
		.qe(),
		.q(reg2hw[78]),
		.qs(intrpt_fall_status_intrpt_fall_status_14_qs)
	);
	// Trace: design.sv:64832:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_15_we),
		.wd(intrpt_fall_status_intrpt_fall_status_15_wd),
		.de(hw2reg[158]),
		.d(hw2reg[159]),
		.qe(),
		.q(reg2hw[79]),
		.qs(intrpt_fall_status_intrpt_fall_status_15_qs)
	);
	// Trace: design.sv:64858:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_16_we),
		.wd(intrpt_fall_status_intrpt_fall_status_16_wd),
		.de(hw2reg[160]),
		.d(hw2reg[161]),
		.qe(),
		.q(reg2hw[80]),
		.qs(intrpt_fall_status_intrpt_fall_status_16_qs)
	);
	// Trace: design.sv:64884:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_17_we),
		.wd(intrpt_fall_status_intrpt_fall_status_17_wd),
		.de(hw2reg[162]),
		.d(hw2reg[163]),
		.qe(),
		.q(reg2hw[81]),
		.qs(intrpt_fall_status_intrpt_fall_status_17_qs)
	);
	// Trace: design.sv:64910:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_18_we),
		.wd(intrpt_fall_status_intrpt_fall_status_18_wd),
		.de(hw2reg[164]),
		.d(hw2reg[165]),
		.qe(),
		.q(reg2hw[82]),
		.qs(intrpt_fall_status_intrpt_fall_status_18_qs)
	);
	// Trace: design.sv:64936:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_19_we),
		.wd(intrpt_fall_status_intrpt_fall_status_19_wd),
		.de(hw2reg[166]),
		.d(hw2reg[167]),
		.qe(),
		.q(reg2hw[83]),
		.qs(intrpt_fall_status_intrpt_fall_status_19_qs)
	);
	// Trace: design.sv:64962:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_20_we),
		.wd(intrpt_fall_status_intrpt_fall_status_20_wd),
		.de(hw2reg[168]),
		.d(hw2reg[169]),
		.qe(),
		.q(reg2hw[84]),
		.qs(intrpt_fall_status_intrpt_fall_status_20_qs)
	);
	// Trace: design.sv:64988:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_21_we),
		.wd(intrpt_fall_status_intrpt_fall_status_21_wd),
		.de(hw2reg[170]),
		.d(hw2reg[171]),
		.qe(),
		.q(reg2hw[85]),
		.qs(intrpt_fall_status_intrpt_fall_status_21_qs)
	);
	// Trace: design.sv:65014:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_22_we),
		.wd(intrpt_fall_status_intrpt_fall_status_22_wd),
		.de(hw2reg[172]),
		.d(hw2reg[173]),
		.qe(),
		.q(reg2hw[86]),
		.qs(intrpt_fall_status_intrpt_fall_status_22_qs)
	);
	// Trace: design.sv:65040:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_23_we),
		.wd(intrpt_fall_status_intrpt_fall_status_23_wd),
		.de(hw2reg[174]),
		.d(hw2reg[175]),
		.qe(),
		.q(reg2hw[87]),
		.qs(intrpt_fall_status_intrpt_fall_status_23_qs)
	);
	// Trace: design.sv:65066:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_24_we),
		.wd(intrpt_fall_status_intrpt_fall_status_24_wd),
		.de(hw2reg[176]),
		.d(hw2reg[177]),
		.qe(),
		.q(reg2hw[88]),
		.qs(intrpt_fall_status_intrpt_fall_status_24_qs)
	);
	// Trace: design.sv:65092:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_25_we),
		.wd(intrpt_fall_status_intrpt_fall_status_25_wd),
		.de(hw2reg[178]),
		.d(hw2reg[179]),
		.qe(),
		.q(reg2hw[89]),
		.qs(intrpt_fall_status_intrpt_fall_status_25_qs)
	);
	// Trace: design.sv:65118:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_26_we),
		.wd(intrpt_fall_status_intrpt_fall_status_26_wd),
		.de(hw2reg[180]),
		.d(hw2reg[181]),
		.qe(),
		.q(reg2hw[90]),
		.qs(intrpt_fall_status_intrpt_fall_status_26_qs)
	);
	// Trace: design.sv:65144:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_27_we),
		.wd(intrpt_fall_status_intrpt_fall_status_27_wd),
		.de(hw2reg[182]),
		.d(hw2reg[183]),
		.qe(),
		.q(reg2hw[91]),
		.qs(intrpt_fall_status_intrpt_fall_status_27_qs)
	);
	// Trace: design.sv:65170:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_28_we),
		.wd(intrpt_fall_status_intrpt_fall_status_28_wd),
		.de(hw2reg[184]),
		.d(hw2reg[185]),
		.qe(),
		.q(reg2hw[92]),
		.qs(intrpt_fall_status_intrpt_fall_status_28_qs)
	);
	// Trace: design.sv:65196:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_29_we),
		.wd(intrpt_fall_status_intrpt_fall_status_29_wd),
		.de(hw2reg[186]),
		.d(hw2reg[187]),
		.qe(),
		.q(reg2hw[93]),
		.qs(intrpt_fall_status_intrpt_fall_status_29_qs)
	);
	// Trace: design.sv:65222:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_30_we),
		.wd(intrpt_fall_status_intrpt_fall_status_30_wd),
		.de(hw2reg[188]),
		.d(hw2reg[189]),
		.qe(),
		.q(reg2hw[94]),
		.qs(intrpt_fall_status_intrpt_fall_status_30_qs)
	);
	// Trace: design.sv:65248:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_fall_status_intrpt_fall_status_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_fall_status_intrpt_fall_status_31_we),
		.wd(intrpt_fall_status_intrpt_fall_status_31_wd),
		.de(hw2reg[190]),
		.d(hw2reg[191]),
		.qe(),
		.q(reg2hw[95]),
		.qs(intrpt_fall_status_intrpt_fall_status_31_qs)
	);
	// Trace: design.sv:65279:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_0_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_0_wd),
		.de(hw2reg[64]),
		.d(hw2reg[65]),
		.qe(),
		.q(reg2hw[32]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_0_qs)
	);
	// Trace: design.sv:65305:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_1_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_1_wd),
		.de(hw2reg[66]),
		.d(hw2reg[67]),
		.qe(),
		.q(reg2hw[33]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_1_qs)
	);
	// Trace: design.sv:65331:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_2_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_2_wd),
		.de(hw2reg[68]),
		.d(hw2reg[69]),
		.qe(),
		.q(reg2hw[34]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_2_qs)
	);
	// Trace: design.sv:65357:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_3_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_3_wd),
		.de(hw2reg[70]),
		.d(hw2reg[71]),
		.qe(),
		.q(reg2hw[35]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_3_qs)
	);
	// Trace: design.sv:65383:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_4_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_4_wd),
		.de(hw2reg[72]),
		.d(hw2reg[73]),
		.qe(),
		.q(reg2hw[36]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_4_qs)
	);
	// Trace: design.sv:65409:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_5_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_5_wd),
		.de(hw2reg[74]),
		.d(hw2reg[75]),
		.qe(),
		.q(reg2hw[37]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_5_qs)
	);
	// Trace: design.sv:65435:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_6_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_6_wd),
		.de(hw2reg[76]),
		.d(hw2reg[77]),
		.qe(),
		.q(reg2hw[38]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_6_qs)
	);
	// Trace: design.sv:65461:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_7_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_7_wd),
		.de(hw2reg[78]),
		.d(hw2reg[79]),
		.qe(),
		.q(reg2hw[39]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_7_qs)
	);
	// Trace: design.sv:65487:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_8_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_8_wd),
		.de(hw2reg[80]),
		.d(hw2reg[81]),
		.qe(),
		.q(reg2hw[40]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_8_qs)
	);
	// Trace: design.sv:65513:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_9_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_9_wd),
		.de(hw2reg[82]),
		.d(hw2reg[83]),
		.qe(),
		.q(reg2hw[41]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_9_qs)
	);
	// Trace: design.sv:65539:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_10_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_10_wd),
		.de(hw2reg[84]),
		.d(hw2reg[85]),
		.qe(),
		.q(reg2hw[42]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_10_qs)
	);
	// Trace: design.sv:65565:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_11_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_11_wd),
		.de(hw2reg[86]),
		.d(hw2reg[87]),
		.qe(),
		.q(reg2hw[43]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_11_qs)
	);
	// Trace: design.sv:65591:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_12_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_12_wd),
		.de(hw2reg[88]),
		.d(hw2reg[89]),
		.qe(),
		.q(reg2hw[44]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_12_qs)
	);
	// Trace: design.sv:65617:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_13_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_13_wd),
		.de(hw2reg[90]),
		.d(hw2reg[91]),
		.qe(),
		.q(reg2hw[45]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_13_qs)
	);
	// Trace: design.sv:65643:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_14_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_14_wd),
		.de(hw2reg[92]),
		.d(hw2reg[93]),
		.qe(),
		.q(reg2hw[46]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_14_qs)
	);
	// Trace: design.sv:65669:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_15_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_15_wd),
		.de(hw2reg[94]),
		.d(hw2reg[95]),
		.qe(),
		.q(reg2hw[47]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_15_qs)
	);
	// Trace: design.sv:65695:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_16_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_16_wd),
		.de(hw2reg[96]),
		.d(hw2reg[97]),
		.qe(),
		.q(reg2hw[48]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_16_qs)
	);
	// Trace: design.sv:65721:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_17_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_17_wd),
		.de(hw2reg[98]),
		.d(hw2reg[99]),
		.qe(),
		.q(reg2hw[49]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_17_qs)
	);
	// Trace: design.sv:65747:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_18_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_18_wd),
		.de(hw2reg[100]),
		.d(hw2reg[101]),
		.qe(),
		.q(reg2hw[50]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_18_qs)
	);
	// Trace: design.sv:65773:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_19_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_19_wd),
		.de(hw2reg[102]),
		.d(hw2reg[103]),
		.qe(),
		.q(reg2hw[51]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_19_qs)
	);
	// Trace: design.sv:65799:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_20_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_20_wd),
		.de(hw2reg[104]),
		.d(hw2reg[105]),
		.qe(),
		.q(reg2hw[52]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_20_qs)
	);
	// Trace: design.sv:65825:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_21_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_21_wd),
		.de(hw2reg[106]),
		.d(hw2reg[107]),
		.qe(),
		.q(reg2hw[53]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_21_qs)
	);
	// Trace: design.sv:65851:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_22_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_22_wd),
		.de(hw2reg[108]),
		.d(hw2reg[109]),
		.qe(),
		.q(reg2hw[54]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_22_qs)
	);
	// Trace: design.sv:65877:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_23_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_23_wd),
		.de(hw2reg[110]),
		.d(hw2reg[111]),
		.qe(),
		.q(reg2hw[55]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_23_qs)
	);
	// Trace: design.sv:65903:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_24_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_24_wd),
		.de(hw2reg[112]),
		.d(hw2reg[113]),
		.qe(),
		.q(reg2hw[56]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_24_qs)
	);
	// Trace: design.sv:65929:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_25_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_25_wd),
		.de(hw2reg[114]),
		.d(hw2reg[115]),
		.qe(),
		.q(reg2hw[57]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_25_qs)
	);
	// Trace: design.sv:65955:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_26_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_26_wd),
		.de(hw2reg[116]),
		.d(hw2reg[117]),
		.qe(),
		.q(reg2hw[58]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_26_qs)
	);
	// Trace: design.sv:65981:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_27_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_27_wd),
		.de(hw2reg[118]),
		.d(hw2reg[119]),
		.qe(),
		.q(reg2hw[59]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_27_qs)
	);
	// Trace: design.sv:66007:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_28_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_28_wd),
		.de(hw2reg[120]),
		.d(hw2reg[121]),
		.qe(),
		.q(reg2hw[60]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_28_qs)
	);
	// Trace: design.sv:66033:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_29_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_29_wd),
		.de(hw2reg[122]),
		.d(hw2reg[123]),
		.qe(),
		.q(reg2hw[61]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_29_qs)
	);
	// Trace: design.sv:66059:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_30_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_30_wd),
		.de(hw2reg[124]),
		.d(hw2reg[125]),
		.qe(),
		.q(reg2hw[62]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_30_qs)
	);
	// Trace: design.sv:66085:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_high_status_intrpt_lvl_high_status_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_high_status_intrpt_lvl_high_status_31_we),
		.wd(intrpt_lvl_high_status_intrpt_lvl_high_status_31_wd),
		.de(hw2reg[126]),
		.d(hw2reg[127]),
		.qe(),
		.q(reg2hw[63]),
		.qs(intrpt_lvl_high_status_intrpt_lvl_high_status_31_qs)
	);
	// Trace: design.sv:66116:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_0_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_0_wd),
		.de(hw2reg[0]),
		.d(hw2reg[1]),
		.qe(),
		.q(reg2hw[0]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_0_qs)
	);
	// Trace: design.sv:66142:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_1_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_1_wd),
		.de(hw2reg[2]),
		.d(hw2reg[3]),
		.qe(),
		.q(reg2hw[1]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_1_qs)
	);
	// Trace: design.sv:66168:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_2_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_2_wd),
		.de(hw2reg[4]),
		.d(hw2reg[5]),
		.qe(),
		.q(reg2hw[2]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_2_qs)
	);
	// Trace: design.sv:66194:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_3_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_3_wd),
		.de(hw2reg[6]),
		.d(hw2reg[7]),
		.qe(),
		.q(reg2hw[3]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_3_qs)
	);
	// Trace: design.sv:66220:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_4_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_4_wd),
		.de(hw2reg[8]),
		.d(hw2reg[9]),
		.qe(),
		.q(reg2hw[4]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_4_qs)
	);
	// Trace: design.sv:66246:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_5_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_5_wd),
		.de(hw2reg[10]),
		.d(hw2reg[11]),
		.qe(),
		.q(reg2hw[5]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_5_qs)
	);
	// Trace: design.sv:66272:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_6_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_6_wd),
		.de(hw2reg[12]),
		.d(hw2reg[13]),
		.qe(),
		.q(reg2hw[6]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_6_qs)
	);
	// Trace: design.sv:66298:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_7_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_7_wd),
		.de(hw2reg[14]),
		.d(hw2reg[15]),
		.qe(),
		.q(reg2hw[7]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_7_qs)
	);
	// Trace: design.sv:66324:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_8_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_8_wd),
		.de(hw2reg[16]),
		.d(hw2reg[17]),
		.qe(),
		.q(reg2hw[8]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_8_qs)
	);
	// Trace: design.sv:66350:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_9_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_9_wd),
		.de(hw2reg[18]),
		.d(hw2reg[19]),
		.qe(),
		.q(reg2hw[9]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_9_qs)
	);
	// Trace: design.sv:66376:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_10_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_10_wd),
		.de(hw2reg[20]),
		.d(hw2reg[21]),
		.qe(),
		.q(reg2hw[10]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_10_qs)
	);
	// Trace: design.sv:66402:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_11_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_11_wd),
		.de(hw2reg[22]),
		.d(hw2reg[23]),
		.qe(),
		.q(reg2hw[11]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_11_qs)
	);
	// Trace: design.sv:66428:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_12_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_12_wd),
		.de(hw2reg[24]),
		.d(hw2reg[25]),
		.qe(),
		.q(reg2hw[12]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_12_qs)
	);
	// Trace: design.sv:66454:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_13_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_13_wd),
		.de(hw2reg[26]),
		.d(hw2reg[27]),
		.qe(),
		.q(reg2hw[13]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_13_qs)
	);
	// Trace: design.sv:66480:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_14_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_14_wd),
		.de(hw2reg[28]),
		.d(hw2reg[29]),
		.qe(),
		.q(reg2hw[14]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_14_qs)
	);
	// Trace: design.sv:66506:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_15_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_15_wd),
		.de(hw2reg[30]),
		.d(hw2reg[31]),
		.qe(),
		.q(reg2hw[15]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_15_qs)
	);
	// Trace: design.sv:66532:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_16_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_16_wd),
		.de(hw2reg[32]),
		.d(hw2reg[33]),
		.qe(),
		.q(reg2hw[16]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_16_qs)
	);
	// Trace: design.sv:66558:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_17_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_17_wd),
		.de(hw2reg[34]),
		.d(hw2reg[35]),
		.qe(),
		.q(reg2hw[17]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_17_qs)
	);
	// Trace: design.sv:66584:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_18_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_18_wd),
		.de(hw2reg[36]),
		.d(hw2reg[37]),
		.qe(),
		.q(reg2hw[18]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_18_qs)
	);
	// Trace: design.sv:66610:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_19_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_19_wd),
		.de(hw2reg[38]),
		.d(hw2reg[39]),
		.qe(),
		.q(reg2hw[19]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_19_qs)
	);
	// Trace: design.sv:66636:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_20_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_20_wd),
		.de(hw2reg[40]),
		.d(hw2reg[41]),
		.qe(),
		.q(reg2hw[20]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_20_qs)
	);
	// Trace: design.sv:66662:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_21_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_21_wd),
		.de(hw2reg[42]),
		.d(hw2reg[43]),
		.qe(),
		.q(reg2hw[21]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_21_qs)
	);
	// Trace: design.sv:66688:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_22_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_22_wd),
		.de(hw2reg[44]),
		.d(hw2reg[45]),
		.qe(),
		.q(reg2hw[22]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_22_qs)
	);
	// Trace: design.sv:66714:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_23_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_23_wd),
		.de(hw2reg[46]),
		.d(hw2reg[47]),
		.qe(),
		.q(reg2hw[23]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_23_qs)
	);
	// Trace: design.sv:66740:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_24_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_24_wd),
		.de(hw2reg[48]),
		.d(hw2reg[49]),
		.qe(),
		.q(reg2hw[24]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_24_qs)
	);
	// Trace: design.sv:66766:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_25_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_25_wd),
		.de(hw2reg[50]),
		.d(hw2reg[51]),
		.qe(),
		.q(reg2hw[25]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_25_qs)
	);
	// Trace: design.sv:66792:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_26_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_26_wd),
		.de(hw2reg[52]),
		.d(hw2reg[53]),
		.qe(),
		.q(reg2hw[26]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_26_qs)
	);
	// Trace: design.sv:66818:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_27_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_27_wd),
		.de(hw2reg[54]),
		.d(hw2reg[55]),
		.qe(),
		.q(reg2hw[27]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_27_qs)
	);
	// Trace: design.sv:66844:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_28_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_28_wd),
		.de(hw2reg[56]),
		.d(hw2reg[57]),
		.qe(),
		.q(reg2hw[28]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_28_qs)
	);
	// Trace: design.sv:66870:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_29_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_29_wd),
		.de(hw2reg[58]),
		.d(hw2reg[59]),
		.qe(),
		.q(reg2hw[29]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_29_qs)
	);
	// Trace: design.sv:66896:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_30_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_30_wd),
		.de(hw2reg[60]),
		.d(hw2reg[61]),
		.qe(),
		.q(reg2hw[30]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_30_qs)
	);
	// Trace: design.sv:66922:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intrpt_lvl_low_status_intrpt_lvl_low_status_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intrpt_lvl_low_status_intrpt_lvl_low_status_31_we),
		.wd(intrpt_lvl_low_status_intrpt_lvl_low_status_31_wd),
		.de(hw2reg[62]),
		.d(hw2reg[63]),
		.qe(),
		.q(reg2hw[31]),
		.qs(intrpt_lvl_low_status_intrpt_lvl_low_status_31_qs)
	);
	// Trace: design.sv:66950:3
	reg [18:0] addr_hit;
	// Trace: design.sv:66951:3
	localparam signed [31:0] gpio_reg_pkg_BlockAw = 11;
	localparam [10:0] gpio_reg_pkg_GPIO_CFG_OFFSET = 11'h004;
	localparam [10:0] gpio_reg_pkg_GPIO_GPIO_CLEAR_OFFSET = 11'h280;
	localparam [10:0] gpio_reg_pkg_GPIO_GPIO_EN_OFFSET = 11'h080;
	localparam [10:0] gpio_reg_pkg_GPIO_GPIO_IN_OFFSET = 11'h100;
	localparam [10:0] gpio_reg_pkg_GPIO_GPIO_MODE_0_OFFSET = 11'h008;
	localparam [10:0] gpio_reg_pkg_GPIO_GPIO_MODE_1_OFFSET = 11'h00c;
	localparam [10:0] gpio_reg_pkg_GPIO_GPIO_OUT_OFFSET = 11'h180;
	localparam [10:0] gpio_reg_pkg_GPIO_GPIO_SET_OFFSET = 11'h200;
	localparam [10:0] gpio_reg_pkg_GPIO_GPIO_TOGGLE_OFFSET = 11'h300;
	localparam [10:0] gpio_reg_pkg_GPIO_INFO_OFFSET = 11'h000;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_FALL_EN_OFFSET = 11'h400;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_FALL_STATUS_OFFSET = 11'h680;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_LVL_HIGH_EN_OFFSET = 11'h480;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_LVL_HIGH_STATUS_OFFSET = 11'h700;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_LVL_LOW_EN_OFFSET = 11'h500;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_LVL_LOW_STATUS_OFFSET = 11'h780;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_RISE_EN_OFFSET = 11'h380;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_RISE_STATUS_OFFSET = 11'h600;
	localparam [10:0] gpio_reg_pkg_GPIO_INTRPT_STATUS_OFFSET = 11'h580;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:66952:5
		addr_hit = 1'sb0;
		// Trace: design.sv:66953:5
		addr_hit[0] = reg_addr == gpio_reg_pkg_GPIO_INFO_OFFSET;
		// Trace: design.sv:66954:5
		addr_hit[1] = reg_addr == gpio_reg_pkg_GPIO_CFG_OFFSET;
		// Trace: design.sv:66955:5
		addr_hit[2] = reg_addr == gpio_reg_pkg_GPIO_GPIO_MODE_0_OFFSET;
		// Trace: design.sv:66956:5
		addr_hit[3] = reg_addr == gpio_reg_pkg_GPIO_GPIO_MODE_1_OFFSET;
		// Trace: design.sv:66957:5
		addr_hit[4] = reg_addr == gpio_reg_pkg_GPIO_GPIO_EN_OFFSET;
		// Trace: design.sv:66958:5
		addr_hit[5] = reg_addr == gpio_reg_pkg_GPIO_GPIO_IN_OFFSET;
		// Trace: design.sv:66959:5
		addr_hit[6] = reg_addr == gpio_reg_pkg_GPIO_GPIO_OUT_OFFSET;
		// Trace: design.sv:66960:5
		addr_hit[7] = reg_addr == gpio_reg_pkg_GPIO_GPIO_SET_OFFSET;
		// Trace: design.sv:66961:5
		addr_hit[8] = reg_addr == gpio_reg_pkg_GPIO_GPIO_CLEAR_OFFSET;
		// Trace: design.sv:66962:5
		addr_hit[9] = reg_addr == gpio_reg_pkg_GPIO_GPIO_TOGGLE_OFFSET;
		// Trace: design.sv:66963:5
		addr_hit[10] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_RISE_EN_OFFSET;
		// Trace: design.sv:66964:5
		addr_hit[11] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_FALL_EN_OFFSET;
		// Trace: design.sv:66965:5
		addr_hit[12] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_LVL_HIGH_EN_OFFSET;
		// Trace: design.sv:66966:5
		addr_hit[13] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_LVL_LOW_EN_OFFSET;
		// Trace: design.sv:66967:5
		addr_hit[14] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_STATUS_OFFSET;
		// Trace: design.sv:66968:5
		addr_hit[15] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_RISE_STATUS_OFFSET;
		// Trace: design.sv:66969:5
		addr_hit[16] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_FALL_STATUS_OFFSET;
		// Trace: design.sv:66970:5
		addr_hit[17] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_LVL_HIGH_STATUS_OFFSET;
		// Trace: design.sv:66971:5
		addr_hit[18] = reg_addr == gpio_reg_pkg_GPIO_INTRPT_LVL_LOW_STATUS_OFFSET;
	end
	// Trace: design.sv:66974:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:66977:3
	localparam [75:0] gpio_reg_pkg_GPIO_PERMIT = 76'b0111000111111111111111111111111111111111111111111111111111111111111111111111;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:66978:5
		wr_err = reg_we & (((((((((((((((((((addr_hit[0] & |(gpio_reg_pkg_GPIO_PERMIT[72+:4] & ~reg_be)) | (addr_hit[1] & |(gpio_reg_pkg_GPIO_PERMIT[68+:4] & ~reg_be))) | (addr_hit[2] & |(gpio_reg_pkg_GPIO_PERMIT[64+:4] & ~reg_be))) | (addr_hit[3] & |(gpio_reg_pkg_GPIO_PERMIT[60+:4] & ~reg_be))) | (addr_hit[4] & |(gpio_reg_pkg_GPIO_PERMIT[56+:4] & ~reg_be))) | (addr_hit[5] & |(gpio_reg_pkg_GPIO_PERMIT[52+:4] & ~reg_be))) | (addr_hit[6] & |(gpio_reg_pkg_GPIO_PERMIT[48+:4] & ~reg_be))) | (addr_hit[7] & |(gpio_reg_pkg_GPIO_PERMIT[44+:4] & ~reg_be))) | (addr_hit[8] & |(gpio_reg_pkg_GPIO_PERMIT[40+:4] & ~reg_be))) | (addr_hit[9] & |(gpio_reg_pkg_GPIO_PERMIT[36+:4] & ~reg_be))) | (addr_hit[10] & |(gpio_reg_pkg_GPIO_PERMIT[32+:4] & ~reg_be))) | (addr_hit[11] & |(gpio_reg_pkg_GPIO_PERMIT[28+:4] & ~reg_be))) | (addr_hit[12] & |(gpio_reg_pkg_GPIO_PERMIT[24+:4] & ~reg_be))) | (addr_hit[13] & |(gpio_reg_pkg_GPIO_PERMIT[20+:4] & ~reg_be))) | (addr_hit[14] & |(gpio_reg_pkg_GPIO_PERMIT[16+:4] & ~reg_be))) | (addr_hit[15] & |(gpio_reg_pkg_GPIO_PERMIT[12+:4] & ~reg_be))) | (addr_hit[16] & |(gpio_reg_pkg_GPIO_PERMIT[8+:4] & ~reg_be))) | (addr_hit[17] & |(gpio_reg_pkg_GPIO_PERMIT[4+:4] & ~reg_be))) | (addr_hit[18] & |(gpio_reg_pkg_GPIO_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:67000:3
	assign info_gpio_cnt_re = (addr_hit[0] & reg_re) & !reg_error;
	// Trace: design.sv:67002:3
	assign info_version_re = (addr_hit[0] & reg_re) & !reg_error;
	// Trace: design.sv:67004:3
	assign cfg_glbl_intrpt_mode_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:67005:3
	assign cfg_glbl_intrpt_mode_wd = reg_wdata[0];
	// Trace: design.sv:67007:3
	assign cfg_pin_lvl_intrpt_mode_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:67008:3
	assign cfg_pin_lvl_intrpt_mode_wd = reg_wdata[0];
	// Trace: design.sv:67010:3
	assign cfg_reserved_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:67011:3
	assign cfg_reserved_wd = reg_wdata[1];
	// Trace: design.sv:67013:3
	assign gpio_mode_0_mode_0_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67014:3
	assign gpio_mode_0_mode_0_wd = reg_wdata[1:0];
	// Trace: design.sv:67016:3
	assign gpio_mode_0_mode_1_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67017:3
	assign gpio_mode_0_mode_1_wd = reg_wdata[3:2];
	// Trace: design.sv:67019:3
	assign gpio_mode_0_mode_2_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67020:3
	assign gpio_mode_0_mode_2_wd = reg_wdata[5:4];
	// Trace: design.sv:67022:3
	assign gpio_mode_0_mode_3_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67023:3
	assign gpio_mode_0_mode_3_wd = reg_wdata[7:6];
	// Trace: design.sv:67025:3
	assign gpio_mode_0_mode_4_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67026:3
	assign gpio_mode_0_mode_4_wd = reg_wdata[9:8];
	// Trace: design.sv:67028:3
	assign gpio_mode_0_mode_5_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67029:3
	assign gpio_mode_0_mode_5_wd = reg_wdata[11:10];
	// Trace: design.sv:67031:3
	assign gpio_mode_0_mode_6_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67032:3
	assign gpio_mode_0_mode_6_wd = reg_wdata[13:12];
	// Trace: design.sv:67034:3
	assign gpio_mode_0_mode_7_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67035:3
	assign gpio_mode_0_mode_7_wd = reg_wdata[15:14];
	// Trace: design.sv:67037:3
	assign gpio_mode_0_mode_8_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67038:3
	assign gpio_mode_0_mode_8_wd = reg_wdata[17:16];
	// Trace: design.sv:67040:3
	assign gpio_mode_0_mode_9_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67041:3
	assign gpio_mode_0_mode_9_wd = reg_wdata[19:18];
	// Trace: design.sv:67043:3
	assign gpio_mode_0_mode_10_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67044:3
	assign gpio_mode_0_mode_10_wd = reg_wdata[21:20];
	// Trace: design.sv:67046:3
	assign gpio_mode_0_mode_11_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67047:3
	assign gpio_mode_0_mode_11_wd = reg_wdata[23:22];
	// Trace: design.sv:67049:3
	assign gpio_mode_0_mode_12_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67050:3
	assign gpio_mode_0_mode_12_wd = reg_wdata[25:24];
	// Trace: design.sv:67052:3
	assign gpio_mode_0_mode_13_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67053:3
	assign gpio_mode_0_mode_13_wd = reg_wdata[27:26];
	// Trace: design.sv:67055:3
	assign gpio_mode_0_mode_14_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67056:3
	assign gpio_mode_0_mode_14_wd = reg_wdata[29:28];
	// Trace: design.sv:67058:3
	assign gpio_mode_0_mode_15_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:67059:3
	assign gpio_mode_0_mode_15_wd = reg_wdata[31:30];
	// Trace: design.sv:67061:3
	assign gpio_mode_1_mode_16_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67062:3
	assign gpio_mode_1_mode_16_wd = reg_wdata[1:0];
	// Trace: design.sv:67064:3
	assign gpio_mode_1_mode_17_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67065:3
	assign gpio_mode_1_mode_17_wd = reg_wdata[3:2];
	// Trace: design.sv:67067:3
	assign gpio_mode_1_mode_18_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67068:3
	assign gpio_mode_1_mode_18_wd = reg_wdata[5:4];
	// Trace: design.sv:67070:3
	assign gpio_mode_1_mode_19_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67071:3
	assign gpio_mode_1_mode_19_wd = reg_wdata[7:6];
	// Trace: design.sv:67073:3
	assign gpio_mode_1_mode_20_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67074:3
	assign gpio_mode_1_mode_20_wd = reg_wdata[9:8];
	// Trace: design.sv:67076:3
	assign gpio_mode_1_mode_21_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67077:3
	assign gpio_mode_1_mode_21_wd = reg_wdata[11:10];
	// Trace: design.sv:67079:3
	assign gpio_mode_1_mode_22_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67080:3
	assign gpio_mode_1_mode_22_wd = reg_wdata[13:12];
	// Trace: design.sv:67082:3
	assign gpio_mode_1_mode_23_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67083:3
	assign gpio_mode_1_mode_23_wd = reg_wdata[15:14];
	// Trace: design.sv:67085:3
	assign gpio_mode_1_mode_24_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67086:3
	assign gpio_mode_1_mode_24_wd = reg_wdata[17:16];
	// Trace: design.sv:67088:3
	assign gpio_mode_1_mode_25_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67089:3
	assign gpio_mode_1_mode_25_wd = reg_wdata[19:18];
	// Trace: design.sv:67091:3
	assign gpio_mode_1_mode_26_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67092:3
	assign gpio_mode_1_mode_26_wd = reg_wdata[21:20];
	// Trace: design.sv:67094:3
	assign gpio_mode_1_mode_27_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67095:3
	assign gpio_mode_1_mode_27_wd = reg_wdata[23:22];
	// Trace: design.sv:67097:3
	assign gpio_mode_1_mode_28_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67098:3
	assign gpio_mode_1_mode_28_wd = reg_wdata[25:24];
	// Trace: design.sv:67100:3
	assign gpio_mode_1_mode_29_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67101:3
	assign gpio_mode_1_mode_29_wd = reg_wdata[27:26];
	// Trace: design.sv:67103:3
	assign gpio_mode_1_mode_30_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67104:3
	assign gpio_mode_1_mode_30_wd = reg_wdata[29:28];
	// Trace: design.sv:67106:3
	assign gpio_mode_1_mode_31_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:67107:3
	assign gpio_mode_1_mode_31_wd = reg_wdata[31:30];
	// Trace: design.sv:67109:3
	assign gpio_en_gpio_en_0_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67110:3
	assign gpio_en_gpio_en_0_wd = reg_wdata[0];
	// Trace: design.sv:67112:3
	assign gpio_en_gpio_en_1_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67113:3
	assign gpio_en_gpio_en_1_wd = reg_wdata[1];
	// Trace: design.sv:67115:3
	assign gpio_en_gpio_en_2_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67116:3
	assign gpio_en_gpio_en_2_wd = reg_wdata[2];
	// Trace: design.sv:67118:3
	assign gpio_en_gpio_en_3_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67119:3
	assign gpio_en_gpio_en_3_wd = reg_wdata[3];
	// Trace: design.sv:67121:3
	assign gpio_en_gpio_en_4_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67122:3
	assign gpio_en_gpio_en_4_wd = reg_wdata[4];
	// Trace: design.sv:67124:3
	assign gpio_en_gpio_en_5_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67125:3
	assign gpio_en_gpio_en_5_wd = reg_wdata[5];
	// Trace: design.sv:67127:3
	assign gpio_en_gpio_en_6_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67128:3
	assign gpio_en_gpio_en_6_wd = reg_wdata[6];
	// Trace: design.sv:67130:3
	assign gpio_en_gpio_en_7_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67131:3
	assign gpio_en_gpio_en_7_wd = reg_wdata[7];
	// Trace: design.sv:67133:3
	assign gpio_en_gpio_en_8_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67134:3
	assign gpio_en_gpio_en_8_wd = reg_wdata[8];
	// Trace: design.sv:67136:3
	assign gpio_en_gpio_en_9_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67137:3
	assign gpio_en_gpio_en_9_wd = reg_wdata[9];
	// Trace: design.sv:67139:3
	assign gpio_en_gpio_en_10_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67140:3
	assign gpio_en_gpio_en_10_wd = reg_wdata[10];
	// Trace: design.sv:67142:3
	assign gpio_en_gpio_en_11_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67143:3
	assign gpio_en_gpio_en_11_wd = reg_wdata[11];
	// Trace: design.sv:67145:3
	assign gpio_en_gpio_en_12_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67146:3
	assign gpio_en_gpio_en_12_wd = reg_wdata[12];
	// Trace: design.sv:67148:3
	assign gpio_en_gpio_en_13_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67149:3
	assign gpio_en_gpio_en_13_wd = reg_wdata[13];
	// Trace: design.sv:67151:3
	assign gpio_en_gpio_en_14_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67152:3
	assign gpio_en_gpio_en_14_wd = reg_wdata[14];
	// Trace: design.sv:67154:3
	assign gpio_en_gpio_en_15_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67155:3
	assign gpio_en_gpio_en_15_wd = reg_wdata[15];
	// Trace: design.sv:67157:3
	assign gpio_en_gpio_en_16_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67158:3
	assign gpio_en_gpio_en_16_wd = reg_wdata[16];
	// Trace: design.sv:67160:3
	assign gpio_en_gpio_en_17_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67161:3
	assign gpio_en_gpio_en_17_wd = reg_wdata[17];
	// Trace: design.sv:67163:3
	assign gpio_en_gpio_en_18_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67164:3
	assign gpio_en_gpio_en_18_wd = reg_wdata[18];
	// Trace: design.sv:67166:3
	assign gpio_en_gpio_en_19_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67167:3
	assign gpio_en_gpio_en_19_wd = reg_wdata[19];
	// Trace: design.sv:67169:3
	assign gpio_en_gpio_en_20_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67170:3
	assign gpio_en_gpio_en_20_wd = reg_wdata[20];
	// Trace: design.sv:67172:3
	assign gpio_en_gpio_en_21_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67173:3
	assign gpio_en_gpio_en_21_wd = reg_wdata[21];
	// Trace: design.sv:67175:3
	assign gpio_en_gpio_en_22_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67176:3
	assign gpio_en_gpio_en_22_wd = reg_wdata[22];
	// Trace: design.sv:67178:3
	assign gpio_en_gpio_en_23_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67179:3
	assign gpio_en_gpio_en_23_wd = reg_wdata[23];
	// Trace: design.sv:67181:3
	assign gpio_en_gpio_en_24_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67182:3
	assign gpio_en_gpio_en_24_wd = reg_wdata[24];
	// Trace: design.sv:67184:3
	assign gpio_en_gpio_en_25_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67185:3
	assign gpio_en_gpio_en_25_wd = reg_wdata[25];
	// Trace: design.sv:67187:3
	assign gpio_en_gpio_en_26_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67188:3
	assign gpio_en_gpio_en_26_wd = reg_wdata[26];
	// Trace: design.sv:67190:3
	assign gpio_en_gpio_en_27_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67191:3
	assign gpio_en_gpio_en_27_wd = reg_wdata[27];
	// Trace: design.sv:67193:3
	assign gpio_en_gpio_en_28_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67194:3
	assign gpio_en_gpio_en_28_wd = reg_wdata[28];
	// Trace: design.sv:67196:3
	assign gpio_en_gpio_en_29_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67197:3
	assign gpio_en_gpio_en_29_wd = reg_wdata[29];
	// Trace: design.sv:67199:3
	assign gpio_en_gpio_en_30_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67200:3
	assign gpio_en_gpio_en_30_wd = reg_wdata[30];
	// Trace: design.sv:67202:3
	assign gpio_en_gpio_en_31_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:67203:3
	assign gpio_en_gpio_en_31_wd = reg_wdata[31];
	// Trace: design.sv:67205:3
	assign gpio_in_gpio_in_0_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67207:3
	assign gpio_in_gpio_in_1_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67209:3
	assign gpio_in_gpio_in_2_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67211:3
	assign gpio_in_gpio_in_3_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67213:3
	assign gpio_in_gpio_in_4_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67215:3
	assign gpio_in_gpio_in_5_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67217:3
	assign gpio_in_gpio_in_6_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67219:3
	assign gpio_in_gpio_in_7_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67221:3
	assign gpio_in_gpio_in_8_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67223:3
	assign gpio_in_gpio_in_9_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67225:3
	assign gpio_in_gpio_in_10_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67227:3
	assign gpio_in_gpio_in_11_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67229:3
	assign gpio_in_gpio_in_12_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67231:3
	assign gpio_in_gpio_in_13_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67233:3
	assign gpio_in_gpio_in_14_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67235:3
	assign gpio_in_gpio_in_15_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67237:3
	assign gpio_in_gpio_in_16_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67239:3
	assign gpio_in_gpio_in_17_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67241:3
	assign gpio_in_gpio_in_18_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67243:3
	assign gpio_in_gpio_in_19_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67245:3
	assign gpio_in_gpio_in_20_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67247:3
	assign gpio_in_gpio_in_21_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67249:3
	assign gpio_in_gpio_in_22_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67251:3
	assign gpio_in_gpio_in_23_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67253:3
	assign gpio_in_gpio_in_24_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67255:3
	assign gpio_in_gpio_in_25_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67257:3
	assign gpio_in_gpio_in_26_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67259:3
	assign gpio_in_gpio_in_27_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67261:3
	assign gpio_in_gpio_in_28_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67263:3
	assign gpio_in_gpio_in_29_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67265:3
	assign gpio_in_gpio_in_30_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67267:3
	assign gpio_in_gpio_in_31_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:67269:3
	assign gpio_out_gpio_out_0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67270:3
	assign gpio_out_gpio_out_0_wd = reg_wdata[0];
	// Trace: design.sv:67272:3
	assign gpio_out_gpio_out_1_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67273:3
	assign gpio_out_gpio_out_1_wd = reg_wdata[1];
	// Trace: design.sv:67275:3
	assign gpio_out_gpio_out_2_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67276:3
	assign gpio_out_gpio_out_2_wd = reg_wdata[2];
	// Trace: design.sv:67278:3
	assign gpio_out_gpio_out_3_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67279:3
	assign gpio_out_gpio_out_3_wd = reg_wdata[3];
	// Trace: design.sv:67281:3
	assign gpio_out_gpio_out_4_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67282:3
	assign gpio_out_gpio_out_4_wd = reg_wdata[4];
	// Trace: design.sv:67284:3
	assign gpio_out_gpio_out_5_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67285:3
	assign gpio_out_gpio_out_5_wd = reg_wdata[5];
	// Trace: design.sv:67287:3
	assign gpio_out_gpio_out_6_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67288:3
	assign gpio_out_gpio_out_6_wd = reg_wdata[6];
	// Trace: design.sv:67290:3
	assign gpio_out_gpio_out_7_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67291:3
	assign gpio_out_gpio_out_7_wd = reg_wdata[7];
	// Trace: design.sv:67293:3
	assign gpio_out_gpio_out_8_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67294:3
	assign gpio_out_gpio_out_8_wd = reg_wdata[8];
	// Trace: design.sv:67296:3
	assign gpio_out_gpio_out_9_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67297:3
	assign gpio_out_gpio_out_9_wd = reg_wdata[9];
	// Trace: design.sv:67299:3
	assign gpio_out_gpio_out_10_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67300:3
	assign gpio_out_gpio_out_10_wd = reg_wdata[10];
	// Trace: design.sv:67302:3
	assign gpio_out_gpio_out_11_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67303:3
	assign gpio_out_gpio_out_11_wd = reg_wdata[11];
	// Trace: design.sv:67305:3
	assign gpio_out_gpio_out_12_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67306:3
	assign gpio_out_gpio_out_12_wd = reg_wdata[12];
	// Trace: design.sv:67308:3
	assign gpio_out_gpio_out_13_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67309:3
	assign gpio_out_gpio_out_13_wd = reg_wdata[13];
	// Trace: design.sv:67311:3
	assign gpio_out_gpio_out_14_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67312:3
	assign gpio_out_gpio_out_14_wd = reg_wdata[14];
	// Trace: design.sv:67314:3
	assign gpio_out_gpio_out_15_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67315:3
	assign gpio_out_gpio_out_15_wd = reg_wdata[15];
	// Trace: design.sv:67317:3
	assign gpio_out_gpio_out_16_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67318:3
	assign gpio_out_gpio_out_16_wd = reg_wdata[16];
	// Trace: design.sv:67320:3
	assign gpio_out_gpio_out_17_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67321:3
	assign gpio_out_gpio_out_17_wd = reg_wdata[17];
	// Trace: design.sv:67323:3
	assign gpio_out_gpio_out_18_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67324:3
	assign gpio_out_gpio_out_18_wd = reg_wdata[18];
	// Trace: design.sv:67326:3
	assign gpio_out_gpio_out_19_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67327:3
	assign gpio_out_gpio_out_19_wd = reg_wdata[19];
	// Trace: design.sv:67329:3
	assign gpio_out_gpio_out_20_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67330:3
	assign gpio_out_gpio_out_20_wd = reg_wdata[20];
	// Trace: design.sv:67332:3
	assign gpio_out_gpio_out_21_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67333:3
	assign gpio_out_gpio_out_21_wd = reg_wdata[21];
	// Trace: design.sv:67335:3
	assign gpio_out_gpio_out_22_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67336:3
	assign gpio_out_gpio_out_22_wd = reg_wdata[22];
	// Trace: design.sv:67338:3
	assign gpio_out_gpio_out_23_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67339:3
	assign gpio_out_gpio_out_23_wd = reg_wdata[23];
	// Trace: design.sv:67341:3
	assign gpio_out_gpio_out_24_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67342:3
	assign gpio_out_gpio_out_24_wd = reg_wdata[24];
	// Trace: design.sv:67344:3
	assign gpio_out_gpio_out_25_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67345:3
	assign gpio_out_gpio_out_25_wd = reg_wdata[25];
	// Trace: design.sv:67347:3
	assign gpio_out_gpio_out_26_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67348:3
	assign gpio_out_gpio_out_26_wd = reg_wdata[26];
	// Trace: design.sv:67350:3
	assign gpio_out_gpio_out_27_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67351:3
	assign gpio_out_gpio_out_27_wd = reg_wdata[27];
	// Trace: design.sv:67353:3
	assign gpio_out_gpio_out_28_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67354:3
	assign gpio_out_gpio_out_28_wd = reg_wdata[28];
	// Trace: design.sv:67356:3
	assign gpio_out_gpio_out_29_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67357:3
	assign gpio_out_gpio_out_29_wd = reg_wdata[29];
	// Trace: design.sv:67359:3
	assign gpio_out_gpio_out_30_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67360:3
	assign gpio_out_gpio_out_30_wd = reg_wdata[30];
	// Trace: design.sv:67362:3
	assign gpio_out_gpio_out_31_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:67363:3
	assign gpio_out_gpio_out_31_wd = reg_wdata[31];
	// Trace: design.sv:67365:3
	assign gpio_set_gpio_set_0_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67366:3
	assign gpio_set_gpio_set_0_wd = reg_wdata[0];
	// Trace: design.sv:67368:3
	assign gpio_set_gpio_set_1_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67369:3
	assign gpio_set_gpio_set_1_wd = reg_wdata[1];
	// Trace: design.sv:67371:3
	assign gpio_set_gpio_set_2_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67372:3
	assign gpio_set_gpio_set_2_wd = reg_wdata[2];
	// Trace: design.sv:67374:3
	assign gpio_set_gpio_set_3_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67375:3
	assign gpio_set_gpio_set_3_wd = reg_wdata[3];
	// Trace: design.sv:67377:3
	assign gpio_set_gpio_set_4_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67378:3
	assign gpio_set_gpio_set_4_wd = reg_wdata[4];
	// Trace: design.sv:67380:3
	assign gpio_set_gpio_set_5_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67381:3
	assign gpio_set_gpio_set_5_wd = reg_wdata[5];
	// Trace: design.sv:67383:3
	assign gpio_set_gpio_set_6_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67384:3
	assign gpio_set_gpio_set_6_wd = reg_wdata[6];
	// Trace: design.sv:67386:3
	assign gpio_set_gpio_set_7_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67387:3
	assign gpio_set_gpio_set_7_wd = reg_wdata[7];
	// Trace: design.sv:67389:3
	assign gpio_set_gpio_set_8_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67390:3
	assign gpio_set_gpio_set_8_wd = reg_wdata[8];
	// Trace: design.sv:67392:3
	assign gpio_set_gpio_set_9_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67393:3
	assign gpio_set_gpio_set_9_wd = reg_wdata[9];
	// Trace: design.sv:67395:3
	assign gpio_set_gpio_set_10_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67396:3
	assign gpio_set_gpio_set_10_wd = reg_wdata[10];
	// Trace: design.sv:67398:3
	assign gpio_set_gpio_set_11_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67399:3
	assign gpio_set_gpio_set_11_wd = reg_wdata[11];
	// Trace: design.sv:67401:3
	assign gpio_set_gpio_set_12_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67402:3
	assign gpio_set_gpio_set_12_wd = reg_wdata[12];
	// Trace: design.sv:67404:3
	assign gpio_set_gpio_set_13_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67405:3
	assign gpio_set_gpio_set_13_wd = reg_wdata[13];
	// Trace: design.sv:67407:3
	assign gpio_set_gpio_set_14_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67408:3
	assign gpio_set_gpio_set_14_wd = reg_wdata[14];
	// Trace: design.sv:67410:3
	assign gpio_set_gpio_set_15_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67411:3
	assign gpio_set_gpio_set_15_wd = reg_wdata[15];
	// Trace: design.sv:67413:3
	assign gpio_set_gpio_set_16_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67414:3
	assign gpio_set_gpio_set_16_wd = reg_wdata[16];
	// Trace: design.sv:67416:3
	assign gpio_set_gpio_set_17_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67417:3
	assign gpio_set_gpio_set_17_wd = reg_wdata[17];
	// Trace: design.sv:67419:3
	assign gpio_set_gpio_set_18_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67420:3
	assign gpio_set_gpio_set_18_wd = reg_wdata[18];
	// Trace: design.sv:67422:3
	assign gpio_set_gpio_set_19_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67423:3
	assign gpio_set_gpio_set_19_wd = reg_wdata[19];
	// Trace: design.sv:67425:3
	assign gpio_set_gpio_set_20_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67426:3
	assign gpio_set_gpio_set_20_wd = reg_wdata[20];
	// Trace: design.sv:67428:3
	assign gpio_set_gpio_set_21_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67429:3
	assign gpio_set_gpio_set_21_wd = reg_wdata[21];
	// Trace: design.sv:67431:3
	assign gpio_set_gpio_set_22_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67432:3
	assign gpio_set_gpio_set_22_wd = reg_wdata[22];
	// Trace: design.sv:67434:3
	assign gpio_set_gpio_set_23_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67435:3
	assign gpio_set_gpio_set_23_wd = reg_wdata[23];
	// Trace: design.sv:67437:3
	assign gpio_set_gpio_set_24_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67438:3
	assign gpio_set_gpio_set_24_wd = reg_wdata[24];
	// Trace: design.sv:67440:3
	assign gpio_set_gpio_set_25_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67441:3
	assign gpio_set_gpio_set_25_wd = reg_wdata[25];
	// Trace: design.sv:67443:3
	assign gpio_set_gpio_set_26_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67444:3
	assign gpio_set_gpio_set_26_wd = reg_wdata[26];
	// Trace: design.sv:67446:3
	assign gpio_set_gpio_set_27_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67447:3
	assign gpio_set_gpio_set_27_wd = reg_wdata[27];
	// Trace: design.sv:67449:3
	assign gpio_set_gpio_set_28_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67450:3
	assign gpio_set_gpio_set_28_wd = reg_wdata[28];
	// Trace: design.sv:67452:3
	assign gpio_set_gpio_set_29_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67453:3
	assign gpio_set_gpio_set_29_wd = reg_wdata[29];
	// Trace: design.sv:67455:3
	assign gpio_set_gpio_set_30_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67456:3
	assign gpio_set_gpio_set_30_wd = reg_wdata[30];
	// Trace: design.sv:67458:3
	assign gpio_set_gpio_set_31_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:67459:3
	assign gpio_set_gpio_set_31_wd = reg_wdata[31];
	// Trace: design.sv:67461:3
	assign gpio_clear_gpio_clear_0_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67462:3
	assign gpio_clear_gpio_clear_0_wd = reg_wdata[0];
	// Trace: design.sv:67464:3
	assign gpio_clear_gpio_clear_1_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67465:3
	assign gpio_clear_gpio_clear_1_wd = reg_wdata[1];
	// Trace: design.sv:67467:3
	assign gpio_clear_gpio_clear_2_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67468:3
	assign gpio_clear_gpio_clear_2_wd = reg_wdata[2];
	// Trace: design.sv:67470:3
	assign gpio_clear_gpio_clear_3_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67471:3
	assign gpio_clear_gpio_clear_3_wd = reg_wdata[3];
	// Trace: design.sv:67473:3
	assign gpio_clear_gpio_clear_4_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67474:3
	assign gpio_clear_gpio_clear_4_wd = reg_wdata[4];
	// Trace: design.sv:67476:3
	assign gpio_clear_gpio_clear_5_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67477:3
	assign gpio_clear_gpio_clear_5_wd = reg_wdata[5];
	// Trace: design.sv:67479:3
	assign gpio_clear_gpio_clear_6_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67480:3
	assign gpio_clear_gpio_clear_6_wd = reg_wdata[6];
	// Trace: design.sv:67482:3
	assign gpio_clear_gpio_clear_7_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67483:3
	assign gpio_clear_gpio_clear_7_wd = reg_wdata[7];
	// Trace: design.sv:67485:3
	assign gpio_clear_gpio_clear_8_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67486:3
	assign gpio_clear_gpio_clear_8_wd = reg_wdata[8];
	// Trace: design.sv:67488:3
	assign gpio_clear_gpio_clear_9_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67489:3
	assign gpio_clear_gpio_clear_9_wd = reg_wdata[9];
	// Trace: design.sv:67491:3
	assign gpio_clear_gpio_clear_10_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67492:3
	assign gpio_clear_gpio_clear_10_wd = reg_wdata[10];
	// Trace: design.sv:67494:3
	assign gpio_clear_gpio_clear_11_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67495:3
	assign gpio_clear_gpio_clear_11_wd = reg_wdata[11];
	// Trace: design.sv:67497:3
	assign gpio_clear_gpio_clear_12_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67498:3
	assign gpio_clear_gpio_clear_12_wd = reg_wdata[12];
	// Trace: design.sv:67500:3
	assign gpio_clear_gpio_clear_13_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67501:3
	assign gpio_clear_gpio_clear_13_wd = reg_wdata[13];
	// Trace: design.sv:67503:3
	assign gpio_clear_gpio_clear_14_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67504:3
	assign gpio_clear_gpio_clear_14_wd = reg_wdata[14];
	// Trace: design.sv:67506:3
	assign gpio_clear_gpio_clear_15_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67507:3
	assign gpio_clear_gpio_clear_15_wd = reg_wdata[15];
	// Trace: design.sv:67509:3
	assign gpio_clear_gpio_clear_16_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67510:3
	assign gpio_clear_gpio_clear_16_wd = reg_wdata[16];
	// Trace: design.sv:67512:3
	assign gpio_clear_gpio_clear_17_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67513:3
	assign gpio_clear_gpio_clear_17_wd = reg_wdata[17];
	// Trace: design.sv:67515:3
	assign gpio_clear_gpio_clear_18_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67516:3
	assign gpio_clear_gpio_clear_18_wd = reg_wdata[18];
	// Trace: design.sv:67518:3
	assign gpio_clear_gpio_clear_19_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67519:3
	assign gpio_clear_gpio_clear_19_wd = reg_wdata[19];
	// Trace: design.sv:67521:3
	assign gpio_clear_gpio_clear_20_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67522:3
	assign gpio_clear_gpio_clear_20_wd = reg_wdata[20];
	// Trace: design.sv:67524:3
	assign gpio_clear_gpio_clear_21_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67525:3
	assign gpio_clear_gpio_clear_21_wd = reg_wdata[21];
	// Trace: design.sv:67527:3
	assign gpio_clear_gpio_clear_22_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67528:3
	assign gpio_clear_gpio_clear_22_wd = reg_wdata[22];
	// Trace: design.sv:67530:3
	assign gpio_clear_gpio_clear_23_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67531:3
	assign gpio_clear_gpio_clear_23_wd = reg_wdata[23];
	// Trace: design.sv:67533:3
	assign gpio_clear_gpio_clear_24_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67534:3
	assign gpio_clear_gpio_clear_24_wd = reg_wdata[24];
	// Trace: design.sv:67536:3
	assign gpio_clear_gpio_clear_25_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67537:3
	assign gpio_clear_gpio_clear_25_wd = reg_wdata[25];
	// Trace: design.sv:67539:3
	assign gpio_clear_gpio_clear_26_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67540:3
	assign gpio_clear_gpio_clear_26_wd = reg_wdata[26];
	// Trace: design.sv:67542:3
	assign gpio_clear_gpio_clear_27_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67543:3
	assign gpio_clear_gpio_clear_27_wd = reg_wdata[27];
	// Trace: design.sv:67545:3
	assign gpio_clear_gpio_clear_28_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67546:3
	assign gpio_clear_gpio_clear_28_wd = reg_wdata[28];
	// Trace: design.sv:67548:3
	assign gpio_clear_gpio_clear_29_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67549:3
	assign gpio_clear_gpio_clear_29_wd = reg_wdata[29];
	// Trace: design.sv:67551:3
	assign gpio_clear_gpio_clear_30_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67552:3
	assign gpio_clear_gpio_clear_30_wd = reg_wdata[30];
	// Trace: design.sv:67554:3
	assign gpio_clear_gpio_clear_31_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:67555:3
	assign gpio_clear_gpio_clear_31_wd = reg_wdata[31];
	// Trace: design.sv:67557:3
	assign gpio_toggle_gpio_toggle_0_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67558:3
	assign gpio_toggle_gpio_toggle_0_wd = reg_wdata[0];
	// Trace: design.sv:67560:3
	assign gpio_toggle_gpio_toggle_1_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67561:3
	assign gpio_toggle_gpio_toggle_1_wd = reg_wdata[1];
	// Trace: design.sv:67563:3
	assign gpio_toggle_gpio_toggle_2_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67564:3
	assign gpio_toggle_gpio_toggle_2_wd = reg_wdata[2];
	// Trace: design.sv:67566:3
	assign gpio_toggle_gpio_toggle_3_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67567:3
	assign gpio_toggle_gpio_toggle_3_wd = reg_wdata[3];
	// Trace: design.sv:67569:3
	assign gpio_toggle_gpio_toggle_4_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67570:3
	assign gpio_toggle_gpio_toggle_4_wd = reg_wdata[4];
	// Trace: design.sv:67572:3
	assign gpio_toggle_gpio_toggle_5_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67573:3
	assign gpio_toggle_gpio_toggle_5_wd = reg_wdata[5];
	// Trace: design.sv:67575:3
	assign gpio_toggle_gpio_toggle_6_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67576:3
	assign gpio_toggle_gpio_toggle_6_wd = reg_wdata[6];
	// Trace: design.sv:67578:3
	assign gpio_toggle_gpio_toggle_7_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67579:3
	assign gpio_toggle_gpio_toggle_7_wd = reg_wdata[7];
	// Trace: design.sv:67581:3
	assign gpio_toggle_gpio_toggle_8_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67582:3
	assign gpio_toggle_gpio_toggle_8_wd = reg_wdata[8];
	// Trace: design.sv:67584:3
	assign gpio_toggle_gpio_toggle_9_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67585:3
	assign gpio_toggle_gpio_toggle_9_wd = reg_wdata[9];
	// Trace: design.sv:67587:3
	assign gpio_toggle_gpio_toggle_10_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67588:3
	assign gpio_toggle_gpio_toggle_10_wd = reg_wdata[10];
	// Trace: design.sv:67590:3
	assign gpio_toggle_gpio_toggle_11_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67591:3
	assign gpio_toggle_gpio_toggle_11_wd = reg_wdata[11];
	// Trace: design.sv:67593:3
	assign gpio_toggle_gpio_toggle_12_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67594:3
	assign gpio_toggle_gpio_toggle_12_wd = reg_wdata[12];
	// Trace: design.sv:67596:3
	assign gpio_toggle_gpio_toggle_13_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67597:3
	assign gpio_toggle_gpio_toggle_13_wd = reg_wdata[13];
	// Trace: design.sv:67599:3
	assign gpio_toggle_gpio_toggle_14_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67600:3
	assign gpio_toggle_gpio_toggle_14_wd = reg_wdata[14];
	// Trace: design.sv:67602:3
	assign gpio_toggle_gpio_toggle_15_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67603:3
	assign gpio_toggle_gpio_toggle_15_wd = reg_wdata[15];
	// Trace: design.sv:67605:3
	assign gpio_toggle_gpio_toggle_16_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67606:3
	assign gpio_toggle_gpio_toggle_16_wd = reg_wdata[16];
	// Trace: design.sv:67608:3
	assign gpio_toggle_gpio_toggle_17_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67609:3
	assign gpio_toggle_gpio_toggle_17_wd = reg_wdata[17];
	// Trace: design.sv:67611:3
	assign gpio_toggle_gpio_toggle_18_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67612:3
	assign gpio_toggle_gpio_toggle_18_wd = reg_wdata[18];
	// Trace: design.sv:67614:3
	assign gpio_toggle_gpio_toggle_19_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67615:3
	assign gpio_toggle_gpio_toggle_19_wd = reg_wdata[19];
	// Trace: design.sv:67617:3
	assign gpio_toggle_gpio_toggle_20_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67618:3
	assign gpio_toggle_gpio_toggle_20_wd = reg_wdata[20];
	// Trace: design.sv:67620:3
	assign gpio_toggle_gpio_toggle_21_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67621:3
	assign gpio_toggle_gpio_toggle_21_wd = reg_wdata[21];
	// Trace: design.sv:67623:3
	assign gpio_toggle_gpio_toggle_22_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67624:3
	assign gpio_toggle_gpio_toggle_22_wd = reg_wdata[22];
	// Trace: design.sv:67626:3
	assign gpio_toggle_gpio_toggle_23_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67627:3
	assign gpio_toggle_gpio_toggle_23_wd = reg_wdata[23];
	// Trace: design.sv:67629:3
	assign gpio_toggle_gpio_toggle_24_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67630:3
	assign gpio_toggle_gpio_toggle_24_wd = reg_wdata[24];
	// Trace: design.sv:67632:3
	assign gpio_toggle_gpio_toggle_25_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67633:3
	assign gpio_toggle_gpio_toggle_25_wd = reg_wdata[25];
	// Trace: design.sv:67635:3
	assign gpio_toggle_gpio_toggle_26_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67636:3
	assign gpio_toggle_gpio_toggle_26_wd = reg_wdata[26];
	// Trace: design.sv:67638:3
	assign gpio_toggle_gpio_toggle_27_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67639:3
	assign gpio_toggle_gpio_toggle_27_wd = reg_wdata[27];
	// Trace: design.sv:67641:3
	assign gpio_toggle_gpio_toggle_28_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67642:3
	assign gpio_toggle_gpio_toggle_28_wd = reg_wdata[28];
	// Trace: design.sv:67644:3
	assign gpio_toggle_gpio_toggle_29_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67645:3
	assign gpio_toggle_gpio_toggle_29_wd = reg_wdata[29];
	// Trace: design.sv:67647:3
	assign gpio_toggle_gpio_toggle_30_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67648:3
	assign gpio_toggle_gpio_toggle_30_wd = reg_wdata[30];
	// Trace: design.sv:67650:3
	assign gpio_toggle_gpio_toggle_31_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:67651:3
	assign gpio_toggle_gpio_toggle_31_wd = reg_wdata[31];
	// Trace: design.sv:67653:3
	assign intrpt_rise_en_intrpt_rise_en_0_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67654:3
	assign intrpt_rise_en_intrpt_rise_en_0_wd = reg_wdata[0];
	// Trace: design.sv:67656:3
	assign intrpt_rise_en_intrpt_rise_en_1_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67657:3
	assign intrpt_rise_en_intrpt_rise_en_1_wd = reg_wdata[1];
	// Trace: design.sv:67659:3
	assign intrpt_rise_en_intrpt_rise_en_2_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67660:3
	assign intrpt_rise_en_intrpt_rise_en_2_wd = reg_wdata[2];
	// Trace: design.sv:67662:3
	assign intrpt_rise_en_intrpt_rise_en_3_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67663:3
	assign intrpt_rise_en_intrpt_rise_en_3_wd = reg_wdata[3];
	// Trace: design.sv:67665:3
	assign intrpt_rise_en_intrpt_rise_en_4_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67666:3
	assign intrpt_rise_en_intrpt_rise_en_4_wd = reg_wdata[4];
	// Trace: design.sv:67668:3
	assign intrpt_rise_en_intrpt_rise_en_5_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67669:3
	assign intrpt_rise_en_intrpt_rise_en_5_wd = reg_wdata[5];
	// Trace: design.sv:67671:3
	assign intrpt_rise_en_intrpt_rise_en_6_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67672:3
	assign intrpt_rise_en_intrpt_rise_en_6_wd = reg_wdata[6];
	// Trace: design.sv:67674:3
	assign intrpt_rise_en_intrpt_rise_en_7_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67675:3
	assign intrpt_rise_en_intrpt_rise_en_7_wd = reg_wdata[7];
	// Trace: design.sv:67677:3
	assign intrpt_rise_en_intrpt_rise_en_8_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67678:3
	assign intrpt_rise_en_intrpt_rise_en_8_wd = reg_wdata[8];
	// Trace: design.sv:67680:3
	assign intrpt_rise_en_intrpt_rise_en_9_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67681:3
	assign intrpt_rise_en_intrpt_rise_en_9_wd = reg_wdata[9];
	// Trace: design.sv:67683:3
	assign intrpt_rise_en_intrpt_rise_en_10_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67684:3
	assign intrpt_rise_en_intrpt_rise_en_10_wd = reg_wdata[10];
	// Trace: design.sv:67686:3
	assign intrpt_rise_en_intrpt_rise_en_11_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67687:3
	assign intrpt_rise_en_intrpt_rise_en_11_wd = reg_wdata[11];
	// Trace: design.sv:67689:3
	assign intrpt_rise_en_intrpt_rise_en_12_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67690:3
	assign intrpt_rise_en_intrpt_rise_en_12_wd = reg_wdata[12];
	// Trace: design.sv:67692:3
	assign intrpt_rise_en_intrpt_rise_en_13_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67693:3
	assign intrpt_rise_en_intrpt_rise_en_13_wd = reg_wdata[13];
	// Trace: design.sv:67695:3
	assign intrpt_rise_en_intrpt_rise_en_14_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67696:3
	assign intrpt_rise_en_intrpt_rise_en_14_wd = reg_wdata[14];
	// Trace: design.sv:67698:3
	assign intrpt_rise_en_intrpt_rise_en_15_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67699:3
	assign intrpt_rise_en_intrpt_rise_en_15_wd = reg_wdata[15];
	// Trace: design.sv:67701:3
	assign intrpt_rise_en_intrpt_rise_en_16_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67702:3
	assign intrpt_rise_en_intrpt_rise_en_16_wd = reg_wdata[16];
	// Trace: design.sv:67704:3
	assign intrpt_rise_en_intrpt_rise_en_17_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67705:3
	assign intrpt_rise_en_intrpt_rise_en_17_wd = reg_wdata[17];
	// Trace: design.sv:67707:3
	assign intrpt_rise_en_intrpt_rise_en_18_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67708:3
	assign intrpt_rise_en_intrpt_rise_en_18_wd = reg_wdata[18];
	// Trace: design.sv:67710:3
	assign intrpt_rise_en_intrpt_rise_en_19_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67711:3
	assign intrpt_rise_en_intrpt_rise_en_19_wd = reg_wdata[19];
	// Trace: design.sv:67713:3
	assign intrpt_rise_en_intrpt_rise_en_20_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67714:3
	assign intrpt_rise_en_intrpt_rise_en_20_wd = reg_wdata[20];
	// Trace: design.sv:67716:3
	assign intrpt_rise_en_intrpt_rise_en_21_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67717:3
	assign intrpt_rise_en_intrpt_rise_en_21_wd = reg_wdata[21];
	// Trace: design.sv:67719:3
	assign intrpt_rise_en_intrpt_rise_en_22_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67720:3
	assign intrpt_rise_en_intrpt_rise_en_22_wd = reg_wdata[22];
	// Trace: design.sv:67722:3
	assign intrpt_rise_en_intrpt_rise_en_23_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67723:3
	assign intrpt_rise_en_intrpt_rise_en_23_wd = reg_wdata[23];
	// Trace: design.sv:67725:3
	assign intrpt_rise_en_intrpt_rise_en_24_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67726:3
	assign intrpt_rise_en_intrpt_rise_en_24_wd = reg_wdata[24];
	// Trace: design.sv:67728:3
	assign intrpt_rise_en_intrpt_rise_en_25_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67729:3
	assign intrpt_rise_en_intrpt_rise_en_25_wd = reg_wdata[25];
	// Trace: design.sv:67731:3
	assign intrpt_rise_en_intrpt_rise_en_26_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67732:3
	assign intrpt_rise_en_intrpt_rise_en_26_wd = reg_wdata[26];
	// Trace: design.sv:67734:3
	assign intrpt_rise_en_intrpt_rise_en_27_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67735:3
	assign intrpt_rise_en_intrpt_rise_en_27_wd = reg_wdata[27];
	// Trace: design.sv:67737:3
	assign intrpt_rise_en_intrpt_rise_en_28_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67738:3
	assign intrpt_rise_en_intrpt_rise_en_28_wd = reg_wdata[28];
	// Trace: design.sv:67740:3
	assign intrpt_rise_en_intrpt_rise_en_29_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67741:3
	assign intrpt_rise_en_intrpt_rise_en_29_wd = reg_wdata[29];
	// Trace: design.sv:67743:3
	assign intrpt_rise_en_intrpt_rise_en_30_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67744:3
	assign intrpt_rise_en_intrpt_rise_en_30_wd = reg_wdata[30];
	// Trace: design.sv:67746:3
	assign intrpt_rise_en_intrpt_rise_en_31_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:67747:3
	assign intrpt_rise_en_intrpt_rise_en_31_wd = reg_wdata[31];
	// Trace: design.sv:67749:3
	assign intrpt_fall_en_intrpt_fall_en_0_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67750:3
	assign intrpt_fall_en_intrpt_fall_en_0_wd = reg_wdata[0];
	// Trace: design.sv:67752:3
	assign intrpt_fall_en_intrpt_fall_en_1_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67753:3
	assign intrpt_fall_en_intrpt_fall_en_1_wd = reg_wdata[1];
	// Trace: design.sv:67755:3
	assign intrpt_fall_en_intrpt_fall_en_2_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67756:3
	assign intrpt_fall_en_intrpt_fall_en_2_wd = reg_wdata[2];
	// Trace: design.sv:67758:3
	assign intrpt_fall_en_intrpt_fall_en_3_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67759:3
	assign intrpt_fall_en_intrpt_fall_en_3_wd = reg_wdata[3];
	// Trace: design.sv:67761:3
	assign intrpt_fall_en_intrpt_fall_en_4_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67762:3
	assign intrpt_fall_en_intrpt_fall_en_4_wd = reg_wdata[4];
	// Trace: design.sv:67764:3
	assign intrpt_fall_en_intrpt_fall_en_5_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67765:3
	assign intrpt_fall_en_intrpt_fall_en_5_wd = reg_wdata[5];
	// Trace: design.sv:67767:3
	assign intrpt_fall_en_intrpt_fall_en_6_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67768:3
	assign intrpt_fall_en_intrpt_fall_en_6_wd = reg_wdata[6];
	// Trace: design.sv:67770:3
	assign intrpt_fall_en_intrpt_fall_en_7_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67771:3
	assign intrpt_fall_en_intrpt_fall_en_7_wd = reg_wdata[7];
	// Trace: design.sv:67773:3
	assign intrpt_fall_en_intrpt_fall_en_8_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67774:3
	assign intrpt_fall_en_intrpt_fall_en_8_wd = reg_wdata[8];
	// Trace: design.sv:67776:3
	assign intrpt_fall_en_intrpt_fall_en_9_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67777:3
	assign intrpt_fall_en_intrpt_fall_en_9_wd = reg_wdata[9];
	// Trace: design.sv:67779:3
	assign intrpt_fall_en_intrpt_fall_en_10_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67780:3
	assign intrpt_fall_en_intrpt_fall_en_10_wd = reg_wdata[10];
	// Trace: design.sv:67782:3
	assign intrpt_fall_en_intrpt_fall_en_11_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67783:3
	assign intrpt_fall_en_intrpt_fall_en_11_wd = reg_wdata[11];
	// Trace: design.sv:67785:3
	assign intrpt_fall_en_intrpt_fall_en_12_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67786:3
	assign intrpt_fall_en_intrpt_fall_en_12_wd = reg_wdata[12];
	// Trace: design.sv:67788:3
	assign intrpt_fall_en_intrpt_fall_en_13_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67789:3
	assign intrpt_fall_en_intrpt_fall_en_13_wd = reg_wdata[13];
	// Trace: design.sv:67791:3
	assign intrpt_fall_en_intrpt_fall_en_14_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67792:3
	assign intrpt_fall_en_intrpt_fall_en_14_wd = reg_wdata[14];
	// Trace: design.sv:67794:3
	assign intrpt_fall_en_intrpt_fall_en_15_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67795:3
	assign intrpt_fall_en_intrpt_fall_en_15_wd = reg_wdata[15];
	// Trace: design.sv:67797:3
	assign intrpt_fall_en_intrpt_fall_en_16_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67798:3
	assign intrpt_fall_en_intrpt_fall_en_16_wd = reg_wdata[16];
	// Trace: design.sv:67800:3
	assign intrpt_fall_en_intrpt_fall_en_17_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67801:3
	assign intrpt_fall_en_intrpt_fall_en_17_wd = reg_wdata[17];
	// Trace: design.sv:67803:3
	assign intrpt_fall_en_intrpt_fall_en_18_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67804:3
	assign intrpt_fall_en_intrpt_fall_en_18_wd = reg_wdata[18];
	// Trace: design.sv:67806:3
	assign intrpt_fall_en_intrpt_fall_en_19_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67807:3
	assign intrpt_fall_en_intrpt_fall_en_19_wd = reg_wdata[19];
	// Trace: design.sv:67809:3
	assign intrpt_fall_en_intrpt_fall_en_20_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67810:3
	assign intrpt_fall_en_intrpt_fall_en_20_wd = reg_wdata[20];
	// Trace: design.sv:67812:3
	assign intrpt_fall_en_intrpt_fall_en_21_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67813:3
	assign intrpt_fall_en_intrpt_fall_en_21_wd = reg_wdata[21];
	// Trace: design.sv:67815:3
	assign intrpt_fall_en_intrpt_fall_en_22_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67816:3
	assign intrpt_fall_en_intrpt_fall_en_22_wd = reg_wdata[22];
	// Trace: design.sv:67818:3
	assign intrpt_fall_en_intrpt_fall_en_23_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67819:3
	assign intrpt_fall_en_intrpt_fall_en_23_wd = reg_wdata[23];
	// Trace: design.sv:67821:3
	assign intrpt_fall_en_intrpt_fall_en_24_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67822:3
	assign intrpt_fall_en_intrpt_fall_en_24_wd = reg_wdata[24];
	// Trace: design.sv:67824:3
	assign intrpt_fall_en_intrpt_fall_en_25_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67825:3
	assign intrpt_fall_en_intrpt_fall_en_25_wd = reg_wdata[25];
	// Trace: design.sv:67827:3
	assign intrpt_fall_en_intrpt_fall_en_26_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67828:3
	assign intrpt_fall_en_intrpt_fall_en_26_wd = reg_wdata[26];
	// Trace: design.sv:67830:3
	assign intrpt_fall_en_intrpt_fall_en_27_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67831:3
	assign intrpt_fall_en_intrpt_fall_en_27_wd = reg_wdata[27];
	// Trace: design.sv:67833:3
	assign intrpt_fall_en_intrpt_fall_en_28_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67834:3
	assign intrpt_fall_en_intrpt_fall_en_28_wd = reg_wdata[28];
	// Trace: design.sv:67836:3
	assign intrpt_fall_en_intrpt_fall_en_29_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67837:3
	assign intrpt_fall_en_intrpt_fall_en_29_wd = reg_wdata[29];
	// Trace: design.sv:67839:3
	assign intrpt_fall_en_intrpt_fall_en_30_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67840:3
	assign intrpt_fall_en_intrpt_fall_en_30_wd = reg_wdata[30];
	// Trace: design.sv:67842:3
	assign intrpt_fall_en_intrpt_fall_en_31_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:67843:3
	assign intrpt_fall_en_intrpt_fall_en_31_wd = reg_wdata[31];
	// Trace: design.sv:67845:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_0_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67846:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_0_wd = reg_wdata[0];
	// Trace: design.sv:67848:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_1_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67849:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_1_wd = reg_wdata[1];
	// Trace: design.sv:67851:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_2_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67852:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_2_wd = reg_wdata[2];
	// Trace: design.sv:67854:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_3_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67855:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_3_wd = reg_wdata[3];
	// Trace: design.sv:67857:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_4_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67858:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_4_wd = reg_wdata[4];
	// Trace: design.sv:67860:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_5_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67861:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_5_wd = reg_wdata[5];
	// Trace: design.sv:67863:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_6_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67864:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_6_wd = reg_wdata[6];
	// Trace: design.sv:67866:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_7_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67867:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_7_wd = reg_wdata[7];
	// Trace: design.sv:67869:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_8_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67870:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_8_wd = reg_wdata[8];
	// Trace: design.sv:67872:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_9_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67873:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_9_wd = reg_wdata[9];
	// Trace: design.sv:67875:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_10_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67876:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_10_wd = reg_wdata[10];
	// Trace: design.sv:67878:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_11_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67879:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_11_wd = reg_wdata[11];
	// Trace: design.sv:67881:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_12_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67882:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_12_wd = reg_wdata[12];
	// Trace: design.sv:67884:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_13_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67885:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_13_wd = reg_wdata[13];
	// Trace: design.sv:67887:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_14_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67888:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_14_wd = reg_wdata[14];
	// Trace: design.sv:67890:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_15_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67891:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_15_wd = reg_wdata[15];
	// Trace: design.sv:67893:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_16_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67894:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_16_wd = reg_wdata[16];
	// Trace: design.sv:67896:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_17_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67897:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_17_wd = reg_wdata[17];
	// Trace: design.sv:67899:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_18_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67900:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_18_wd = reg_wdata[18];
	// Trace: design.sv:67902:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_19_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67903:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_19_wd = reg_wdata[19];
	// Trace: design.sv:67905:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_20_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67906:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_20_wd = reg_wdata[20];
	// Trace: design.sv:67908:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_21_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67909:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_21_wd = reg_wdata[21];
	// Trace: design.sv:67911:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_22_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67912:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_22_wd = reg_wdata[22];
	// Trace: design.sv:67914:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_23_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67915:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_23_wd = reg_wdata[23];
	// Trace: design.sv:67917:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_24_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67918:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_24_wd = reg_wdata[24];
	// Trace: design.sv:67920:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_25_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67921:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_25_wd = reg_wdata[25];
	// Trace: design.sv:67923:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_26_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67924:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_26_wd = reg_wdata[26];
	// Trace: design.sv:67926:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_27_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67927:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_27_wd = reg_wdata[27];
	// Trace: design.sv:67929:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_28_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67930:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_28_wd = reg_wdata[28];
	// Trace: design.sv:67932:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_29_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67933:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_29_wd = reg_wdata[29];
	// Trace: design.sv:67935:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_30_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67936:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_30_wd = reg_wdata[30];
	// Trace: design.sv:67938:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_31_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:67939:3
	assign intrpt_lvl_high_en_intrpt_lvl_high_en_31_wd = reg_wdata[31];
	// Trace: design.sv:67941:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_0_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67942:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_0_wd = reg_wdata[0];
	// Trace: design.sv:67944:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_1_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67945:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_1_wd = reg_wdata[1];
	// Trace: design.sv:67947:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_2_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67948:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_2_wd = reg_wdata[2];
	// Trace: design.sv:67950:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_3_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67951:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_3_wd = reg_wdata[3];
	// Trace: design.sv:67953:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_4_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67954:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_4_wd = reg_wdata[4];
	// Trace: design.sv:67956:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_5_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67957:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_5_wd = reg_wdata[5];
	// Trace: design.sv:67959:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_6_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67960:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_6_wd = reg_wdata[6];
	// Trace: design.sv:67962:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_7_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67963:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_7_wd = reg_wdata[7];
	// Trace: design.sv:67965:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_8_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67966:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_8_wd = reg_wdata[8];
	// Trace: design.sv:67968:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_9_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67969:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_9_wd = reg_wdata[9];
	// Trace: design.sv:67971:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_10_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67972:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_10_wd = reg_wdata[10];
	// Trace: design.sv:67974:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_11_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67975:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_11_wd = reg_wdata[11];
	// Trace: design.sv:67977:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_12_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67978:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_12_wd = reg_wdata[12];
	// Trace: design.sv:67980:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_13_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67981:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_13_wd = reg_wdata[13];
	// Trace: design.sv:67983:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_14_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67984:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_14_wd = reg_wdata[14];
	// Trace: design.sv:67986:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_15_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67987:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_15_wd = reg_wdata[15];
	// Trace: design.sv:67989:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_16_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67990:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_16_wd = reg_wdata[16];
	// Trace: design.sv:67992:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_17_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67993:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_17_wd = reg_wdata[17];
	// Trace: design.sv:67995:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_18_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67996:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_18_wd = reg_wdata[18];
	// Trace: design.sv:67998:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_19_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:67999:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_19_wd = reg_wdata[19];
	// Trace: design.sv:68001:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_20_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68002:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_20_wd = reg_wdata[20];
	// Trace: design.sv:68004:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_21_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68005:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_21_wd = reg_wdata[21];
	// Trace: design.sv:68007:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_22_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68008:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_22_wd = reg_wdata[22];
	// Trace: design.sv:68010:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_23_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68011:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_23_wd = reg_wdata[23];
	// Trace: design.sv:68013:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_24_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68014:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_24_wd = reg_wdata[24];
	// Trace: design.sv:68016:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_25_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68017:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_25_wd = reg_wdata[25];
	// Trace: design.sv:68019:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_26_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68020:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_26_wd = reg_wdata[26];
	// Trace: design.sv:68022:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_27_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68023:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_27_wd = reg_wdata[27];
	// Trace: design.sv:68025:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_28_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68026:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_28_wd = reg_wdata[28];
	// Trace: design.sv:68028:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_29_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68029:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_29_wd = reg_wdata[29];
	// Trace: design.sv:68031:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_30_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68032:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_30_wd = reg_wdata[30];
	// Trace: design.sv:68034:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_31_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:68035:3
	assign intrpt_lvl_low_en_intrpt_lvl_low_en_31_wd = reg_wdata[31];
	// Trace: design.sv:68037:3
	assign intrpt_status_intrpt_status_0_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68038:3
	assign intrpt_status_intrpt_status_0_wd = reg_wdata[0];
	// Trace: design.sv:68039:3
	assign intrpt_status_intrpt_status_0_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68041:3
	assign intrpt_status_intrpt_status_1_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68042:3
	assign intrpt_status_intrpt_status_1_wd = reg_wdata[1];
	// Trace: design.sv:68043:3
	assign intrpt_status_intrpt_status_1_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68045:3
	assign intrpt_status_intrpt_status_2_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68046:3
	assign intrpt_status_intrpt_status_2_wd = reg_wdata[2];
	// Trace: design.sv:68047:3
	assign intrpt_status_intrpt_status_2_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68049:3
	assign intrpt_status_intrpt_status_3_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68050:3
	assign intrpt_status_intrpt_status_3_wd = reg_wdata[3];
	// Trace: design.sv:68051:3
	assign intrpt_status_intrpt_status_3_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68053:3
	assign intrpt_status_intrpt_status_4_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68054:3
	assign intrpt_status_intrpt_status_4_wd = reg_wdata[4];
	// Trace: design.sv:68055:3
	assign intrpt_status_intrpt_status_4_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68057:3
	assign intrpt_status_intrpt_status_5_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68058:3
	assign intrpt_status_intrpt_status_5_wd = reg_wdata[5];
	// Trace: design.sv:68059:3
	assign intrpt_status_intrpt_status_5_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68061:3
	assign intrpt_status_intrpt_status_6_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68062:3
	assign intrpt_status_intrpt_status_6_wd = reg_wdata[6];
	// Trace: design.sv:68063:3
	assign intrpt_status_intrpt_status_6_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68065:3
	assign intrpt_status_intrpt_status_7_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68066:3
	assign intrpt_status_intrpt_status_7_wd = reg_wdata[7];
	// Trace: design.sv:68067:3
	assign intrpt_status_intrpt_status_7_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68069:3
	assign intrpt_status_intrpt_status_8_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68070:3
	assign intrpt_status_intrpt_status_8_wd = reg_wdata[8];
	// Trace: design.sv:68071:3
	assign intrpt_status_intrpt_status_8_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68073:3
	assign intrpt_status_intrpt_status_9_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68074:3
	assign intrpt_status_intrpt_status_9_wd = reg_wdata[9];
	// Trace: design.sv:68075:3
	assign intrpt_status_intrpt_status_9_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68077:3
	assign intrpt_status_intrpt_status_10_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68078:3
	assign intrpt_status_intrpt_status_10_wd = reg_wdata[10];
	// Trace: design.sv:68079:3
	assign intrpt_status_intrpt_status_10_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68081:3
	assign intrpt_status_intrpt_status_11_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68082:3
	assign intrpt_status_intrpt_status_11_wd = reg_wdata[11];
	// Trace: design.sv:68083:3
	assign intrpt_status_intrpt_status_11_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68085:3
	assign intrpt_status_intrpt_status_12_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68086:3
	assign intrpt_status_intrpt_status_12_wd = reg_wdata[12];
	// Trace: design.sv:68087:3
	assign intrpt_status_intrpt_status_12_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68089:3
	assign intrpt_status_intrpt_status_13_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68090:3
	assign intrpt_status_intrpt_status_13_wd = reg_wdata[13];
	// Trace: design.sv:68091:3
	assign intrpt_status_intrpt_status_13_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68093:3
	assign intrpt_status_intrpt_status_14_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68094:3
	assign intrpt_status_intrpt_status_14_wd = reg_wdata[14];
	// Trace: design.sv:68095:3
	assign intrpt_status_intrpt_status_14_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68097:3
	assign intrpt_status_intrpt_status_15_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68098:3
	assign intrpt_status_intrpt_status_15_wd = reg_wdata[15];
	// Trace: design.sv:68099:3
	assign intrpt_status_intrpt_status_15_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68101:3
	assign intrpt_status_intrpt_status_16_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68102:3
	assign intrpt_status_intrpt_status_16_wd = reg_wdata[16];
	// Trace: design.sv:68103:3
	assign intrpt_status_intrpt_status_16_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68105:3
	assign intrpt_status_intrpt_status_17_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68106:3
	assign intrpt_status_intrpt_status_17_wd = reg_wdata[17];
	// Trace: design.sv:68107:3
	assign intrpt_status_intrpt_status_17_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68109:3
	assign intrpt_status_intrpt_status_18_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68110:3
	assign intrpt_status_intrpt_status_18_wd = reg_wdata[18];
	// Trace: design.sv:68111:3
	assign intrpt_status_intrpt_status_18_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68113:3
	assign intrpt_status_intrpt_status_19_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68114:3
	assign intrpt_status_intrpt_status_19_wd = reg_wdata[19];
	// Trace: design.sv:68115:3
	assign intrpt_status_intrpt_status_19_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68117:3
	assign intrpt_status_intrpt_status_20_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68118:3
	assign intrpt_status_intrpt_status_20_wd = reg_wdata[20];
	// Trace: design.sv:68119:3
	assign intrpt_status_intrpt_status_20_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68121:3
	assign intrpt_status_intrpt_status_21_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68122:3
	assign intrpt_status_intrpt_status_21_wd = reg_wdata[21];
	// Trace: design.sv:68123:3
	assign intrpt_status_intrpt_status_21_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68125:3
	assign intrpt_status_intrpt_status_22_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68126:3
	assign intrpt_status_intrpt_status_22_wd = reg_wdata[22];
	// Trace: design.sv:68127:3
	assign intrpt_status_intrpt_status_22_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68129:3
	assign intrpt_status_intrpt_status_23_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68130:3
	assign intrpt_status_intrpt_status_23_wd = reg_wdata[23];
	// Trace: design.sv:68131:3
	assign intrpt_status_intrpt_status_23_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68133:3
	assign intrpt_status_intrpt_status_24_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68134:3
	assign intrpt_status_intrpt_status_24_wd = reg_wdata[24];
	// Trace: design.sv:68135:3
	assign intrpt_status_intrpt_status_24_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68137:3
	assign intrpt_status_intrpt_status_25_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68138:3
	assign intrpt_status_intrpt_status_25_wd = reg_wdata[25];
	// Trace: design.sv:68139:3
	assign intrpt_status_intrpt_status_25_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68141:3
	assign intrpt_status_intrpt_status_26_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68142:3
	assign intrpt_status_intrpt_status_26_wd = reg_wdata[26];
	// Trace: design.sv:68143:3
	assign intrpt_status_intrpt_status_26_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68145:3
	assign intrpt_status_intrpt_status_27_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68146:3
	assign intrpt_status_intrpt_status_27_wd = reg_wdata[27];
	// Trace: design.sv:68147:3
	assign intrpt_status_intrpt_status_27_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68149:3
	assign intrpt_status_intrpt_status_28_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68150:3
	assign intrpt_status_intrpt_status_28_wd = reg_wdata[28];
	// Trace: design.sv:68151:3
	assign intrpt_status_intrpt_status_28_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68153:3
	assign intrpt_status_intrpt_status_29_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68154:3
	assign intrpt_status_intrpt_status_29_wd = reg_wdata[29];
	// Trace: design.sv:68155:3
	assign intrpt_status_intrpt_status_29_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68157:3
	assign intrpt_status_intrpt_status_30_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68158:3
	assign intrpt_status_intrpt_status_30_wd = reg_wdata[30];
	// Trace: design.sv:68159:3
	assign intrpt_status_intrpt_status_30_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68161:3
	assign intrpt_status_intrpt_status_31_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:68162:3
	assign intrpt_status_intrpt_status_31_wd = reg_wdata[31];
	// Trace: design.sv:68163:3
	assign intrpt_status_intrpt_status_31_re = (addr_hit[14] & reg_re) & !reg_error;
	// Trace: design.sv:68165:3
	assign intrpt_rise_status_intrpt_rise_status_0_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68166:3
	assign intrpt_rise_status_intrpt_rise_status_0_wd = reg_wdata[0];
	// Trace: design.sv:68168:3
	assign intrpt_rise_status_intrpt_rise_status_1_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68169:3
	assign intrpt_rise_status_intrpt_rise_status_1_wd = reg_wdata[1];
	// Trace: design.sv:68171:3
	assign intrpt_rise_status_intrpt_rise_status_2_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68172:3
	assign intrpt_rise_status_intrpt_rise_status_2_wd = reg_wdata[2];
	// Trace: design.sv:68174:3
	assign intrpt_rise_status_intrpt_rise_status_3_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68175:3
	assign intrpt_rise_status_intrpt_rise_status_3_wd = reg_wdata[3];
	// Trace: design.sv:68177:3
	assign intrpt_rise_status_intrpt_rise_status_4_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68178:3
	assign intrpt_rise_status_intrpt_rise_status_4_wd = reg_wdata[4];
	// Trace: design.sv:68180:3
	assign intrpt_rise_status_intrpt_rise_status_5_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68181:3
	assign intrpt_rise_status_intrpt_rise_status_5_wd = reg_wdata[5];
	// Trace: design.sv:68183:3
	assign intrpt_rise_status_intrpt_rise_status_6_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68184:3
	assign intrpt_rise_status_intrpt_rise_status_6_wd = reg_wdata[6];
	// Trace: design.sv:68186:3
	assign intrpt_rise_status_intrpt_rise_status_7_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68187:3
	assign intrpt_rise_status_intrpt_rise_status_7_wd = reg_wdata[7];
	// Trace: design.sv:68189:3
	assign intrpt_rise_status_intrpt_rise_status_8_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68190:3
	assign intrpt_rise_status_intrpt_rise_status_8_wd = reg_wdata[8];
	// Trace: design.sv:68192:3
	assign intrpt_rise_status_intrpt_rise_status_9_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68193:3
	assign intrpt_rise_status_intrpt_rise_status_9_wd = reg_wdata[9];
	// Trace: design.sv:68195:3
	assign intrpt_rise_status_intrpt_rise_status_10_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68196:3
	assign intrpt_rise_status_intrpt_rise_status_10_wd = reg_wdata[10];
	// Trace: design.sv:68198:3
	assign intrpt_rise_status_intrpt_rise_status_11_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68199:3
	assign intrpt_rise_status_intrpt_rise_status_11_wd = reg_wdata[11];
	// Trace: design.sv:68201:3
	assign intrpt_rise_status_intrpt_rise_status_12_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68202:3
	assign intrpt_rise_status_intrpt_rise_status_12_wd = reg_wdata[12];
	// Trace: design.sv:68204:3
	assign intrpt_rise_status_intrpt_rise_status_13_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68205:3
	assign intrpt_rise_status_intrpt_rise_status_13_wd = reg_wdata[13];
	// Trace: design.sv:68207:3
	assign intrpt_rise_status_intrpt_rise_status_14_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68208:3
	assign intrpt_rise_status_intrpt_rise_status_14_wd = reg_wdata[14];
	// Trace: design.sv:68210:3
	assign intrpt_rise_status_intrpt_rise_status_15_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68211:3
	assign intrpt_rise_status_intrpt_rise_status_15_wd = reg_wdata[15];
	// Trace: design.sv:68213:3
	assign intrpt_rise_status_intrpt_rise_status_16_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68214:3
	assign intrpt_rise_status_intrpt_rise_status_16_wd = reg_wdata[16];
	// Trace: design.sv:68216:3
	assign intrpt_rise_status_intrpt_rise_status_17_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68217:3
	assign intrpt_rise_status_intrpt_rise_status_17_wd = reg_wdata[17];
	// Trace: design.sv:68219:3
	assign intrpt_rise_status_intrpt_rise_status_18_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68220:3
	assign intrpt_rise_status_intrpt_rise_status_18_wd = reg_wdata[18];
	// Trace: design.sv:68222:3
	assign intrpt_rise_status_intrpt_rise_status_19_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68223:3
	assign intrpt_rise_status_intrpt_rise_status_19_wd = reg_wdata[19];
	// Trace: design.sv:68225:3
	assign intrpt_rise_status_intrpt_rise_status_20_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68226:3
	assign intrpt_rise_status_intrpt_rise_status_20_wd = reg_wdata[20];
	// Trace: design.sv:68228:3
	assign intrpt_rise_status_intrpt_rise_status_21_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68229:3
	assign intrpt_rise_status_intrpt_rise_status_21_wd = reg_wdata[21];
	// Trace: design.sv:68231:3
	assign intrpt_rise_status_intrpt_rise_status_22_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68232:3
	assign intrpt_rise_status_intrpt_rise_status_22_wd = reg_wdata[22];
	// Trace: design.sv:68234:3
	assign intrpt_rise_status_intrpt_rise_status_23_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68235:3
	assign intrpt_rise_status_intrpt_rise_status_23_wd = reg_wdata[23];
	// Trace: design.sv:68237:3
	assign intrpt_rise_status_intrpt_rise_status_24_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68238:3
	assign intrpt_rise_status_intrpt_rise_status_24_wd = reg_wdata[24];
	// Trace: design.sv:68240:3
	assign intrpt_rise_status_intrpt_rise_status_25_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68241:3
	assign intrpt_rise_status_intrpt_rise_status_25_wd = reg_wdata[25];
	// Trace: design.sv:68243:3
	assign intrpt_rise_status_intrpt_rise_status_26_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68244:3
	assign intrpt_rise_status_intrpt_rise_status_26_wd = reg_wdata[26];
	// Trace: design.sv:68246:3
	assign intrpt_rise_status_intrpt_rise_status_27_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68247:3
	assign intrpt_rise_status_intrpt_rise_status_27_wd = reg_wdata[27];
	// Trace: design.sv:68249:3
	assign intrpt_rise_status_intrpt_rise_status_28_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68250:3
	assign intrpt_rise_status_intrpt_rise_status_28_wd = reg_wdata[28];
	// Trace: design.sv:68252:3
	assign intrpt_rise_status_intrpt_rise_status_29_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68253:3
	assign intrpt_rise_status_intrpt_rise_status_29_wd = reg_wdata[29];
	// Trace: design.sv:68255:3
	assign intrpt_rise_status_intrpt_rise_status_30_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68256:3
	assign intrpt_rise_status_intrpt_rise_status_30_wd = reg_wdata[30];
	// Trace: design.sv:68258:3
	assign intrpt_rise_status_intrpt_rise_status_31_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:68259:3
	assign intrpt_rise_status_intrpt_rise_status_31_wd = reg_wdata[31];
	// Trace: design.sv:68261:3
	assign intrpt_fall_status_intrpt_fall_status_0_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68262:3
	assign intrpt_fall_status_intrpt_fall_status_0_wd = reg_wdata[0];
	// Trace: design.sv:68264:3
	assign intrpt_fall_status_intrpt_fall_status_1_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68265:3
	assign intrpt_fall_status_intrpt_fall_status_1_wd = reg_wdata[1];
	// Trace: design.sv:68267:3
	assign intrpt_fall_status_intrpt_fall_status_2_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68268:3
	assign intrpt_fall_status_intrpt_fall_status_2_wd = reg_wdata[2];
	// Trace: design.sv:68270:3
	assign intrpt_fall_status_intrpt_fall_status_3_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68271:3
	assign intrpt_fall_status_intrpt_fall_status_3_wd = reg_wdata[3];
	// Trace: design.sv:68273:3
	assign intrpt_fall_status_intrpt_fall_status_4_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68274:3
	assign intrpt_fall_status_intrpt_fall_status_4_wd = reg_wdata[4];
	// Trace: design.sv:68276:3
	assign intrpt_fall_status_intrpt_fall_status_5_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68277:3
	assign intrpt_fall_status_intrpt_fall_status_5_wd = reg_wdata[5];
	// Trace: design.sv:68279:3
	assign intrpt_fall_status_intrpt_fall_status_6_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68280:3
	assign intrpt_fall_status_intrpt_fall_status_6_wd = reg_wdata[6];
	// Trace: design.sv:68282:3
	assign intrpt_fall_status_intrpt_fall_status_7_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68283:3
	assign intrpt_fall_status_intrpt_fall_status_7_wd = reg_wdata[7];
	// Trace: design.sv:68285:3
	assign intrpt_fall_status_intrpt_fall_status_8_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68286:3
	assign intrpt_fall_status_intrpt_fall_status_8_wd = reg_wdata[8];
	// Trace: design.sv:68288:3
	assign intrpt_fall_status_intrpt_fall_status_9_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68289:3
	assign intrpt_fall_status_intrpt_fall_status_9_wd = reg_wdata[9];
	// Trace: design.sv:68291:3
	assign intrpt_fall_status_intrpt_fall_status_10_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68292:3
	assign intrpt_fall_status_intrpt_fall_status_10_wd = reg_wdata[10];
	// Trace: design.sv:68294:3
	assign intrpt_fall_status_intrpt_fall_status_11_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68295:3
	assign intrpt_fall_status_intrpt_fall_status_11_wd = reg_wdata[11];
	// Trace: design.sv:68297:3
	assign intrpt_fall_status_intrpt_fall_status_12_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68298:3
	assign intrpt_fall_status_intrpt_fall_status_12_wd = reg_wdata[12];
	// Trace: design.sv:68300:3
	assign intrpt_fall_status_intrpt_fall_status_13_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68301:3
	assign intrpt_fall_status_intrpt_fall_status_13_wd = reg_wdata[13];
	// Trace: design.sv:68303:3
	assign intrpt_fall_status_intrpt_fall_status_14_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68304:3
	assign intrpt_fall_status_intrpt_fall_status_14_wd = reg_wdata[14];
	// Trace: design.sv:68306:3
	assign intrpt_fall_status_intrpt_fall_status_15_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68307:3
	assign intrpt_fall_status_intrpt_fall_status_15_wd = reg_wdata[15];
	// Trace: design.sv:68309:3
	assign intrpt_fall_status_intrpt_fall_status_16_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68310:3
	assign intrpt_fall_status_intrpt_fall_status_16_wd = reg_wdata[16];
	// Trace: design.sv:68312:3
	assign intrpt_fall_status_intrpt_fall_status_17_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68313:3
	assign intrpt_fall_status_intrpt_fall_status_17_wd = reg_wdata[17];
	// Trace: design.sv:68315:3
	assign intrpt_fall_status_intrpt_fall_status_18_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68316:3
	assign intrpt_fall_status_intrpt_fall_status_18_wd = reg_wdata[18];
	// Trace: design.sv:68318:3
	assign intrpt_fall_status_intrpt_fall_status_19_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68319:3
	assign intrpt_fall_status_intrpt_fall_status_19_wd = reg_wdata[19];
	// Trace: design.sv:68321:3
	assign intrpt_fall_status_intrpt_fall_status_20_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68322:3
	assign intrpt_fall_status_intrpt_fall_status_20_wd = reg_wdata[20];
	// Trace: design.sv:68324:3
	assign intrpt_fall_status_intrpt_fall_status_21_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68325:3
	assign intrpt_fall_status_intrpt_fall_status_21_wd = reg_wdata[21];
	// Trace: design.sv:68327:3
	assign intrpt_fall_status_intrpt_fall_status_22_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68328:3
	assign intrpt_fall_status_intrpt_fall_status_22_wd = reg_wdata[22];
	// Trace: design.sv:68330:3
	assign intrpt_fall_status_intrpt_fall_status_23_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68331:3
	assign intrpt_fall_status_intrpt_fall_status_23_wd = reg_wdata[23];
	// Trace: design.sv:68333:3
	assign intrpt_fall_status_intrpt_fall_status_24_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68334:3
	assign intrpt_fall_status_intrpt_fall_status_24_wd = reg_wdata[24];
	// Trace: design.sv:68336:3
	assign intrpt_fall_status_intrpt_fall_status_25_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68337:3
	assign intrpt_fall_status_intrpt_fall_status_25_wd = reg_wdata[25];
	// Trace: design.sv:68339:3
	assign intrpt_fall_status_intrpt_fall_status_26_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68340:3
	assign intrpt_fall_status_intrpt_fall_status_26_wd = reg_wdata[26];
	// Trace: design.sv:68342:3
	assign intrpt_fall_status_intrpt_fall_status_27_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68343:3
	assign intrpt_fall_status_intrpt_fall_status_27_wd = reg_wdata[27];
	// Trace: design.sv:68345:3
	assign intrpt_fall_status_intrpt_fall_status_28_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68346:3
	assign intrpt_fall_status_intrpt_fall_status_28_wd = reg_wdata[28];
	// Trace: design.sv:68348:3
	assign intrpt_fall_status_intrpt_fall_status_29_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68349:3
	assign intrpt_fall_status_intrpt_fall_status_29_wd = reg_wdata[29];
	// Trace: design.sv:68351:3
	assign intrpt_fall_status_intrpt_fall_status_30_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68352:3
	assign intrpt_fall_status_intrpt_fall_status_30_wd = reg_wdata[30];
	// Trace: design.sv:68354:3
	assign intrpt_fall_status_intrpt_fall_status_31_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:68355:3
	assign intrpt_fall_status_intrpt_fall_status_31_wd = reg_wdata[31];
	// Trace: design.sv:68357:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_0_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68358:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_0_wd = reg_wdata[0];
	// Trace: design.sv:68360:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_1_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68361:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_1_wd = reg_wdata[1];
	// Trace: design.sv:68363:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_2_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68364:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_2_wd = reg_wdata[2];
	// Trace: design.sv:68366:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_3_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68367:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_3_wd = reg_wdata[3];
	// Trace: design.sv:68369:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_4_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68370:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_4_wd = reg_wdata[4];
	// Trace: design.sv:68372:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_5_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68373:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_5_wd = reg_wdata[5];
	// Trace: design.sv:68375:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_6_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68376:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_6_wd = reg_wdata[6];
	// Trace: design.sv:68378:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_7_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68379:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_7_wd = reg_wdata[7];
	// Trace: design.sv:68381:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_8_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68382:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_8_wd = reg_wdata[8];
	// Trace: design.sv:68384:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_9_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68385:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_9_wd = reg_wdata[9];
	// Trace: design.sv:68387:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_10_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68388:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_10_wd = reg_wdata[10];
	// Trace: design.sv:68390:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_11_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68391:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_11_wd = reg_wdata[11];
	// Trace: design.sv:68393:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_12_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68394:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_12_wd = reg_wdata[12];
	// Trace: design.sv:68396:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_13_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68397:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_13_wd = reg_wdata[13];
	// Trace: design.sv:68399:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_14_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68400:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_14_wd = reg_wdata[14];
	// Trace: design.sv:68402:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_15_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68403:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_15_wd = reg_wdata[15];
	// Trace: design.sv:68405:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_16_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68406:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_16_wd = reg_wdata[16];
	// Trace: design.sv:68408:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_17_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68409:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_17_wd = reg_wdata[17];
	// Trace: design.sv:68411:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_18_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68412:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_18_wd = reg_wdata[18];
	// Trace: design.sv:68414:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_19_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68415:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_19_wd = reg_wdata[19];
	// Trace: design.sv:68417:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_20_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68418:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_20_wd = reg_wdata[20];
	// Trace: design.sv:68420:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_21_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68421:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_21_wd = reg_wdata[21];
	// Trace: design.sv:68423:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_22_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68424:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_22_wd = reg_wdata[22];
	// Trace: design.sv:68426:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_23_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68427:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_23_wd = reg_wdata[23];
	// Trace: design.sv:68429:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_24_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68430:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_24_wd = reg_wdata[24];
	// Trace: design.sv:68432:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_25_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68433:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_25_wd = reg_wdata[25];
	// Trace: design.sv:68435:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_26_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68436:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_26_wd = reg_wdata[26];
	// Trace: design.sv:68438:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_27_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68439:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_27_wd = reg_wdata[27];
	// Trace: design.sv:68441:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_28_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68442:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_28_wd = reg_wdata[28];
	// Trace: design.sv:68444:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_29_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68445:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_29_wd = reg_wdata[29];
	// Trace: design.sv:68447:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_30_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68448:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_30_wd = reg_wdata[30];
	// Trace: design.sv:68450:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_31_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:68451:3
	assign intrpt_lvl_high_status_intrpt_lvl_high_status_31_wd = reg_wdata[31];
	// Trace: design.sv:68453:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_0_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68454:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_0_wd = reg_wdata[0];
	// Trace: design.sv:68456:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_1_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68457:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_1_wd = reg_wdata[1];
	// Trace: design.sv:68459:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_2_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68460:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_2_wd = reg_wdata[2];
	// Trace: design.sv:68462:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_3_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68463:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_3_wd = reg_wdata[3];
	// Trace: design.sv:68465:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_4_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68466:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_4_wd = reg_wdata[4];
	// Trace: design.sv:68468:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_5_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68469:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_5_wd = reg_wdata[5];
	// Trace: design.sv:68471:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_6_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68472:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_6_wd = reg_wdata[6];
	// Trace: design.sv:68474:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_7_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68475:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_7_wd = reg_wdata[7];
	// Trace: design.sv:68477:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_8_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68478:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_8_wd = reg_wdata[8];
	// Trace: design.sv:68480:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_9_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68481:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_9_wd = reg_wdata[9];
	// Trace: design.sv:68483:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_10_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68484:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_10_wd = reg_wdata[10];
	// Trace: design.sv:68486:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_11_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68487:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_11_wd = reg_wdata[11];
	// Trace: design.sv:68489:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_12_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68490:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_12_wd = reg_wdata[12];
	// Trace: design.sv:68492:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_13_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68493:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_13_wd = reg_wdata[13];
	// Trace: design.sv:68495:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_14_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68496:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_14_wd = reg_wdata[14];
	// Trace: design.sv:68498:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_15_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68499:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_15_wd = reg_wdata[15];
	// Trace: design.sv:68501:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_16_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68502:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_16_wd = reg_wdata[16];
	// Trace: design.sv:68504:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_17_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68505:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_17_wd = reg_wdata[17];
	// Trace: design.sv:68507:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_18_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68508:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_18_wd = reg_wdata[18];
	// Trace: design.sv:68510:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_19_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68511:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_19_wd = reg_wdata[19];
	// Trace: design.sv:68513:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_20_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68514:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_20_wd = reg_wdata[20];
	// Trace: design.sv:68516:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_21_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68517:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_21_wd = reg_wdata[21];
	// Trace: design.sv:68519:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_22_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68520:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_22_wd = reg_wdata[22];
	// Trace: design.sv:68522:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_23_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68523:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_23_wd = reg_wdata[23];
	// Trace: design.sv:68525:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_24_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68526:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_24_wd = reg_wdata[24];
	// Trace: design.sv:68528:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_25_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68529:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_25_wd = reg_wdata[25];
	// Trace: design.sv:68531:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_26_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68532:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_26_wd = reg_wdata[26];
	// Trace: design.sv:68534:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_27_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68535:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_27_wd = reg_wdata[27];
	// Trace: design.sv:68537:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_28_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68538:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_28_wd = reg_wdata[28];
	// Trace: design.sv:68540:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_29_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68541:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_29_wd = reg_wdata[29];
	// Trace: design.sv:68543:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_30_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68544:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_30_wd = reg_wdata[30];
	// Trace: design.sv:68546:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_31_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:68547:3
	assign intrpt_lvl_low_status_intrpt_lvl_low_status_31_wd = reg_wdata[31];
	// Trace: design.sv:68550:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:68551:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:68552:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]: begin
				// Trace: design.sv:68554:9
				reg_rdata_next[9:0] = info_gpio_cnt_qs;
				// Trace: design.sv:68555:9
				reg_rdata_next[19:10] = info_version_qs;
			end
			addr_hit[1]: begin
				// Trace: design.sv:68559:9
				reg_rdata_next[0] = cfg_glbl_intrpt_mode_qs;
				// Trace: design.sv:68560:9
				reg_rdata_next[0] = cfg_pin_lvl_intrpt_mode_qs;
				// Trace: design.sv:68561:9
				reg_rdata_next[1] = cfg_reserved_qs;
			end
			addr_hit[2]: begin
				// Trace: design.sv:68565:9
				reg_rdata_next[1:0] = gpio_mode_0_mode_0_qs;
				// Trace: design.sv:68566:9
				reg_rdata_next[3:2] = gpio_mode_0_mode_1_qs;
				// Trace: design.sv:68567:9
				reg_rdata_next[5:4] = gpio_mode_0_mode_2_qs;
				// Trace: design.sv:68568:9
				reg_rdata_next[7:6] = gpio_mode_0_mode_3_qs;
				// Trace: design.sv:68569:9
				reg_rdata_next[9:8] = gpio_mode_0_mode_4_qs;
				// Trace: design.sv:68570:9
				reg_rdata_next[11:10] = gpio_mode_0_mode_5_qs;
				// Trace: design.sv:68571:9
				reg_rdata_next[13:12] = gpio_mode_0_mode_6_qs;
				// Trace: design.sv:68572:9
				reg_rdata_next[15:14] = gpio_mode_0_mode_7_qs;
				// Trace: design.sv:68573:9
				reg_rdata_next[17:16] = gpio_mode_0_mode_8_qs;
				// Trace: design.sv:68574:9
				reg_rdata_next[19:18] = gpio_mode_0_mode_9_qs;
				// Trace: design.sv:68575:9
				reg_rdata_next[21:20] = gpio_mode_0_mode_10_qs;
				// Trace: design.sv:68576:9
				reg_rdata_next[23:22] = gpio_mode_0_mode_11_qs;
				// Trace: design.sv:68577:9
				reg_rdata_next[25:24] = gpio_mode_0_mode_12_qs;
				// Trace: design.sv:68578:9
				reg_rdata_next[27:26] = gpio_mode_0_mode_13_qs;
				// Trace: design.sv:68579:9
				reg_rdata_next[29:28] = gpio_mode_0_mode_14_qs;
				// Trace: design.sv:68580:9
				reg_rdata_next[31:30] = gpio_mode_0_mode_15_qs;
			end
			addr_hit[3]: begin
				// Trace: design.sv:68584:9
				reg_rdata_next[1:0] = gpio_mode_1_mode_16_qs;
				// Trace: design.sv:68585:9
				reg_rdata_next[3:2] = gpio_mode_1_mode_17_qs;
				// Trace: design.sv:68586:9
				reg_rdata_next[5:4] = gpio_mode_1_mode_18_qs;
				// Trace: design.sv:68587:9
				reg_rdata_next[7:6] = gpio_mode_1_mode_19_qs;
				// Trace: design.sv:68588:9
				reg_rdata_next[9:8] = gpio_mode_1_mode_20_qs;
				// Trace: design.sv:68589:9
				reg_rdata_next[11:10] = gpio_mode_1_mode_21_qs;
				// Trace: design.sv:68590:9
				reg_rdata_next[13:12] = gpio_mode_1_mode_22_qs;
				// Trace: design.sv:68591:9
				reg_rdata_next[15:14] = gpio_mode_1_mode_23_qs;
				// Trace: design.sv:68592:9
				reg_rdata_next[17:16] = gpio_mode_1_mode_24_qs;
				// Trace: design.sv:68593:9
				reg_rdata_next[19:18] = gpio_mode_1_mode_25_qs;
				// Trace: design.sv:68594:9
				reg_rdata_next[21:20] = gpio_mode_1_mode_26_qs;
				// Trace: design.sv:68595:9
				reg_rdata_next[23:22] = gpio_mode_1_mode_27_qs;
				// Trace: design.sv:68596:9
				reg_rdata_next[25:24] = gpio_mode_1_mode_28_qs;
				// Trace: design.sv:68597:9
				reg_rdata_next[27:26] = gpio_mode_1_mode_29_qs;
				// Trace: design.sv:68598:9
				reg_rdata_next[29:28] = gpio_mode_1_mode_30_qs;
				// Trace: design.sv:68599:9
				reg_rdata_next[31:30] = gpio_mode_1_mode_31_qs;
			end
			addr_hit[4]: begin
				// Trace: design.sv:68603:9
				reg_rdata_next[0] = gpio_en_gpio_en_0_qs;
				// Trace: design.sv:68604:9
				reg_rdata_next[1] = gpio_en_gpio_en_1_qs;
				// Trace: design.sv:68605:9
				reg_rdata_next[2] = gpio_en_gpio_en_2_qs;
				// Trace: design.sv:68606:9
				reg_rdata_next[3] = gpio_en_gpio_en_3_qs;
				// Trace: design.sv:68607:9
				reg_rdata_next[4] = gpio_en_gpio_en_4_qs;
				// Trace: design.sv:68608:9
				reg_rdata_next[5] = gpio_en_gpio_en_5_qs;
				// Trace: design.sv:68609:9
				reg_rdata_next[6] = gpio_en_gpio_en_6_qs;
				// Trace: design.sv:68610:9
				reg_rdata_next[7] = gpio_en_gpio_en_7_qs;
				// Trace: design.sv:68611:9
				reg_rdata_next[8] = gpio_en_gpio_en_8_qs;
				// Trace: design.sv:68612:9
				reg_rdata_next[9] = gpio_en_gpio_en_9_qs;
				// Trace: design.sv:68613:9
				reg_rdata_next[10] = gpio_en_gpio_en_10_qs;
				// Trace: design.sv:68614:9
				reg_rdata_next[11] = gpio_en_gpio_en_11_qs;
				// Trace: design.sv:68615:9
				reg_rdata_next[12] = gpio_en_gpio_en_12_qs;
				// Trace: design.sv:68616:9
				reg_rdata_next[13] = gpio_en_gpio_en_13_qs;
				// Trace: design.sv:68617:9
				reg_rdata_next[14] = gpio_en_gpio_en_14_qs;
				// Trace: design.sv:68618:9
				reg_rdata_next[15] = gpio_en_gpio_en_15_qs;
				// Trace: design.sv:68619:9
				reg_rdata_next[16] = gpio_en_gpio_en_16_qs;
				// Trace: design.sv:68620:9
				reg_rdata_next[17] = gpio_en_gpio_en_17_qs;
				// Trace: design.sv:68621:9
				reg_rdata_next[18] = gpio_en_gpio_en_18_qs;
				// Trace: design.sv:68622:9
				reg_rdata_next[19] = gpio_en_gpio_en_19_qs;
				// Trace: design.sv:68623:9
				reg_rdata_next[20] = gpio_en_gpio_en_20_qs;
				// Trace: design.sv:68624:9
				reg_rdata_next[21] = gpio_en_gpio_en_21_qs;
				// Trace: design.sv:68625:9
				reg_rdata_next[22] = gpio_en_gpio_en_22_qs;
				// Trace: design.sv:68626:9
				reg_rdata_next[23] = gpio_en_gpio_en_23_qs;
				// Trace: design.sv:68627:9
				reg_rdata_next[24] = gpio_en_gpio_en_24_qs;
				// Trace: design.sv:68628:9
				reg_rdata_next[25] = gpio_en_gpio_en_25_qs;
				// Trace: design.sv:68629:9
				reg_rdata_next[26] = gpio_en_gpio_en_26_qs;
				// Trace: design.sv:68630:9
				reg_rdata_next[27] = gpio_en_gpio_en_27_qs;
				// Trace: design.sv:68631:9
				reg_rdata_next[28] = gpio_en_gpio_en_28_qs;
				// Trace: design.sv:68632:9
				reg_rdata_next[29] = gpio_en_gpio_en_29_qs;
				// Trace: design.sv:68633:9
				reg_rdata_next[30] = gpio_en_gpio_en_30_qs;
				// Trace: design.sv:68634:9
				reg_rdata_next[31] = gpio_en_gpio_en_31_qs;
			end
			addr_hit[5]: begin
				// Trace: design.sv:68638:9
				reg_rdata_next[0] = gpio_in_gpio_in_0_qs;
				// Trace: design.sv:68639:9
				reg_rdata_next[1] = gpio_in_gpio_in_1_qs;
				// Trace: design.sv:68640:9
				reg_rdata_next[2] = gpio_in_gpio_in_2_qs;
				// Trace: design.sv:68641:9
				reg_rdata_next[3] = gpio_in_gpio_in_3_qs;
				// Trace: design.sv:68642:9
				reg_rdata_next[4] = gpio_in_gpio_in_4_qs;
				// Trace: design.sv:68643:9
				reg_rdata_next[5] = gpio_in_gpio_in_5_qs;
				// Trace: design.sv:68644:9
				reg_rdata_next[6] = gpio_in_gpio_in_6_qs;
				// Trace: design.sv:68645:9
				reg_rdata_next[7] = gpio_in_gpio_in_7_qs;
				// Trace: design.sv:68646:9
				reg_rdata_next[8] = gpio_in_gpio_in_8_qs;
				// Trace: design.sv:68647:9
				reg_rdata_next[9] = gpio_in_gpio_in_9_qs;
				// Trace: design.sv:68648:9
				reg_rdata_next[10] = gpio_in_gpio_in_10_qs;
				// Trace: design.sv:68649:9
				reg_rdata_next[11] = gpio_in_gpio_in_11_qs;
				// Trace: design.sv:68650:9
				reg_rdata_next[12] = gpio_in_gpio_in_12_qs;
				// Trace: design.sv:68651:9
				reg_rdata_next[13] = gpio_in_gpio_in_13_qs;
				// Trace: design.sv:68652:9
				reg_rdata_next[14] = gpio_in_gpio_in_14_qs;
				// Trace: design.sv:68653:9
				reg_rdata_next[15] = gpio_in_gpio_in_15_qs;
				// Trace: design.sv:68654:9
				reg_rdata_next[16] = gpio_in_gpio_in_16_qs;
				// Trace: design.sv:68655:9
				reg_rdata_next[17] = gpio_in_gpio_in_17_qs;
				// Trace: design.sv:68656:9
				reg_rdata_next[18] = gpio_in_gpio_in_18_qs;
				// Trace: design.sv:68657:9
				reg_rdata_next[19] = gpio_in_gpio_in_19_qs;
				// Trace: design.sv:68658:9
				reg_rdata_next[20] = gpio_in_gpio_in_20_qs;
				// Trace: design.sv:68659:9
				reg_rdata_next[21] = gpio_in_gpio_in_21_qs;
				// Trace: design.sv:68660:9
				reg_rdata_next[22] = gpio_in_gpio_in_22_qs;
				// Trace: design.sv:68661:9
				reg_rdata_next[23] = gpio_in_gpio_in_23_qs;
				// Trace: design.sv:68662:9
				reg_rdata_next[24] = gpio_in_gpio_in_24_qs;
				// Trace: design.sv:68663:9
				reg_rdata_next[25] = gpio_in_gpio_in_25_qs;
				// Trace: design.sv:68664:9
				reg_rdata_next[26] = gpio_in_gpio_in_26_qs;
				// Trace: design.sv:68665:9
				reg_rdata_next[27] = gpio_in_gpio_in_27_qs;
				// Trace: design.sv:68666:9
				reg_rdata_next[28] = gpio_in_gpio_in_28_qs;
				// Trace: design.sv:68667:9
				reg_rdata_next[29] = gpio_in_gpio_in_29_qs;
				// Trace: design.sv:68668:9
				reg_rdata_next[30] = gpio_in_gpio_in_30_qs;
				// Trace: design.sv:68669:9
				reg_rdata_next[31] = gpio_in_gpio_in_31_qs;
			end
			addr_hit[6]: begin
				// Trace: design.sv:68673:9
				reg_rdata_next[0] = gpio_out_gpio_out_0_qs;
				// Trace: design.sv:68674:9
				reg_rdata_next[1] = gpio_out_gpio_out_1_qs;
				// Trace: design.sv:68675:9
				reg_rdata_next[2] = gpio_out_gpio_out_2_qs;
				// Trace: design.sv:68676:9
				reg_rdata_next[3] = gpio_out_gpio_out_3_qs;
				// Trace: design.sv:68677:9
				reg_rdata_next[4] = gpio_out_gpio_out_4_qs;
				// Trace: design.sv:68678:9
				reg_rdata_next[5] = gpio_out_gpio_out_5_qs;
				// Trace: design.sv:68679:9
				reg_rdata_next[6] = gpio_out_gpio_out_6_qs;
				// Trace: design.sv:68680:9
				reg_rdata_next[7] = gpio_out_gpio_out_7_qs;
				// Trace: design.sv:68681:9
				reg_rdata_next[8] = gpio_out_gpio_out_8_qs;
				// Trace: design.sv:68682:9
				reg_rdata_next[9] = gpio_out_gpio_out_9_qs;
				// Trace: design.sv:68683:9
				reg_rdata_next[10] = gpio_out_gpio_out_10_qs;
				// Trace: design.sv:68684:9
				reg_rdata_next[11] = gpio_out_gpio_out_11_qs;
				// Trace: design.sv:68685:9
				reg_rdata_next[12] = gpio_out_gpio_out_12_qs;
				// Trace: design.sv:68686:9
				reg_rdata_next[13] = gpio_out_gpio_out_13_qs;
				// Trace: design.sv:68687:9
				reg_rdata_next[14] = gpio_out_gpio_out_14_qs;
				// Trace: design.sv:68688:9
				reg_rdata_next[15] = gpio_out_gpio_out_15_qs;
				// Trace: design.sv:68689:9
				reg_rdata_next[16] = gpio_out_gpio_out_16_qs;
				// Trace: design.sv:68690:9
				reg_rdata_next[17] = gpio_out_gpio_out_17_qs;
				// Trace: design.sv:68691:9
				reg_rdata_next[18] = gpio_out_gpio_out_18_qs;
				// Trace: design.sv:68692:9
				reg_rdata_next[19] = gpio_out_gpio_out_19_qs;
				// Trace: design.sv:68693:9
				reg_rdata_next[20] = gpio_out_gpio_out_20_qs;
				// Trace: design.sv:68694:9
				reg_rdata_next[21] = gpio_out_gpio_out_21_qs;
				// Trace: design.sv:68695:9
				reg_rdata_next[22] = gpio_out_gpio_out_22_qs;
				// Trace: design.sv:68696:9
				reg_rdata_next[23] = gpio_out_gpio_out_23_qs;
				// Trace: design.sv:68697:9
				reg_rdata_next[24] = gpio_out_gpio_out_24_qs;
				// Trace: design.sv:68698:9
				reg_rdata_next[25] = gpio_out_gpio_out_25_qs;
				// Trace: design.sv:68699:9
				reg_rdata_next[26] = gpio_out_gpio_out_26_qs;
				// Trace: design.sv:68700:9
				reg_rdata_next[27] = gpio_out_gpio_out_27_qs;
				// Trace: design.sv:68701:9
				reg_rdata_next[28] = gpio_out_gpio_out_28_qs;
				// Trace: design.sv:68702:9
				reg_rdata_next[29] = gpio_out_gpio_out_29_qs;
				// Trace: design.sv:68703:9
				reg_rdata_next[30] = gpio_out_gpio_out_30_qs;
				// Trace: design.sv:68704:9
				reg_rdata_next[31] = gpio_out_gpio_out_31_qs;
			end
			addr_hit[7]: begin
				// Trace: design.sv:68708:9
				reg_rdata_next[0] = 1'sb0;
				// Trace: design.sv:68709:9
				reg_rdata_next[1] = 1'sb0;
				// Trace: design.sv:68710:9
				reg_rdata_next[2] = 1'sb0;
				// Trace: design.sv:68711:9
				reg_rdata_next[3] = 1'sb0;
				// Trace: design.sv:68712:9
				reg_rdata_next[4] = 1'sb0;
				// Trace: design.sv:68713:9
				reg_rdata_next[5] = 1'sb0;
				// Trace: design.sv:68714:9
				reg_rdata_next[6] = 1'sb0;
				// Trace: design.sv:68715:9
				reg_rdata_next[7] = 1'sb0;
				// Trace: design.sv:68716:9
				reg_rdata_next[8] = 1'sb0;
				// Trace: design.sv:68717:9
				reg_rdata_next[9] = 1'sb0;
				// Trace: design.sv:68718:9
				reg_rdata_next[10] = 1'sb0;
				// Trace: design.sv:68719:9
				reg_rdata_next[11] = 1'sb0;
				// Trace: design.sv:68720:9
				reg_rdata_next[12] = 1'sb0;
				// Trace: design.sv:68721:9
				reg_rdata_next[13] = 1'sb0;
				// Trace: design.sv:68722:9
				reg_rdata_next[14] = 1'sb0;
				// Trace: design.sv:68723:9
				reg_rdata_next[15] = 1'sb0;
				// Trace: design.sv:68724:9
				reg_rdata_next[16] = 1'sb0;
				// Trace: design.sv:68725:9
				reg_rdata_next[17] = 1'sb0;
				// Trace: design.sv:68726:9
				reg_rdata_next[18] = 1'sb0;
				// Trace: design.sv:68727:9
				reg_rdata_next[19] = 1'sb0;
				// Trace: design.sv:68728:9
				reg_rdata_next[20] = 1'sb0;
				// Trace: design.sv:68729:9
				reg_rdata_next[21] = 1'sb0;
				// Trace: design.sv:68730:9
				reg_rdata_next[22] = 1'sb0;
				// Trace: design.sv:68731:9
				reg_rdata_next[23] = 1'sb0;
				// Trace: design.sv:68732:9
				reg_rdata_next[24] = 1'sb0;
				// Trace: design.sv:68733:9
				reg_rdata_next[25] = 1'sb0;
				// Trace: design.sv:68734:9
				reg_rdata_next[26] = 1'sb0;
				// Trace: design.sv:68735:9
				reg_rdata_next[27] = 1'sb0;
				// Trace: design.sv:68736:9
				reg_rdata_next[28] = 1'sb0;
				// Trace: design.sv:68737:9
				reg_rdata_next[29] = 1'sb0;
				// Trace: design.sv:68738:9
				reg_rdata_next[30] = 1'sb0;
				// Trace: design.sv:68739:9
				reg_rdata_next[31] = 1'sb0;
			end
			addr_hit[8]: begin
				// Trace: design.sv:68743:9
				reg_rdata_next[0] = 1'sb0;
				// Trace: design.sv:68744:9
				reg_rdata_next[1] = 1'sb0;
				// Trace: design.sv:68745:9
				reg_rdata_next[2] = 1'sb0;
				// Trace: design.sv:68746:9
				reg_rdata_next[3] = 1'sb0;
				// Trace: design.sv:68747:9
				reg_rdata_next[4] = 1'sb0;
				// Trace: design.sv:68748:9
				reg_rdata_next[5] = 1'sb0;
				// Trace: design.sv:68749:9
				reg_rdata_next[6] = 1'sb0;
				// Trace: design.sv:68750:9
				reg_rdata_next[7] = 1'sb0;
				// Trace: design.sv:68751:9
				reg_rdata_next[8] = 1'sb0;
				// Trace: design.sv:68752:9
				reg_rdata_next[9] = 1'sb0;
				// Trace: design.sv:68753:9
				reg_rdata_next[10] = 1'sb0;
				// Trace: design.sv:68754:9
				reg_rdata_next[11] = 1'sb0;
				// Trace: design.sv:68755:9
				reg_rdata_next[12] = 1'sb0;
				// Trace: design.sv:68756:9
				reg_rdata_next[13] = 1'sb0;
				// Trace: design.sv:68757:9
				reg_rdata_next[14] = 1'sb0;
				// Trace: design.sv:68758:9
				reg_rdata_next[15] = 1'sb0;
				// Trace: design.sv:68759:9
				reg_rdata_next[16] = 1'sb0;
				// Trace: design.sv:68760:9
				reg_rdata_next[17] = 1'sb0;
				// Trace: design.sv:68761:9
				reg_rdata_next[18] = 1'sb0;
				// Trace: design.sv:68762:9
				reg_rdata_next[19] = 1'sb0;
				// Trace: design.sv:68763:9
				reg_rdata_next[20] = 1'sb0;
				// Trace: design.sv:68764:9
				reg_rdata_next[21] = 1'sb0;
				// Trace: design.sv:68765:9
				reg_rdata_next[22] = 1'sb0;
				// Trace: design.sv:68766:9
				reg_rdata_next[23] = 1'sb0;
				// Trace: design.sv:68767:9
				reg_rdata_next[24] = 1'sb0;
				// Trace: design.sv:68768:9
				reg_rdata_next[25] = 1'sb0;
				// Trace: design.sv:68769:9
				reg_rdata_next[26] = 1'sb0;
				// Trace: design.sv:68770:9
				reg_rdata_next[27] = 1'sb0;
				// Trace: design.sv:68771:9
				reg_rdata_next[28] = 1'sb0;
				// Trace: design.sv:68772:9
				reg_rdata_next[29] = 1'sb0;
				// Trace: design.sv:68773:9
				reg_rdata_next[30] = 1'sb0;
				// Trace: design.sv:68774:9
				reg_rdata_next[31] = 1'sb0;
			end
			addr_hit[9]: begin
				// Trace: design.sv:68778:9
				reg_rdata_next[0] = 1'sb0;
				// Trace: design.sv:68779:9
				reg_rdata_next[1] = 1'sb0;
				// Trace: design.sv:68780:9
				reg_rdata_next[2] = 1'sb0;
				// Trace: design.sv:68781:9
				reg_rdata_next[3] = 1'sb0;
				// Trace: design.sv:68782:9
				reg_rdata_next[4] = 1'sb0;
				// Trace: design.sv:68783:9
				reg_rdata_next[5] = 1'sb0;
				// Trace: design.sv:68784:9
				reg_rdata_next[6] = 1'sb0;
				// Trace: design.sv:68785:9
				reg_rdata_next[7] = 1'sb0;
				// Trace: design.sv:68786:9
				reg_rdata_next[8] = 1'sb0;
				// Trace: design.sv:68787:9
				reg_rdata_next[9] = 1'sb0;
				// Trace: design.sv:68788:9
				reg_rdata_next[10] = 1'sb0;
				// Trace: design.sv:68789:9
				reg_rdata_next[11] = 1'sb0;
				// Trace: design.sv:68790:9
				reg_rdata_next[12] = 1'sb0;
				// Trace: design.sv:68791:9
				reg_rdata_next[13] = 1'sb0;
				// Trace: design.sv:68792:9
				reg_rdata_next[14] = 1'sb0;
				// Trace: design.sv:68793:9
				reg_rdata_next[15] = 1'sb0;
				// Trace: design.sv:68794:9
				reg_rdata_next[16] = 1'sb0;
				// Trace: design.sv:68795:9
				reg_rdata_next[17] = 1'sb0;
				// Trace: design.sv:68796:9
				reg_rdata_next[18] = 1'sb0;
				// Trace: design.sv:68797:9
				reg_rdata_next[19] = 1'sb0;
				// Trace: design.sv:68798:9
				reg_rdata_next[20] = 1'sb0;
				// Trace: design.sv:68799:9
				reg_rdata_next[21] = 1'sb0;
				// Trace: design.sv:68800:9
				reg_rdata_next[22] = 1'sb0;
				// Trace: design.sv:68801:9
				reg_rdata_next[23] = 1'sb0;
				// Trace: design.sv:68802:9
				reg_rdata_next[24] = 1'sb0;
				// Trace: design.sv:68803:9
				reg_rdata_next[25] = 1'sb0;
				// Trace: design.sv:68804:9
				reg_rdata_next[26] = 1'sb0;
				// Trace: design.sv:68805:9
				reg_rdata_next[27] = 1'sb0;
				// Trace: design.sv:68806:9
				reg_rdata_next[28] = 1'sb0;
				// Trace: design.sv:68807:9
				reg_rdata_next[29] = 1'sb0;
				// Trace: design.sv:68808:9
				reg_rdata_next[30] = 1'sb0;
				// Trace: design.sv:68809:9
				reg_rdata_next[31] = 1'sb0;
			end
			addr_hit[10]: begin
				// Trace: design.sv:68813:9
				reg_rdata_next[0] = intrpt_rise_en_intrpt_rise_en_0_qs;
				// Trace: design.sv:68814:9
				reg_rdata_next[1] = intrpt_rise_en_intrpt_rise_en_1_qs;
				// Trace: design.sv:68815:9
				reg_rdata_next[2] = intrpt_rise_en_intrpt_rise_en_2_qs;
				// Trace: design.sv:68816:9
				reg_rdata_next[3] = intrpt_rise_en_intrpt_rise_en_3_qs;
				// Trace: design.sv:68817:9
				reg_rdata_next[4] = intrpt_rise_en_intrpt_rise_en_4_qs;
				// Trace: design.sv:68818:9
				reg_rdata_next[5] = intrpt_rise_en_intrpt_rise_en_5_qs;
				// Trace: design.sv:68819:9
				reg_rdata_next[6] = intrpt_rise_en_intrpt_rise_en_6_qs;
				// Trace: design.sv:68820:9
				reg_rdata_next[7] = intrpt_rise_en_intrpt_rise_en_7_qs;
				// Trace: design.sv:68821:9
				reg_rdata_next[8] = intrpt_rise_en_intrpt_rise_en_8_qs;
				// Trace: design.sv:68822:9
				reg_rdata_next[9] = intrpt_rise_en_intrpt_rise_en_9_qs;
				// Trace: design.sv:68823:9
				reg_rdata_next[10] = intrpt_rise_en_intrpt_rise_en_10_qs;
				// Trace: design.sv:68824:9
				reg_rdata_next[11] = intrpt_rise_en_intrpt_rise_en_11_qs;
				// Trace: design.sv:68825:9
				reg_rdata_next[12] = intrpt_rise_en_intrpt_rise_en_12_qs;
				// Trace: design.sv:68826:9
				reg_rdata_next[13] = intrpt_rise_en_intrpt_rise_en_13_qs;
				// Trace: design.sv:68827:9
				reg_rdata_next[14] = intrpt_rise_en_intrpt_rise_en_14_qs;
				// Trace: design.sv:68828:9
				reg_rdata_next[15] = intrpt_rise_en_intrpt_rise_en_15_qs;
				// Trace: design.sv:68829:9
				reg_rdata_next[16] = intrpt_rise_en_intrpt_rise_en_16_qs;
				// Trace: design.sv:68830:9
				reg_rdata_next[17] = intrpt_rise_en_intrpt_rise_en_17_qs;
				// Trace: design.sv:68831:9
				reg_rdata_next[18] = intrpt_rise_en_intrpt_rise_en_18_qs;
				// Trace: design.sv:68832:9
				reg_rdata_next[19] = intrpt_rise_en_intrpt_rise_en_19_qs;
				// Trace: design.sv:68833:9
				reg_rdata_next[20] = intrpt_rise_en_intrpt_rise_en_20_qs;
				// Trace: design.sv:68834:9
				reg_rdata_next[21] = intrpt_rise_en_intrpt_rise_en_21_qs;
				// Trace: design.sv:68835:9
				reg_rdata_next[22] = intrpt_rise_en_intrpt_rise_en_22_qs;
				// Trace: design.sv:68836:9
				reg_rdata_next[23] = intrpt_rise_en_intrpt_rise_en_23_qs;
				// Trace: design.sv:68837:9
				reg_rdata_next[24] = intrpt_rise_en_intrpt_rise_en_24_qs;
				// Trace: design.sv:68838:9
				reg_rdata_next[25] = intrpt_rise_en_intrpt_rise_en_25_qs;
				// Trace: design.sv:68839:9
				reg_rdata_next[26] = intrpt_rise_en_intrpt_rise_en_26_qs;
				// Trace: design.sv:68840:9
				reg_rdata_next[27] = intrpt_rise_en_intrpt_rise_en_27_qs;
				// Trace: design.sv:68841:9
				reg_rdata_next[28] = intrpt_rise_en_intrpt_rise_en_28_qs;
				// Trace: design.sv:68842:9
				reg_rdata_next[29] = intrpt_rise_en_intrpt_rise_en_29_qs;
				// Trace: design.sv:68843:9
				reg_rdata_next[30] = intrpt_rise_en_intrpt_rise_en_30_qs;
				// Trace: design.sv:68844:9
				reg_rdata_next[31] = intrpt_rise_en_intrpt_rise_en_31_qs;
			end
			addr_hit[11]: begin
				// Trace: design.sv:68848:9
				reg_rdata_next[0] = intrpt_fall_en_intrpt_fall_en_0_qs;
				// Trace: design.sv:68849:9
				reg_rdata_next[1] = intrpt_fall_en_intrpt_fall_en_1_qs;
				// Trace: design.sv:68850:9
				reg_rdata_next[2] = intrpt_fall_en_intrpt_fall_en_2_qs;
				// Trace: design.sv:68851:9
				reg_rdata_next[3] = intrpt_fall_en_intrpt_fall_en_3_qs;
				// Trace: design.sv:68852:9
				reg_rdata_next[4] = intrpt_fall_en_intrpt_fall_en_4_qs;
				// Trace: design.sv:68853:9
				reg_rdata_next[5] = intrpt_fall_en_intrpt_fall_en_5_qs;
				// Trace: design.sv:68854:9
				reg_rdata_next[6] = intrpt_fall_en_intrpt_fall_en_6_qs;
				// Trace: design.sv:68855:9
				reg_rdata_next[7] = intrpt_fall_en_intrpt_fall_en_7_qs;
				// Trace: design.sv:68856:9
				reg_rdata_next[8] = intrpt_fall_en_intrpt_fall_en_8_qs;
				// Trace: design.sv:68857:9
				reg_rdata_next[9] = intrpt_fall_en_intrpt_fall_en_9_qs;
				// Trace: design.sv:68858:9
				reg_rdata_next[10] = intrpt_fall_en_intrpt_fall_en_10_qs;
				// Trace: design.sv:68859:9
				reg_rdata_next[11] = intrpt_fall_en_intrpt_fall_en_11_qs;
				// Trace: design.sv:68860:9
				reg_rdata_next[12] = intrpt_fall_en_intrpt_fall_en_12_qs;
				// Trace: design.sv:68861:9
				reg_rdata_next[13] = intrpt_fall_en_intrpt_fall_en_13_qs;
				// Trace: design.sv:68862:9
				reg_rdata_next[14] = intrpt_fall_en_intrpt_fall_en_14_qs;
				// Trace: design.sv:68863:9
				reg_rdata_next[15] = intrpt_fall_en_intrpt_fall_en_15_qs;
				// Trace: design.sv:68864:9
				reg_rdata_next[16] = intrpt_fall_en_intrpt_fall_en_16_qs;
				// Trace: design.sv:68865:9
				reg_rdata_next[17] = intrpt_fall_en_intrpt_fall_en_17_qs;
				// Trace: design.sv:68866:9
				reg_rdata_next[18] = intrpt_fall_en_intrpt_fall_en_18_qs;
				// Trace: design.sv:68867:9
				reg_rdata_next[19] = intrpt_fall_en_intrpt_fall_en_19_qs;
				// Trace: design.sv:68868:9
				reg_rdata_next[20] = intrpt_fall_en_intrpt_fall_en_20_qs;
				// Trace: design.sv:68869:9
				reg_rdata_next[21] = intrpt_fall_en_intrpt_fall_en_21_qs;
				// Trace: design.sv:68870:9
				reg_rdata_next[22] = intrpt_fall_en_intrpt_fall_en_22_qs;
				// Trace: design.sv:68871:9
				reg_rdata_next[23] = intrpt_fall_en_intrpt_fall_en_23_qs;
				// Trace: design.sv:68872:9
				reg_rdata_next[24] = intrpt_fall_en_intrpt_fall_en_24_qs;
				// Trace: design.sv:68873:9
				reg_rdata_next[25] = intrpt_fall_en_intrpt_fall_en_25_qs;
				// Trace: design.sv:68874:9
				reg_rdata_next[26] = intrpt_fall_en_intrpt_fall_en_26_qs;
				// Trace: design.sv:68875:9
				reg_rdata_next[27] = intrpt_fall_en_intrpt_fall_en_27_qs;
				// Trace: design.sv:68876:9
				reg_rdata_next[28] = intrpt_fall_en_intrpt_fall_en_28_qs;
				// Trace: design.sv:68877:9
				reg_rdata_next[29] = intrpt_fall_en_intrpt_fall_en_29_qs;
				// Trace: design.sv:68878:9
				reg_rdata_next[30] = intrpt_fall_en_intrpt_fall_en_30_qs;
				// Trace: design.sv:68879:9
				reg_rdata_next[31] = intrpt_fall_en_intrpt_fall_en_31_qs;
			end
			addr_hit[12]: begin
				// Trace: design.sv:68883:9
				reg_rdata_next[0] = intrpt_lvl_high_en_intrpt_lvl_high_en_0_qs;
				// Trace: design.sv:68884:9
				reg_rdata_next[1] = intrpt_lvl_high_en_intrpt_lvl_high_en_1_qs;
				// Trace: design.sv:68885:9
				reg_rdata_next[2] = intrpt_lvl_high_en_intrpt_lvl_high_en_2_qs;
				// Trace: design.sv:68886:9
				reg_rdata_next[3] = intrpt_lvl_high_en_intrpt_lvl_high_en_3_qs;
				// Trace: design.sv:68887:9
				reg_rdata_next[4] = intrpt_lvl_high_en_intrpt_lvl_high_en_4_qs;
				// Trace: design.sv:68888:9
				reg_rdata_next[5] = intrpt_lvl_high_en_intrpt_lvl_high_en_5_qs;
				// Trace: design.sv:68889:9
				reg_rdata_next[6] = intrpt_lvl_high_en_intrpt_lvl_high_en_6_qs;
				// Trace: design.sv:68890:9
				reg_rdata_next[7] = intrpt_lvl_high_en_intrpt_lvl_high_en_7_qs;
				// Trace: design.sv:68891:9
				reg_rdata_next[8] = intrpt_lvl_high_en_intrpt_lvl_high_en_8_qs;
				// Trace: design.sv:68892:9
				reg_rdata_next[9] = intrpt_lvl_high_en_intrpt_lvl_high_en_9_qs;
				// Trace: design.sv:68893:9
				reg_rdata_next[10] = intrpt_lvl_high_en_intrpt_lvl_high_en_10_qs;
				// Trace: design.sv:68894:9
				reg_rdata_next[11] = intrpt_lvl_high_en_intrpt_lvl_high_en_11_qs;
				// Trace: design.sv:68895:9
				reg_rdata_next[12] = intrpt_lvl_high_en_intrpt_lvl_high_en_12_qs;
				// Trace: design.sv:68896:9
				reg_rdata_next[13] = intrpt_lvl_high_en_intrpt_lvl_high_en_13_qs;
				// Trace: design.sv:68897:9
				reg_rdata_next[14] = intrpt_lvl_high_en_intrpt_lvl_high_en_14_qs;
				// Trace: design.sv:68898:9
				reg_rdata_next[15] = intrpt_lvl_high_en_intrpt_lvl_high_en_15_qs;
				// Trace: design.sv:68899:9
				reg_rdata_next[16] = intrpt_lvl_high_en_intrpt_lvl_high_en_16_qs;
				// Trace: design.sv:68900:9
				reg_rdata_next[17] = intrpt_lvl_high_en_intrpt_lvl_high_en_17_qs;
				// Trace: design.sv:68901:9
				reg_rdata_next[18] = intrpt_lvl_high_en_intrpt_lvl_high_en_18_qs;
				// Trace: design.sv:68902:9
				reg_rdata_next[19] = intrpt_lvl_high_en_intrpt_lvl_high_en_19_qs;
				// Trace: design.sv:68903:9
				reg_rdata_next[20] = intrpt_lvl_high_en_intrpt_lvl_high_en_20_qs;
				// Trace: design.sv:68904:9
				reg_rdata_next[21] = intrpt_lvl_high_en_intrpt_lvl_high_en_21_qs;
				// Trace: design.sv:68905:9
				reg_rdata_next[22] = intrpt_lvl_high_en_intrpt_lvl_high_en_22_qs;
				// Trace: design.sv:68906:9
				reg_rdata_next[23] = intrpt_lvl_high_en_intrpt_lvl_high_en_23_qs;
				// Trace: design.sv:68907:9
				reg_rdata_next[24] = intrpt_lvl_high_en_intrpt_lvl_high_en_24_qs;
				// Trace: design.sv:68908:9
				reg_rdata_next[25] = intrpt_lvl_high_en_intrpt_lvl_high_en_25_qs;
				// Trace: design.sv:68909:9
				reg_rdata_next[26] = intrpt_lvl_high_en_intrpt_lvl_high_en_26_qs;
				// Trace: design.sv:68910:9
				reg_rdata_next[27] = intrpt_lvl_high_en_intrpt_lvl_high_en_27_qs;
				// Trace: design.sv:68911:9
				reg_rdata_next[28] = intrpt_lvl_high_en_intrpt_lvl_high_en_28_qs;
				// Trace: design.sv:68912:9
				reg_rdata_next[29] = intrpt_lvl_high_en_intrpt_lvl_high_en_29_qs;
				// Trace: design.sv:68913:9
				reg_rdata_next[30] = intrpt_lvl_high_en_intrpt_lvl_high_en_30_qs;
				// Trace: design.sv:68914:9
				reg_rdata_next[31] = intrpt_lvl_high_en_intrpt_lvl_high_en_31_qs;
			end
			addr_hit[13]: begin
				// Trace: design.sv:68918:9
				reg_rdata_next[0] = intrpt_lvl_low_en_intrpt_lvl_low_en_0_qs;
				// Trace: design.sv:68919:9
				reg_rdata_next[1] = intrpt_lvl_low_en_intrpt_lvl_low_en_1_qs;
				// Trace: design.sv:68920:9
				reg_rdata_next[2] = intrpt_lvl_low_en_intrpt_lvl_low_en_2_qs;
				// Trace: design.sv:68921:9
				reg_rdata_next[3] = intrpt_lvl_low_en_intrpt_lvl_low_en_3_qs;
				// Trace: design.sv:68922:9
				reg_rdata_next[4] = intrpt_lvl_low_en_intrpt_lvl_low_en_4_qs;
				// Trace: design.sv:68923:9
				reg_rdata_next[5] = intrpt_lvl_low_en_intrpt_lvl_low_en_5_qs;
				// Trace: design.sv:68924:9
				reg_rdata_next[6] = intrpt_lvl_low_en_intrpt_lvl_low_en_6_qs;
				// Trace: design.sv:68925:9
				reg_rdata_next[7] = intrpt_lvl_low_en_intrpt_lvl_low_en_7_qs;
				// Trace: design.sv:68926:9
				reg_rdata_next[8] = intrpt_lvl_low_en_intrpt_lvl_low_en_8_qs;
				// Trace: design.sv:68927:9
				reg_rdata_next[9] = intrpt_lvl_low_en_intrpt_lvl_low_en_9_qs;
				// Trace: design.sv:68928:9
				reg_rdata_next[10] = intrpt_lvl_low_en_intrpt_lvl_low_en_10_qs;
				// Trace: design.sv:68929:9
				reg_rdata_next[11] = intrpt_lvl_low_en_intrpt_lvl_low_en_11_qs;
				// Trace: design.sv:68930:9
				reg_rdata_next[12] = intrpt_lvl_low_en_intrpt_lvl_low_en_12_qs;
				// Trace: design.sv:68931:9
				reg_rdata_next[13] = intrpt_lvl_low_en_intrpt_lvl_low_en_13_qs;
				// Trace: design.sv:68932:9
				reg_rdata_next[14] = intrpt_lvl_low_en_intrpt_lvl_low_en_14_qs;
				// Trace: design.sv:68933:9
				reg_rdata_next[15] = intrpt_lvl_low_en_intrpt_lvl_low_en_15_qs;
				// Trace: design.sv:68934:9
				reg_rdata_next[16] = intrpt_lvl_low_en_intrpt_lvl_low_en_16_qs;
				// Trace: design.sv:68935:9
				reg_rdata_next[17] = intrpt_lvl_low_en_intrpt_lvl_low_en_17_qs;
				// Trace: design.sv:68936:9
				reg_rdata_next[18] = intrpt_lvl_low_en_intrpt_lvl_low_en_18_qs;
				// Trace: design.sv:68937:9
				reg_rdata_next[19] = intrpt_lvl_low_en_intrpt_lvl_low_en_19_qs;
				// Trace: design.sv:68938:9
				reg_rdata_next[20] = intrpt_lvl_low_en_intrpt_lvl_low_en_20_qs;
				// Trace: design.sv:68939:9
				reg_rdata_next[21] = intrpt_lvl_low_en_intrpt_lvl_low_en_21_qs;
				// Trace: design.sv:68940:9
				reg_rdata_next[22] = intrpt_lvl_low_en_intrpt_lvl_low_en_22_qs;
				// Trace: design.sv:68941:9
				reg_rdata_next[23] = intrpt_lvl_low_en_intrpt_lvl_low_en_23_qs;
				// Trace: design.sv:68942:9
				reg_rdata_next[24] = intrpt_lvl_low_en_intrpt_lvl_low_en_24_qs;
				// Trace: design.sv:68943:9
				reg_rdata_next[25] = intrpt_lvl_low_en_intrpt_lvl_low_en_25_qs;
				// Trace: design.sv:68944:9
				reg_rdata_next[26] = intrpt_lvl_low_en_intrpt_lvl_low_en_26_qs;
				// Trace: design.sv:68945:9
				reg_rdata_next[27] = intrpt_lvl_low_en_intrpt_lvl_low_en_27_qs;
				// Trace: design.sv:68946:9
				reg_rdata_next[28] = intrpt_lvl_low_en_intrpt_lvl_low_en_28_qs;
				// Trace: design.sv:68947:9
				reg_rdata_next[29] = intrpt_lvl_low_en_intrpt_lvl_low_en_29_qs;
				// Trace: design.sv:68948:9
				reg_rdata_next[30] = intrpt_lvl_low_en_intrpt_lvl_low_en_30_qs;
				// Trace: design.sv:68949:9
				reg_rdata_next[31] = intrpt_lvl_low_en_intrpt_lvl_low_en_31_qs;
			end
			addr_hit[14]: begin
				// Trace: design.sv:68953:9
				reg_rdata_next[0] = intrpt_status_intrpt_status_0_qs;
				// Trace: design.sv:68954:9
				reg_rdata_next[1] = intrpt_status_intrpt_status_1_qs;
				// Trace: design.sv:68955:9
				reg_rdata_next[2] = intrpt_status_intrpt_status_2_qs;
				// Trace: design.sv:68956:9
				reg_rdata_next[3] = intrpt_status_intrpt_status_3_qs;
				// Trace: design.sv:68957:9
				reg_rdata_next[4] = intrpt_status_intrpt_status_4_qs;
				// Trace: design.sv:68958:9
				reg_rdata_next[5] = intrpt_status_intrpt_status_5_qs;
				// Trace: design.sv:68959:9
				reg_rdata_next[6] = intrpt_status_intrpt_status_6_qs;
				// Trace: design.sv:68960:9
				reg_rdata_next[7] = intrpt_status_intrpt_status_7_qs;
				// Trace: design.sv:68961:9
				reg_rdata_next[8] = intrpt_status_intrpt_status_8_qs;
				// Trace: design.sv:68962:9
				reg_rdata_next[9] = intrpt_status_intrpt_status_9_qs;
				// Trace: design.sv:68963:9
				reg_rdata_next[10] = intrpt_status_intrpt_status_10_qs;
				// Trace: design.sv:68964:9
				reg_rdata_next[11] = intrpt_status_intrpt_status_11_qs;
				// Trace: design.sv:68965:9
				reg_rdata_next[12] = intrpt_status_intrpt_status_12_qs;
				// Trace: design.sv:68966:9
				reg_rdata_next[13] = intrpt_status_intrpt_status_13_qs;
				// Trace: design.sv:68967:9
				reg_rdata_next[14] = intrpt_status_intrpt_status_14_qs;
				// Trace: design.sv:68968:9
				reg_rdata_next[15] = intrpt_status_intrpt_status_15_qs;
				// Trace: design.sv:68969:9
				reg_rdata_next[16] = intrpt_status_intrpt_status_16_qs;
				// Trace: design.sv:68970:9
				reg_rdata_next[17] = intrpt_status_intrpt_status_17_qs;
				// Trace: design.sv:68971:9
				reg_rdata_next[18] = intrpt_status_intrpt_status_18_qs;
				// Trace: design.sv:68972:9
				reg_rdata_next[19] = intrpt_status_intrpt_status_19_qs;
				// Trace: design.sv:68973:9
				reg_rdata_next[20] = intrpt_status_intrpt_status_20_qs;
				// Trace: design.sv:68974:9
				reg_rdata_next[21] = intrpt_status_intrpt_status_21_qs;
				// Trace: design.sv:68975:9
				reg_rdata_next[22] = intrpt_status_intrpt_status_22_qs;
				// Trace: design.sv:68976:9
				reg_rdata_next[23] = intrpt_status_intrpt_status_23_qs;
				// Trace: design.sv:68977:9
				reg_rdata_next[24] = intrpt_status_intrpt_status_24_qs;
				// Trace: design.sv:68978:9
				reg_rdata_next[25] = intrpt_status_intrpt_status_25_qs;
				// Trace: design.sv:68979:9
				reg_rdata_next[26] = intrpt_status_intrpt_status_26_qs;
				// Trace: design.sv:68980:9
				reg_rdata_next[27] = intrpt_status_intrpt_status_27_qs;
				// Trace: design.sv:68981:9
				reg_rdata_next[28] = intrpt_status_intrpt_status_28_qs;
				// Trace: design.sv:68982:9
				reg_rdata_next[29] = intrpt_status_intrpt_status_29_qs;
				// Trace: design.sv:68983:9
				reg_rdata_next[30] = intrpt_status_intrpt_status_30_qs;
				// Trace: design.sv:68984:9
				reg_rdata_next[31] = intrpt_status_intrpt_status_31_qs;
			end
			addr_hit[15]: begin
				// Trace: design.sv:68988:9
				reg_rdata_next[0] = intrpt_rise_status_intrpt_rise_status_0_qs;
				// Trace: design.sv:68989:9
				reg_rdata_next[1] = intrpt_rise_status_intrpt_rise_status_1_qs;
				// Trace: design.sv:68990:9
				reg_rdata_next[2] = intrpt_rise_status_intrpt_rise_status_2_qs;
				// Trace: design.sv:68991:9
				reg_rdata_next[3] = intrpt_rise_status_intrpt_rise_status_3_qs;
				// Trace: design.sv:68992:9
				reg_rdata_next[4] = intrpt_rise_status_intrpt_rise_status_4_qs;
				// Trace: design.sv:68993:9
				reg_rdata_next[5] = intrpt_rise_status_intrpt_rise_status_5_qs;
				// Trace: design.sv:68994:9
				reg_rdata_next[6] = intrpt_rise_status_intrpt_rise_status_6_qs;
				// Trace: design.sv:68995:9
				reg_rdata_next[7] = intrpt_rise_status_intrpt_rise_status_7_qs;
				// Trace: design.sv:68996:9
				reg_rdata_next[8] = intrpt_rise_status_intrpt_rise_status_8_qs;
				// Trace: design.sv:68997:9
				reg_rdata_next[9] = intrpt_rise_status_intrpt_rise_status_9_qs;
				// Trace: design.sv:68998:9
				reg_rdata_next[10] = intrpt_rise_status_intrpt_rise_status_10_qs;
				// Trace: design.sv:68999:9
				reg_rdata_next[11] = intrpt_rise_status_intrpt_rise_status_11_qs;
				// Trace: design.sv:69000:9
				reg_rdata_next[12] = intrpt_rise_status_intrpt_rise_status_12_qs;
				// Trace: design.sv:69001:9
				reg_rdata_next[13] = intrpt_rise_status_intrpt_rise_status_13_qs;
				// Trace: design.sv:69002:9
				reg_rdata_next[14] = intrpt_rise_status_intrpt_rise_status_14_qs;
				// Trace: design.sv:69003:9
				reg_rdata_next[15] = intrpt_rise_status_intrpt_rise_status_15_qs;
				// Trace: design.sv:69004:9
				reg_rdata_next[16] = intrpt_rise_status_intrpt_rise_status_16_qs;
				// Trace: design.sv:69005:9
				reg_rdata_next[17] = intrpt_rise_status_intrpt_rise_status_17_qs;
				// Trace: design.sv:69006:9
				reg_rdata_next[18] = intrpt_rise_status_intrpt_rise_status_18_qs;
				// Trace: design.sv:69007:9
				reg_rdata_next[19] = intrpt_rise_status_intrpt_rise_status_19_qs;
				// Trace: design.sv:69008:9
				reg_rdata_next[20] = intrpt_rise_status_intrpt_rise_status_20_qs;
				// Trace: design.sv:69009:9
				reg_rdata_next[21] = intrpt_rise_status_intrpt_rise_status_21_qs;
				// Trace: design.sv:69010:9
				reg_rdata_next[22] = intrpt_rise_status_intrpt_rise_status_22_qs;
				// Trace: design.sv:69011:9
				reg_rdata_next[23] = intrpt_rise_status_intrpt_rise_status_23_qs;
				// Trace: design.sv:69012:9
				reg_rdata_next[24] = intrpt_rise_status_intrpt_rise_status_24_qs;
				// Trace: design.sv:69013:9
				reg_rdata_next[25] = intrpt_rise_status_intrpt_rise_status_25_qs;
				// Trace: design.sv:69014:9
				reg_rdata_next[26] = intrpt_rise_status_intrpt_rise_status_26_qs;
				// Trace: design.sv:69015:9
				reg_rdata_next[27] = intrpt_rise_status_intrpt_rise_status_27_qs;
				// Trace: design.sv:69016:9
				reg_rdata_next[28] = intrpt_rise_status_intrpt_rise_status_28_qs;
				// Trace: design.sv:69017:9
				reg_rdata_next[29] = intrpt_rise_status_intrpt_rise_status_29_qs;
				// Trace: design.sv:69018:9
				reg_rdata_next[30] = intrpt_rise_status_intrpt_rise_status_30_qs;
				// Trace: design.sv:69019:9
				reg_rdata_next[31] = intrpt_rise_status_intrpt_rise_status_31_qs;
			end
			addr_hit[16]: begin
				// Trace: design.sv:69023:9
				reg_rdata_next[0] = intrpt_fall_status_intrpt_fall_status_0_qs;
				// Trace: design.sv:69024:9
				reg_rdata_next[1] = intrpt_fall_status_intrpt_fall_status_1_qs;
				// Trace: design.sv:69025:9
				reg_rdata_next[2] = intrpt_fall_status_intrpt_fall_status_2_qs;
				// Trace: design.sv:69026:9
				reg_rdata_next[3] = intrpt_fall_status_intrpt_fall_status_3_qs;
				// Trace: design.sv:69027:9
				reg_rdata_next[4] = intrpt_fall_status_intrpt_fall_status_4_qs;
				// Trace: design.sv:69028:9
				reg_rdata_next[5] = intrpt_fall_status_intrpt_fall_status_5_qs;
				// Trace: design.sv:69029:9
				reg_rdata_next[6] = intrpt_fall_status_intrpt_fall_status_6_qs;
				// Trace: design.sv:69030:9
				reg_rdata_next[7] = intrpt_fall_status_intrpt_fall_status_7_qs;
				// Trace: design.sv:69031:9
				reg_rdata_next[8] = intrpt_fall_status_intrpt_fall_status_8_qs;
				// Trace: design.sv:69032:9
				reg_rdata_next[9] = intrpt_fall_status_intrpt_fall_status_9_qs;
				// Trace: design.sv:69033:9
				reg_rdata_next[10] = intrpt_fall_status_intrpt_fall_status_10_qs;
				// Trace: design.sv:69034:9
				reg_rdata_next[11] = intrpt_fall_status_intrpt_fall_status_11_qs;
				// Trace: design.sv:69035:9
				reg_rdata_next[12] = intrpt_fall_status_intrpt_fall_status_12_qs;
				// Trace: design.sv:69036:9
				reg_rdata_next[13] = intrpt_fall_status_intrpt_fall_status_13_qs;
				// Trace: design.sv:69037:9
				reg_rdata_next[14] = intrpt_fall_status_intrpt_fall_status_14_qs;
				// Trace: design.sv:69038:9
				reg_rdata_next[15] = intrpt_fall_status_intrpt_fall_status_15_qs;
				// Trace: design.sv:69039:9
				reg_rdata_next[16] = intrpt_fall_status_intrpt_fall_status_16_qs;
				// Trace: design.sv:69040:9
				reg_rdata_next[17] = intrpt_fall_status_intrpt_fall_status_17_qs;
				// Trace: design.sv:69041:9
				reg_rdata_next[18] = intrpt_fall_status_intrpt_fall_status_18_qs;
				// Trace: design.sv:69042:9
				reg_rdata_next[19] = intrpt_fall_status_intrpt_fall_status_19_qs;
				// Trace: design.sv:69043:9
				reg_rdata_next[20] = intrpt_fall_status_intrpt_fall_status_20_qs;
				// Trace: design.sv:69044:9
				reg_rdata_next[21] = intrpt_fall_status_intrpt_fall_status_21_qs;
				// Trace: design.sv:69045:9
				reg_rdata_next[22] = intrpt_fall_status_intrpt_fall_status_22_qs;
				// Trace: design.sv:69046:9
				reg_rdata_next[23] = intrpt_fall_status_intrpt_fall_status_23_qs;
				// Trace: design.sv:69047:9
				reg_rdata_next[24] = intrpt_fall_status_intrpt_fall_status_24_qs;
				// Trace: design.sv:69048:9
				reg_rdata_next[25] = intrpt_fall_status_intrpt_fall_status_25_qs;
				// Trace: design.sv:69049:9
				reg_rdata_next[26] = intrpt_fall_status_intrpt_fall_status_26_qs;
				// Trace: design.sv:69050:9
				reg_rdata_next[27] = intrpt_fall_status_intrpt_fall_status_27_qs;
				// Trace: design.sv:69051:9
				reg_rdata_next[28] = intrpt_fall_status_intrpt_fall_status_28_qs;
				// Trace: design.sv:69052:9
				reg_rdata_next[29] = intrpt_fall_status_intrpt_fall_status_29_qs;
				// Trace: design.sv:69053:9
				reg_rdata_next[30] = intrpt_fall_status_intrpt_fall_status_30_qs;
				// Trace: design.sv:69054:9
				reg_rdata_next[31] = intrpt_fall_status_intrpt_fall_status_31_qs;
			end
			addr_hit[17]: begin
				// Trace: design.sv:69058:9
				reg_rdata_next[0] = intrpt_lvl_high_status_intrpt_lvl_high_status_0_qs;
				// Trace: design.sv:69059:9
				reg_rdata_next[1] = intrpt_lvl_high_status_intrpt_lvl_high_status_1_qs;
				// Trace: design.sv:69060:9
				reg_rdata_next[2] = intrpt_lvl_high_status_intrpt_lvl_high_status_2_qs;
				// Trace: design.sv:69061:9
				reg_rdata_next[3] = intrpt_lvl_high_status_intrpt_lvl_high_status_3_qs;
				// Trace: design.sv:69062:9
				reg_rdata_next[4] = intrpt_lvl_high_status_intrpt_lvl_high_status_4_qs;
				// Trace: design.sv:69063:9
				reg_rdata_next[5] = intrpt_lvl_high_status_intrpt_lvl_high_status_5_qs;
				// Trace: design.sv:69064:9
				reg_rdata_next[6] = intrpt_lvl_high_status_intrpt_lvl_high_status_6_qs;
				// Trace: design.sv:69065:9
				reg_rdata_next[7] = intrpt_lvl_high_status_intrpt_lvl_high_status_7_qs;
				// Trace: design.sv:69066:9
				reg_rdata_next[8] = intrpt_lvl_high_status_intrpt_lvl_high_status_8_qs;
				// Trace: design.sv:69067:9
				reg_rdata_next[9] = intrpt_lvl_high_status_intrpt_lvl_high_status_9_qs;
				// Trace: design.sv:69068:9
				reg_rdata_next[10] = intrpt_lvl_high_status_intrpt_lvl_high_status_10_qs;
				// Trace: design.sv:69069:9
				reg_rdata_next[11] = intrpt_lvl_high_status_intrpt_lvl_high_status_11_qs;
				// Trace: design.sv:69070:9
				reg_rdata_next[12] = intrpt_lvl_high_status_intrpt_lvl_high_status_12_qs;
				// Trace: design.sv:69071:9
				reg_rdata_next[13] = intrpt_lvl_high_status_intrpt_lvl_high_status_13_qs;
				// Trace: design.sv:69072:9
				reg_rdata_next[14] = intrpt_lvl_high_status_intrpt_lvl_high_status_14_qs;
				// Trace: design.sv:69073:9
				reg_rdata_next[15] = intrpt_lvl_high_status_intrpt_lvl_high_status_15_qs;
				// Trace: design.sv:69074:9
				reg_rdata_next[16] = intrpt_lvl_high_status_intrpt_lvl_high_status_16_qs;
				// Trace: design.sv:69075:9
				reg_rdata_next[17] = intrpt_lvl_high_status_intrpt_lvl_high_status_17_qs;
				// Trace: design.sv:69076:9
				reg_rdata_next[18] = intrpt_lvl_high_status_intrpt_lvl_high_status_18_qs;
				// Trace: design.sv:69077:9
				reg_rdata_next[19] = intrpt_lvl_high_status_intrpt_lvl_high_status_19_qs;
				// Trace: design.sv:69078:9
				reg_rdata_next[20] = intrpt_lvl_high_status_intrpt_lvl_high_status_20_qs;
				// Trace: design.sv:69079:9
				reg_rdata_next[21] = intrpt_lvl_high_status_intrpt_lvl_high_status_21_qs;
				// Trace: design.sv:69080:9
				reg_rdata_next[22] = intrpt_lvl_high_status_intrpt_lvl_high_status_22_qs;
				// Trace: design.sv:69081:9
				reg_rdata_next[23] = intrpt_lvl_high_status_intrpt_lvl_high_status_23_qs;
				// Trace: design.sv:69082:9
				reg_rdata_next[24] = intrpt_lvl_high_status_intrpt_lvl_high_status_24_qs;
				// Trace: design.sv:69083:9
				reg_rdata_next[25] = intrpt_lvl_high_status_intrpt_lvl_high_status_25_qs;
				// Trace: design.sv:69084:9
				reg_rdata_next[26] = intrpt_lvl_high_status_intrpt_lvl_high_status_26_qs;
				// Trace: design.sv:69085:9
				reg_rdata_next[27] = intrpt_lvl_high_status_intrpt_lvl_high_status_27_qs;
				// Trace: design.sv:69086:9
				reg_rdata_next[28] = intrpt_lvl_high_status_intrpt_lvl_high_status_28_qs;
				// Trace: design.sv:69087:9
				reg_rdata_next[29] = intrpt_lvl_high_status_intrpt_lvl_high_status_29_qs;
				// Trace: design.sv:69088:9
				reg_rdata_next[30] = intrpt_lvl_high_status_intrpt_lvl_high_status_30_qs;
				// Trace: design.sv:69089:9
				reg_rdata_next[31] = intrpt_lvl_high_status_intrpt_lvl_high_status_31_qs;
			end
			addr_hit[18]: begin
				// Trace: design.sv:69093:9
				reg_rdata_next[0] = intrpt_lvl_low_status_intrpt_lvl_low_status_0_qs;
				// Trace: design.sv:69094:9
				reg_rdata_next[1] = intrpt_lvl_low_status_intrpt_lvl_low_status_1_qs;
				// Trace: design.sv:69095:9
				reg_rdata_next[2] = intrpt_lvl_low_status_intrpt_lvl_low_status_2_qs;
				// Trace: design.sv:69096:9
				reg_rdata_next[3] = intrpt_lvl_low_status_intrpt_lvl_low_status_3_qs;
				// Trace: design.sv:69097:9
				reg_rdata_next[4] = intrpt_lvl_low_status_intrpt_lvl_low_status_4_qs;
				// Trace: design.sv:69098:9
				reg_rdata_next[5] = intrpt_lvl_low_status_intrpt_lvl_low_status_5_qs;
				// Trace: design.sv:69099:9
				reg_rdata_next[6] = intrpt_lvl_low_status_intrpt_lvl_low_status_6_qs;
				// Trace: design.sv:69100:9
				reg_rdata_next[7] = intrpt_lvl_low_status_intrpt_lvl_low_status_7_qs;
				// Trace: design.sv:69101:9
				reg_rdata_next[8] = intrpt_lvl_low_status_intrpt_lvl_low_status_8_qs;
				// Trace: design.sv:69102:9
				reg_rdata_next[9] = intrpt_lvl_low_status_intrpt_lvl_low_status_9_qs;
				// Trace: design.sv:69103:9
				reg_rdata_next[10] = intrpt_lvl_low_status_intrpt_lvl_low_status_10_qs;
				// Trace: design.sv:69104:9
				reg_rdata_next[11] = intrpt_lvl_low_status_intrpt_lvl_low_status_11_qs;
				// Trace: design.sv:69105:9
				reg_rdata_next[12] = intrpt_lvl_low_status_intrpt_lvl_low_status_12_qs;
				// Trace: design.sv:69106:9
				reg_rdata_next[13] = intrpt_lvl_low_status_intrpt_lvl_low_status_13_qs;
				// Trace: design.sv:69107:9
				reg_rdata_next[14] = intrpt_lvl_low_status_intrpt_lvl_low_status_14_qs;
				// Trace: design.sv:69108:9
				reg_rdata_next[15] = intrpt_lvl_low_status_intrpt_lvl_low_status_15_qs;
				// Trace: design.sv:69109:9
				reg_rdata_next[16] = intrpt_lvl_low_status_intrpt_lvl_low_status_16_qs;
				// Trace: design.sv:69110:9
				reg_rdata_next[17] = intrpt_lvl_low_status_intrpt_lvl_low_status_17_qs;
				// Trace: design.sv:69111:9
				reg_rdata_next[18] = intrpt_lvl_low_status_intrpt_lvl_low_status_18_qs;
				// Trace: design.sv:69112:9
				reg_rdata_next[19] = intrpt_lvl_low_status_intrpt_lvl_low_status_19_qs;
				// Trace: design.sv:69113:9
				reg_rdata_next[20] = intrpt_lvl_low_status_intrpt_lvl_low_status_20_qs;
				// Trace: design.sv:69114:9
				reg_rdata_next[21] = intrpt_lvl_low_status_intrpt_lvl_low_status_21_qs;
				// Trace: design.sv:69115:9
				reg_rdata_next[22] = intrpt_lvl_low_status_intrpt_lvl_low_status_22_qs;
				// Trace: design.sv:69116:9
				reg_rdata_next[23] = intrpt_lvl_low_status_intrpt_lvl_low_status_23_qs;
				// Trace: design.sv:69117:9
				reg_rdata_next[24] = intrpt_lvl_low_status_intrpt_lvl_low_status_24_qs;
				// Trace: design.sv:69118:9
				reg_rdata_next[25] = intrpt_lvl_low_status_intrpt_lvl_low_status_25_qs;
				// Trace: design.sv:69119:9
				reg_rdata_next[26] = intrpt_lvl_low_status_intrpt_lvl_low_status_26_qs;
				// Trace: design.sv:69120:9
				reg_rdata_next[27] = intrpt_lvl_low_status_intrpt_lvl_low_status_27_qs;
				// Trace: design.sv:69121:9
				reg_rdata_next[28] = intrpt_lvl_low_status_intrpt_lvl_low_status_28_qs;
				// Trace: design.sv:69122:9
				reg_rdata_next[29] = intrpt_lvl_low_status_intrpt_lvl_low_status_29_qs;
				// Trace: design.sv:69123:9
				reg_rdata_next[30] = intrpt_lvl_low_status_intrpt_lvl_low_status_30_qs;
				// Trace: design.sv:69124:9
				reg_rdata_next[31] = intrpt_lvl_low_status_intrpt_lvl_low_status_31_qs;
			end
			default:
				// Trace: design.sv:69128:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:69137:3
	wire unused_wdata;
	// Trace: design.sv:69138:3
	wire unused_be;
	// Trace: design.sv:69139:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:69140:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module gpio_B7E66 (
	clk_i,
	rst_ni,
	gpio_in,
	gpio_out,
	gpio_tx_en_o,
	gpio_in_sync_o,
	global_interrupt_o,
	pin_level_interrupts_o,
	reg_req_i,
	reg_rsp_o
);
	reg _sv2v_0;
	// Trace: design.sv:69181:13
	parameter [31:0] DATA_WIDTH = 32;
	// Trace: design.sv:69183:18
	// removed localparam type reg_req_t
	// Trace: design.sv:69185:18
	// removed localparam type reg_rsp_t
	// Trace: design.sv:69190:14
	localparam signed [31:0] gpio_reg_pkg_GPIOCount = 32;
	localparam [31:0] NrGPIOs = gpio_reg_pkg_GPIOCount;
	// Trace: design.sv:69194:3
	input wire clk_i;
	// Trace: design.sv:69196:3
	input wire rst_ni;
	// Trace: design.sv:69198:3
	input wire [31:0] gpio_in;
	// Trace: design.sv:69200:3
	output wire [31:0] gpio_out;
	// Trace: design.sv:69203:3
	output reg [31:0] gpio_tx_en_o;
	// Trace: design.sv:69206:3
	output wire [31:0] gpio_in_sync_o;
	// Trace: design.sv:69209:3
	output wire global_interrupt_o;
	// Trace: design.sv:69210:3
	output wire [31:0] pin_level_interrupts_o;
	// Trace: design.sv:69212:3
	input wire [69:0] reg_req_i;
	// Trace: design.sv:69214:3
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:69217:3
	localparam [9:0] HW_VERSION = 2;
	// Trace: design.sv:69219:3
	// removed import gpio_reg_pkg::*;
	// Trace: design.sv:69222:3
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_cfg_reg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_clear_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_mode_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_out_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_set_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_gpio_toggle_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_fall_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_fall_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_lvl_high_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_lvl_high_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_lvl_low_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_lvl_low_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_rise_en_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_rise_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_intrpt_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_reg2hw_t
	wire [642:0] s_reg2hw;
	// Trace: design.sv:69223:3
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_gpio_in_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_gpio_out_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_info_reg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_fall_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_lvl_high_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_lvl_low_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_rise_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_intrpt_status_mreg_t
	// removed localparam type gpio_reg_pkg_gpio_hw2reg_t
	reg [403:0] s_hw2reg;
	// Trace: design.sv:69226:3
	wire [31:0] s_gpio_in_sync;
	// Trace: design.sv:69230:3
	wire [31:0] s_gpio_rise_edge;
	// Trace: design.sv:69231:3
	wire [31:0] s_gpio_rise_intrpt_mask;
	// Trace: design.sv:69232:3
	wire [31:0] s_gpio_fall_edge;
	// Trace: design.sv:69233:3
	wire [31:0] s_gpio_fall_intrpt_mask;
	// Trace: design.sv:69236:3
	wire [31:0] s_gpio_high_intrpt_mask;
	// Trace: design.sv:69237:3
	wire [31:0] s_gpio_low_intrpt_mask;
	// Trace: design.sv:69239:3
	wire [31:0] s_gpio_rise_intrpt;
	// Trace: design.sv:69240:3
	wire [31:0] s_gpio_fall_intrpt;
	// Trace: design.sv:69241:3
	wire [31:0] s_gpio_high_intrpt;
	// Trace: design.sv:69242:3
	wire [31:0] s_gpio_low_intrpt;
	// Trace: design.sv:69245:3
	wire [31:0] interrupts_edges;
	// Trace: design.sv:69246:3
	wire [31:0] interrupts_pending;
	// Trace: design.sv:69249:3
	gpio_reg_top_04165 i_reg_file(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(reg_req_i),
		.reg_rsp_o(reg_rsp_o),
		.reg2hw(s_reg2hw),
		.hw2reg(s_hw2reg),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:69263:3
	wire [10:1] sv2v_tmp_854C4;
	assign sv2v_tmp_854C4 = HW_VERSION;
	always @(*) s_hw2reg[393-:10] = sv2v_tmp_854C4;
	// Trace: design.sv:69264:3
	wire [10:1] sv2v_tmp_A9BF5;
	assign sv2v_tmp_A9BF5 = NrGPIOs[9:0];
	always @(*) s_hw2reg[403-:10] = sv2v_tmp_A9BF5;
	// Trace: design.sv:69267:3
	assign s_gpio_rise_intrpt = s_gpio_rise_edge & s_gpio_rise_intrpt_mask;
	// Trace: design.sv:69268:3
	assign s_gpio_fall_intrpt = s_gpio_fall_edge & s_gpio_fall_intrpt_mask;
	// Trace: design.sv:69269:3
	assign s_gpio_high_intrpt = s_gpio_in_sync & s_gpio_high_intrpt_mask;
	// Trace: design.sv:69270:3
	assign s_gpio_low_intrpt = ~s_gpio_in_sync & s_gpio_low_intrpt_mask;
	// Trace: design.sv:69274:3
	assign interrupts_edges = ((s_gpio_rise_intrpt | s_gpio_fall_intrpt) | s_gpio_high_intrpt) | s_gpio_low_intrpt;
	// Trace: design.sv:69277:3
	assign interrupts_pending = ((s_reg2hw[127-:32] | s_reg2hw[95-:32]) | s_reg2hw[63-:32]) | s_reg2hw[31-:32];
	// Trace: design.sv:69280:3
	assign global_interrupt_o = (s_reg2hw[642] ? |interrupts_pending : |interrupts_edges);
	// Trace: design.sv:69281:3
	assign pin_level_interrupts_o = (s_reg2hw[641] ? interrupts_pending : interrupts_edges);
	// Trace: design.sv:69284:3
	assign gpio_in_sync_o = s_gpio_in_sync;
	// Trace: design.sv:69287:3
	genvar _gv_gpio_idx_1;
	generate
		for (_gv_gpio_idx_1 = 0; _gv_gpio_idx_1 < NrGPIOs; _gv_gpio_idx_1 = _gv_gpio_idx_1 + 1) begin : gen_gpios
			localparam gpio_idx = _gv_gpio_idx_1;
			// Trace: design.sv:69289:7
			gpio_input_stage #(.NrSyncStages(2)) i_sync_gpio_input(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.en_i(s_reg2hw[544 + gpio_idx] && (s_reg2hw[576 + ((gpio_idx * 2) + 1)-:2] == 0)),
				.serial_i(gpio_in[gpio_idx]),
				.r_edge_o(s_gpio_rise_edge[gpio_idx]),
				.f_edge_o(s_gpio_fall_edge[gpio_idx]),
				.serial_o(s_gpio_in_sync[gpio_idx])
			);
			// Trace: design.sv:69302:7
			wire [1:1] sv2v_tmp_9F468;
			assign sv2v_tmp_9F468 = s_gpio_in_sync[gpio_idx];
			always @(*) s_hw2reg[352 + gpio_idx] = sv2v_tmp_9F468;
			// Trace: design.sv:69305:7
			assign gpio_out[gpio_idx] = s_reg2hw[512 + gpio_idx];
			// Trace: design.sv:69307:7
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:69308:64
				case (s_reg2hw[576 + (gpio_idx * 2)+:2])
					2'b00:
						// Trace: design.sv:69311:13
						gpio_tx_en_o[gpio_idx] = 1'b0;
					2'b01:
						// Trace: design.sv:69314:13
						gpio_tx_en_o[gpio_idx] = 1'b1;
					2'b10:
						// Trace: design.sv:69317:13
						gpio_tx_en_o[gpio_idx] = s_reg2hw[512 + gpio_idx];
					2'b11:
						// Trace: design.sv:69320:13
						gpio_tx_en_o[gpio_idx] = ~s_reg2hw[512 + gpio_idx];
					default:
						// Trace: design.sv:69323:13
						gpio_tx_en_o[gpio_idx] = 1'b0;
				endcase
			end
			// Trace: design.sv:69329:7
			assign s_gpio_rise_intrpt_mask[gpio_idx] = s_reg2hw[288 + gpio_idx];
			// Trace: design.sv:69330:7
			assign s_gpio_fall_intrpt_mask[gpio_idx] = s_reg2hw[256 + gpio_idx];
			// Trace: design.sv:69331:7
			assign s_gpio_high_intrpt_mask[gpio_idx] = s_reg2hw[224 + gpio_idx];
			// Trace: design.sv:69332:7
			assign s_gpio_low_intrpt_mask[gpio_idx] = s_reg2hw[192 + gpio_idx];
			// Trace: design.sv:69335:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:69336:7
				s_hw2reg[288 + ((gpio_idx * 2) + 1)] = s_reg2hw[512 + gpio_idx];
				// Trace: design.sv:69337:7
				s_hw2reg[288 + (gpio_idx * 2)] = 1'b0;
				// Trace: design.sv:69338:7
				if (s_reg2hw[448 + (gpio_idx * 2)] && s_reg2hw[448 + ((gpio_idx * 2) + 1)]) begin
					// Trace: design.sv:69339:99
					// Trace: design.sv:69340:9
					s_hw2reg[288 + ((gpio_idx * 2) + 1)] = 1'b1;
					// Trace: design.sv:69341:9
					s_hw2reg[288 + (gpio_idx * 2)] = 1'b1;
				end
				else if (s_reg2hw[384 + (gpio_idx * 2)] && s_reg2hw[384 + ((gpio_idx * 2) + 1)]) begin
					// Trace: design.sv:69343:103
					// Trace: design.sv:69344:9
					s_hw2reg[288 + ((gpio_idx * 2) + 1)] = 1'b0;
					// Trace: design.sv:69345:9
					s_hw2reg[288 + (gpio_idx * 2)] = 1'b1;
				end
				else if (s_reg2hw[320 + (gpio_idx * 2)] && s_reg2hw[320 + ((gpio_idx * 2) + 1)]) begin
					// Trace: design.sv:69347:105
					// Trace: design.sv:69348:9
					s_hw2reg[288 + ((gpio_idx * 2) + 1)] = ~s_reg2hw[512 + gpio_idx];
					// Trace: design.sv:69349:9
					s_hw2reg[288 + (gpio_idx * 2)] = 1'b1;
				end
				else begin
					// Trace: design.sv:69351:9
					s_hw2reg[288 + ((gpio_idx * 2) + 1)] = s_reg2hw[512 + gpio_idx];
					// Trace: design.sv:69352:9
					s_hw2reg[288 + (gpio_idx * 2)] = 1'b0;
				end
			end
			// Trace: design.sv:69357:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:69358:107
				if (s_reg2hw[128 + (gpio_idx * 2)] & (s_reg2hw[128 + ((gpio_idx * 2) + 1)] == 1)) begin
					// Trace: design.sv:69362:9
					s_hw2reg[192 + ((gpio_idx * 2) + 1)] = 1'sb0;
					// Trace: design.sv:69363:9
					s_hw2reg[192 + (gpio_idx * 2)] = 1'b1;
					// Trace: design.sv:69364:9
					s_hw2reg[128 + ((gpio_idx * 2) + 1)] = 1'sb0;
					// Trace: design.sv:69365:9
					s_hw2reg[128 + (gpio_idx * 2)] = 1'b1;
					// Trace: design.sv:69366:9
					s_hw2reg[64 + ((gpio_idx * 2) + 1)] = 1'sb0;
					// Trace: design.sv:69367:9
					s_hw2reg[64 + (gpio_idx * 2)] = 1'b1;
					// Trace: design.sv:69368:9
					s_hw2reg[0 + ((gpio_idx * 2) + 1)] = 1'sb0;
					// Trace: design.sv:69369:9
					s_hw2reg[0 + (gpio_idx * 2)] = 1'b1;
				end
				else begin
					// Trace: design.sv:69374:9
					s_hw2reg[192 + ((gpio_idx * 2) + 1)] = s_gpio_rise_intrpt[gpio_idx] | s_reg2hw[96 + gpio_idx];
					// Trace: design.sv:69375:9
					s_hw2reg[192 + (gpio_idx * 2)] = |s_gpio_rise_intrpt[gpio_idx];
					// Trace: design.sv:69376:9
					s_hw2reg[128 + ((gpio_idx * 2) + 1)] = s_gpio_fall_intrpt[gpio_idx] | s_reg2hw[64 + gpio_idx];
					// Trace: design.sv:69377:9
					s_hw2reg[128 + (gpio_idx * 2)] = |s_gpio_fall_intrpt[gpio_idx];
					// Trace: design.sv:69378:9
					s_hw2reg[64 + ((gpio_idx * 2) + 1)] = s_gpio_high_intrpt[gpio_idx] | s_reg2hw[32 + gpio_idx];
					// Trace: design.sv:69379:9
					s_hw2reg[64 + (gpio_idx * 2)] = |s_gpio_high_intrpt[gpio_idx];
					// Trace: design.sv:69380:9
					s_hw2reg[0 + ((gpio_idx * 2) + 1)] = s_gpio_low_intrpt[gpio_idx] | s_reg2hw[0 + gpio_idx];
					// Trace: design.sv:69381:9
					s_hw2reg[0 + (gpio_idx * 2)] = |s_gpio_low_intrpt[gpio_idx];
				end
			end
			// Trace: design.sv:69384:5
			wire [1:1] sv2v_tmp_8DE20;
			assign sv2v_tmp_8DE20 = interrupts_pending[gpio_idx];
			always @(*) s_hw2reg[256 + gpio_idx] = sv2v_tmp_8DE20;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
// removed module with interface ports: gpio_intf
module gpio_input_stage (
	clk_i,
	rst_ni,
	en_i,
	serial_i,
	r_edge_o,
	f_edge_o,
	serial_o
);
	// Trace: design.sv:69472:13
	parameter NrSyncStages = 2;
	// Trace: design.sv:69474:4
	input wire clk_i;
	// Trace: design.sv:69475:4
	input wire rst_ni;
	// Trace: design.sv:69476:4
	input wire en_i;
	// Trace: design.sv:69477:4
	input wire serial_i;
	// Trace: design.sv:69478:4
	output wire r_edge_o;
	// Trace: design.sv:69479:4
	output wire f_edge_o;
	// Trace: design.sv:69480:4
	output wire serial_o;
	// Trace: design.sv:69483:3
	wire clk;
	// Trace: design.sv:69484:3
	wire serial;
	reg serial_q;
	// Trace: design.sv:69486:3
	assign serial_o = serial_q;
	// Trace: design.sv:69487:3
	assign f_edge_o = ~serial & serial_q;
	// Trace: design.sv:69488:3
	assign r_edge_o = serial & ~serial_q;
	// Trace: design.sv:69490:3
	tc_clk_gating #(.IS_FUNCTIONAL(0)) i_clk_gate(
		.clk_i(clk_i),
		.en_i(en_i),
		.test_en_i(1'b0),
		.clk_o(clk)
	);
	// Trace: design.sv:69500:3
	sync #(.STAGES(NrSyncStages)) i_sync(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.serial_i(serial_i),
		.serial_o(serial)
	);
	// Trace: design.sv:69509:3
	always @(posedge clk or negedge rst_ni)
		// Trace: design.sv:69510:5
		if (!rst_ni)
			// Trace: design.sv:69511:7
			serial_q <= 1'b0;
		else
			// Trace: design.sv:69513:7
			serial_q <= serial;
endmodule
module boot_rom (
	reg_req_i,
	reg_rsp_o
);
	reg _sv2v_0;
	// removed import reg_pkg::*;
	// Trace: design.sv:69538:5
	// removed localparam type reg_pkg_reg_req_t
	input wire [69:0] reg_req_i;
	// Trace: design.sv:69539:5
	// removed localparam type reg_pkg_reg_rsp_t
	output reg [33:0] reg_rsp_o;
	// Trace: design.sv:69541:3
	// removed import core_v_mini_mcu_pkg::*;
	// Trace: design.sv:69543:3
	localparam [31:0] RomSize = 59;
	// Trace: design.sv:69545:3
	wire [1887:0] mem;
	// Trace: design.sv:69546:3
	assign mem = 1888'h96024990200005b7f2e9f0068693ff7493e3fec49be304910114a0230285a88302048613dfed8b8583d149dc10048b93fe07dfe349dc00010355a2230ff40a930800043700db46630ff40a930900043710000b13448140000693fe07dfe349dc0001d1d8070d11000737fe075fe349d80001d5d8470dfe075fe349d8d1d8070d10000737d5d80ab00713c99800876713f00777134998d1884501cd9807050fff0737c9988f494998a0000537200205b7958218058593400005b7c1884505200285b7c9110145c5039582498cd17500c5c503e5110085c503200005b7950241c8c1190005c503200405b7;
	// Trace: design.sv:69608:3
	localparam [31:0] core_v_mini_mcu_pkg_BOOTROM_SIZE = 32'h00010000;
	wire [$clog2(32'h00010000) - 3:0] word_addr;
	// Trace: design.sv:69609:3
	wire [5:0] rom_addr;
	// Trace: design.sv:69611:3
	assign word_addr = reg_req_i[31 + $clog2(32'h00010000):34];
	// Trace: design.sv:69612:3
	assign rom_addr = word_addr[5:0];
	// Trace: design.sv:69614:3
	wire [1:1] sv2v_tmp_FC5C0;
	assign sv2v_tmp_FC5C0 = 1'b0;
	always @(*) reg_rsp_o[33] = sv2v_tmp_FC5C0;
	// Trace: design.sv:69615:3
	wire [1:1] sv2v_tmp_6CD20;
	assign sv2v_tmp_6CD20 = 1'b1;
	always @(*) reg_rsp_o[32] = sv2v_tmp_6CD20;
	// Trace: design.sv:69617:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:69618:5
		if (word_addr > 58)
			// Trace: design.sv:69619:7
			reg_rsp_o[31-:32] = 1'sb0;
		else
			// Trace: design.sv:69621:7
			reg_rsp_o[31-:32] = mem[rom_addr * 32+:32];
	end
	initial _sv2v_0 = 0;
endmodule
// removed package "dma_reg_pkg"
module dma_reg_top_A4ADD (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	reg2hw,
	hw2reg,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:69728:20
	// removed localparam type reg_req_t
	// Trace: design.sv:69729:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:69730:15
	parameter signed [31:0] AW = 5;
	// Trace: design.sv:69732:5
	input clk_i;
	// Trace: design.sv:69733:5
	input rst_ni;
	// Trace: design.sv:69734:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:69735:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:69737:5
	// removed localparam type dma_reg_pkg_dma_reg2hw_data_type_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_dma_start_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_dst_ptr_inc_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_ptr_in_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_ptr_out_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_spi_mode_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_src_ptr_inc_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_t
	output wire [164:0] reg2hw;
	// Trace: design.sv:69738:5
	// removed localparam type dma_reg_pkg_dma_hw2reg_dma_start_reg_t
	// removed localparam type dma_reg_pkg_dma_hw2reg_done_reg_t
	// removed localparam type dma_reg_pkg_dma_hw2reg_t
	input wire [65:0] hw2reg;
	// Trace: design.sv:69742:5
	input devmode_i;
	// Trace: design.sv:69745:3
	// removed import dma_reg_pkg::*;
	// Trace: design.sv:69747:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:69748:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:69751:3
	wire reg_we;
	// Trace: design.sv:69752:3
	wire reg_re;
	// Trace: design.sv:69753:3
	wire [AW - 1:0] reg_addr;
	// Trace: design.sv:69754:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:69755:3
	wire [3:0] reg_be;
	// Trace: design.sv:69756:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:69757:3
	wire reg_error;
	// Trace: design.sv:69759:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:69761:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:69764:3
	wire [69:0] reg_intf_req;
	// Trace: design.sv:69765:3
	wire [33:0] reg_intf_rsp;
	// Trace: design.sv:69768:3
	assign reg_intf_req = reg_req_i;
	// Trace: design.sv:69769:3
	assign reg_rsp_o = reg_intf_rsp;
	// Trace: design.sv:69772:3
	assign reg_we = reg_intf_req[69] & reg_intf_req[68];
	// Trace: design.sv:69773:3
	assign reg_re = reg_intf_req[69] & ~reg_intf_req[68];
	// Trace: design.sv:69774:3
	assign reg_addr = reg_intf_req[63-:32];
	// Trace: design.sv:69775:3
	assign reg_wdata = reg_intf_req[31-:32];
	// Trace: design.sv:69776:3
	assign reg_be = reg_intf_req[67-:4];
	// Trace: design.sv:69777:3
	assign reg_intf_rsp[31-:32] = reg_rdata;
	// Trace: design.sv:69778:3
	assign reg_intf_rsp[33] = reg_error;
	// Trace: design.sv:69779:3
	assign reg_intf_rsp[32] = 1'b1;
	// Trace: design.sv:69781:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:69782:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:69788:3
	wire [31:0] ptr_in_qs;
	// Trace: design.sv:69789:3
	wire [31:0] ptr_in_wd;
	// Trace: design.sv:69790:3
	wire ptr_in_we;
	// Trace: design.sv:69791:3
	wire [31:0] ptr_out_qs;
	// Trace: design.sv:69792:3
	wire [31:0] ptr_out_wd;
	// Trace: design.sv:69793:3
	wire ptr_out_we;
	// Trace: design.sv:69794:3
	wire [31:0] dma_start_qs;
	// Trace: design.sv:69795:3
	wire [31:0] dma_start_wd;
	// Trace: design.sv:69796:3
	wire dma_start_we;
	// Trace: design.sv:69797:3
	wire [31:0] done_qs;
	// Trace: design.sv:69798:3
	wire [31:0] src_ptr_inc_qs;
	// Trace: design.sv:69799:3
	wire [31:0] src_ptr_inc_wd;
	// Trace: design.sv:69800:3
	wire src_ptr_inc_we;
	// Trace: design.sv:69801:3
	wire [31:0] dst_ptr_inc_qs;
	// Trace: design.sv:69802:3
	wire [31:0] dst_ptr_inc_wd;
	// Trace: design.sv:69803:3
	wire dst_ptr_inc_we;
	// Trace: design.sv:69804:3
	wire [2:0] spi_mode_qs;
	// Trace: design.sv:69805:3
	wire [2:0] spi_mode_wd;
	// Trace: design.sv:69806:3
	wire spi_mode_we;
	// Trace: design.sv:69807:3
	wire [1:0] data_type_qs;
	// Trace: design.sv:69808:3
	wire [1:0] data_type_wd;
	// Trace: design.sv:69809:3
	wire data_type_we;
	// Trace: design.sv:69814:3
	localparam signed [31:0] sv2v_uu_u_ptr_in_DW = 32;
	// removed localparam type sv2v_uu_u_ptr_in_d
	localparam [31:0] sv2v_uu_u_ptr_in_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_ptr_in(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ptr_in_we),
		.wd(ptr_in_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ptr_in_ext_d_0),
		.qe(),
		.q(reg2hw[164-:32]),
		.qs(ptr_in_qs)
	);
	// Trace: design.sv:69841:3
	localparam signed [31:0] sv2v_uu_u_ptr_out_DW = 32;
	// removed localparam type sv2v_uu_u_ptr_out_d
	localparam [31:0] sv2v_uu_u_ptr_out_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_ptr_out(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ptr_out_we),
		.wd(ptr_out_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ptr_out_ext_d_0),
		.qe(),
		.q(reg2hw[132-:32]),
		.qs(ptr_out_qs)
	);
	// Trace: design.sv:69868:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_dma_start(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dma_start_we),
		.wd(dma_start_wd),
		.de(hw2reg[33]),
		.d(hw2reg[65-:32]),
		.qe(),
		.q(reg2hw[100-:32]),
		.qs(dma_start_qs)
	);
	// Trace: design.sv:69895:3
	localparam signed [31:0] sv2v_uu_u_done_DW = 32;
	// removed localparam type sv2v_uu_u_done_wd
	localparam [31:0] sv2v_uu_u_done_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RO"),
		.RESVAL(32'h00000001)
	) u_done(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_done_ext_wd_0),
		.de(hw2reg[0]),
		.d(hw2reg[32-:32]),
		.qe(),
		.q(),
		.qs(done_qs)
	);
	// Trace: design.sv:69921:3
	localparam signed [31:0] sv2v_uu_u_src_ptr_inc_DW = 32;
	// removed localparam type sv2v_uu_u_src_ptr_inc_d
	localparam [31:0] sv2v_uu_u_src_ptr_inc_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000004)
	) u_src_ptr_inc(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(src_ptr_inc_we),
		.wd(src_ptr_inc_wd),
		.de(1'b0),
		.d(sv2v_uu_u_src_ptr_inc_ext_d_0),
		.qe(),
		.q(reg2hw[68-:32]),
		.qs(src_ptr_inc_qs)
	);
	// Trace: design.sv:69948:3
	localparam signed [31:0] sv2v_uu_u_dst_ptr_inc_DW = 32;
	// removed localparam type sv2v_uu_u_dst_ptr_inc_d
	localparam [31:0] sv2v_uu_u_dst_ptr_inc_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000004)
	) u_dst_ptr_inc(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dst_ptr_inc_we),
		.wd(dst_ptr_inc_wd),
		.de(1'b0),
		.d(sv2v_uu_u_dst_ptr_inc_ext_d_0),
		.qe(),
		.q(reg2hw[36-:32]),
		.qs(dst_ptr_inc_qs)
	);
	// Trace: design.sv:69975:3
	localparam signed [31:0] sv2v_uu_u_spi_mode_DW = 3;
	// removed localparam type sv2v_uu_u_spi_mode_d
	localparam [2:0] sv2v_uu_u_spi_mode_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_spi_mode(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(spi_mode_we),
		.wd(spi_mode_wd),
		.de(1'b0),
		.d(sv2v_uu_u_spi_mode_ext_d_0),
		.qe(),
		.q(reg2hw[4-:3]),
		.qs(spi_mode_qs)
	);
	// Trace: design.sv:70002:3
	localparam signed [31:0] sv2v_uu_u_data_type_DW = 2;
	// removed localparam type sv2v_uu_u_data_type_d
	localparam [1:0] sv2v_uu_u_data_type_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_data_type(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(data_type_we),
		.wd(data_type_wd),
		.de(1'b0),
		.d(sv2v_uu_u_data_type_ext_d_0),
		.qe(),
		.q(reg2hw[1-:2]),
		.qs(data_type_qs)
	);
	// Trace: design.sv:70029:3
	reg [7:0] addr_hit;
	// Trace: design.sv:70030:3
	localparam signed [31:0] dma_reg_pkg_BlockAw = 5;
	localparam [4:0] dma_reg_pkg_DMA_DATA_TYPE_OFFSET = 5'h1c;
	localparam [4:0] dma_reg_pkg_DMA_DMA_START_OFFSET = 5'h08;
	localparam [4:0] dma_reg_pkg_DMA_DONE_OFFSET = 5'h0c;
	localparam [4:0] dma_reg_pkg_DMA_DST_PTR_INC_OFFSET = 5'h14;
	localparam [4:0] dma_reg_pkg_DMA_PTR_IN_OFFSET = 5'h00;
	localparam [4:0] dma_reg_pkg_DMA_PTR_OUT_OFFSET = 5'h04;
	localparam [4:0] dma_reg_pkg_DMA_SPI_MODE_OFFSET = 5'h18;
	localparam [4:0] dma_reg_pkg_DMA_SRC_PTR_INC_OFFSET = 5'h10;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:70031:5
		addr_hit = 1'sb0;
		// Trace: design.sv:70032:5
		addr_hit[0] = reg_addr == dma_reg_pkg_DMA_PTR_IN_OFFSET;
		// Trace: design.sv:70033:5
		addr_hit[1] = reg_addr == dma_reg_pkg_DMA_PTR_OUT_OFFSET;
		// Trace: design.sv:70034:5
		addr_hit[2] = reg_addr == dma_reg_pkg_DMA_DMA_START_OFFSET;
		// Trace: design.sv:70035:5
		addr_hit[3] = reg_addr == dma_reg_pkg_DMA_DONE_OFFSET;
		// Trace: design.sv:70036:5
		addr_hit[4] = reg_addr == dma_reg_pkg_DMA_SRC_PTR_INC_OFFSET;
		// Trace: design.sv:70037:5
		addr_hit[5] = reg_addr == dma_reg_pkg_DMA_DST_PTR_INC_OFFSET;
		// Trace: design.sv:70038:5
		addr_hit[6] = reg_addr == dma_reg_pkg_DMA_SPI_MODE_OFFSET;
		// Trace: design.sv:70039:5
		addr_hit[7] = reg_addr == dma_reg_pkg_DMA_DATA_TYPE_OFFSET;
	end
	// Trace: design.sv:70042:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:70045:3
	localparam [31:0] dma_reg_pkg_DMA_PERMIT = 32'b11111111111111111111111100010001;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:70046:5
		wr_err = reg_we & ((((((((addr_hit[0] & |(dma_reg_pkg_DMA_PERMIT[28+:4] & ~reg_be)) | (addr_hit[1] & |(dma_reg_pkg_DMA_PERMIT[24+:4] & ~reg_be))) | (addr_hit[2] & |(dma_reg_pkg_DMA_PERMIT[20+:4] & ~reg_be))) | (addr_hit[3] & |(dma_reg_pkg_DMA_PERMIT[16+:4] & ~reg_be))) | (addr_hit[4] & |(dma_reg_pkg_DMA_PERMIT[12+:4] & ~reg_be))) | (addr_hit[5] & |(dma_reg_pkg_DMA_PERMIT[8+:4] & ~reg_be))) | (addr_hit[6] & |(dma_reg_pkg_DMA_PERMIT[4+:4] & ~reg_be))) | (addr_hit[7] & |(dma_reg_pkg_DMA_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:70057:3
	assign ptr_in_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:70058:3
	assign ptr_in_wd = reg_wdata[31:0];
	// Trace: design.sv:70060:3
	assign ptr_out_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:70061:3
	assign ptr_out_wd = reg_wdata[31:0];
	// Trace: design.sv:70063:3
	assign dma_start_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:70064:3
	assign dma_start_wd = reg_wdata[31:0];
	// Trace: design.sv:70066:3
	assign src_ptr_inc_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:70067:3
	assign src_ptr_inc_wd = reg_wdata[31:0];
	// Trace: design.sv:70069:3
	assign dst_ptr_inc_we = (addr_hit[5] & reg_we) & !reg_error;
	// Trace: design.sv:70070:3
	assign dst_ptr_inc_wd = reg_wdata[31:0];
	// Trace: design.sv:70072:3
	assign spi_mode_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:70073:3
	assign spi_mode_wd = reg_wdata[2:0];
	// Trace: design.sv:70075:3
	assign data_type_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:70076:3
	assign data_type_wd = reg_wdata[1:0];
	// Trace: design.sv:70079:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:70080:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:70081:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]:
				// Trace: design.sv:70083:9
				reg_rdata_next[31:0] = ptr_in_qs;
			addr_hit[1]:
				// Trace: design.sv:70087:9
				reg_rdata_next[31:0] = ptr_out_qs;
			addr_hit[2]:
				// Trace: design.sv:70091:9
				reg_rdata_next[31:0] = dma_start_qs;
			addr_hit[3]:
				// Trace: design.sv:70095:9
				reg_rdata_next[31:0] = done_qs;
			addr_hit[4]:
				// Trace: design.sv:70099:9
				reg_rdata_next[31:0] = src_ptr_inc_qs;
			addr_hit[5]:
				// Trace: design.sv:70103:9
				reg_rdata_next[31:0] = dst_ptr_inc_qs;
			addr_hit[6]:
				// Trace: design.sv:70107:9
				reg_rdata_next[2:0] = spi_mode_qs;
			addr_hit[7]:
				// Trace: design.sv:70111:9
				reg_rdata_next[1:0] = data_type_qs;
			default:
				// Trace: design.sv:70115:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:70124:3
	wire unused_wdata;
	// Trace: design.sv:70125:3
	wire unused_be;
	// Trace: design.sv:70126:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:70127:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module dma_689DF (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	dma_master0_ch0_req_o,
	dma_master0_ch0_resp_i,
	dma_master1_ch0_req_o,
	dma_master1_ch0_resp_i,
	spi_rx_valid_i,
	spi_tx_ready_i,
	spi_flash_rx_valid_i,
	spi_flash_tx_ready_i,
	dma_intr_o
);
	reg _sv2v_0;
	// Trace: design.sv:70140:15
	parameter [31:0] FIFO_DEPTH = 4;
	// Trace: design.sv:70141:20
	// removed localparam type reg_req_t
	// Trace: design.sv:70142:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:70143:20
	// removed localparam type obi_req_t
	// Trace: design.sv:70144:20
	// removed localparam type obi_resp_t
	// Trace: design.sv:70146:5
	input wire clk_i;
	// Trace: design.sv:70147:5
	input wire rst_ni;
	// Trace: design.sv:70149:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:70150:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:70152:5
	output wire [69:0] dma_master0_ch0_req_o;
	// Trace: design.sv:70153:5
	input wire [33:0] dma_master0_ch0_resp_i;
	// Trace: design.sv:70155:5
	output wire [69:0] dma_master1_ch0_req_o;
	// Trace: design.sv:70156:5
	input wire [33:0] dma_master1_ch0_resp_i;
	// Trace: design.sv:70158:5
	input wire spi_rx_valid_i;
	// Trace: design.sv:70159:5
	input wire spi_tx_ready_i;
	// Trace: design.sv:70160:5
	input wire spi_flash_rx_valid_i;
	// Trace: design.sv:70161:5
	input wire spi_flash_tx_ready_i;
	// Trace: design.sv:70163:5
	output wire dma_intr_o;
	// Trace: design.sv:70166:3
	// removed import dma_reg_pkg::*;
	// Trace: design.sv:70168:3
	localparam [31:0] LastFifoUsage = FIFO_DEPTH - 1;
	// Trace: design.sv:70169:3
	localparam [31:0] Addr_Fifo_Depth = (FIFO_DEPTH > 1 ? $clog2(FIFO_DEPTH) : 1);
	// Trace: design.sv:70171:3
	// removed localparam type dma_reg_pkg_dma_reg2hw_data_type_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_dma_start_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_dst_ptr_inc_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_ptr_in_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_ptr_out_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_spi_mode_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_src_ptr_inc_reg_t
	// removed localparam type dma_reg_pkg_dma_reg2hw_t
	wire [164:0] reg2hw;
	// Trace: design.sv:70172:3
	// removed localparam type dma_reg_pkg_dma_hw2reg_dma_start_reg_t
	// removed localparam type dma_reg_pkg_dma_hw2reg_done_reg_t
	// removed localparam type dma_reg_pkg_dma_hw2reg_t
	wire [65:0] hw2reg;
	// Trace: design.sv:70174:3
	reg [31:0] read_ptr_reg;
	// Trace: design.sv:70175:3
	reg [31:0] read_ptr_valid_reg;
	// Trace: design.sv:70176:3
	reg [31:0] write_ptr_reg;
	// Trace: design.sv:70177:3
	reg [31:0] dma_cnt;
	// Trace: design.sv:70178:3
	reg [31:0] dma_cnt_dec;
	// Trace: design.sv:70179:3
	reg dma_start;
	// Trace: design.sv:70180:3
	reg dma_done;
	// Trace: design.sv:70182:3
	wire [Addr_Fifo_Depth - 1:0] fifo_usage;
	// Trace: design.sv:70183:3
	wire fifo_alm_full;
	// Trace: design.sv:70185:3
	reg data_in_req;
	// Trace: design.sv:70186:3
	reg data_in_we;
	// Trace: design.sv:70187:3
	reg [3:0] data_in_be;
	// Trace: design.sv:70188:3
	reg [31:0] data_in_addr;
	// Trace: design.sv:70189:3
	wire data_in_gnt;
	// Trace: design.sv:70190:3
	wire data_in_rvalid;
	// Trace: design.sv:70191:3
	wire [31:0] data_in_rdata;
	// Trace: design.sv:70193:3
	reg data_out_req;
	// Trace: design.sv:70194:3
	reg data_out_we;
	// Trace: design.sv:70195:3
	reg [3:0] data_out_be;
	// Trace: design.sv:70196:3
	reg [31:0] data_out_addr;
	// Trace: design.sv:70197:3
	reg [31:0] data_out_wdata;
	// Trace: design.sv:70198:3
	wire data_out_gnt;
	// Trace: design.sv:70199:3
	wire data_out_rvalid;
	// Trace: design.sv:70200:3
	wire [31:0] data_out_rdata;
	// Trace: design.sv:70202:3
	reg fifo_flush;
	// Trace: design.sv:70203:3
	wire fifo_full;
	// Trace: design.sv:70204:3
	wire fifo_empty;
	// Trace: design.sv:70206:3
	wire [2:0] spi_dma_mode;
	// Trace: design.sv:70207:3
	wire wait_for_rx_spi;
	// Trace: design.sv:70208:3
	wire wait_for_tx_spi;
	// Trace: design.sv:70210:3
	wire [1:0] data_type;
	// Trace: design.sv:70212:3
	reg [31:0] fifo_input;
	// Trace: design.sv:70213:3
	wire [31:0] fifo_output;
	// Trace: design.sv:70215:3
	reg [3:0] byte_enable_out;
	// Trace: design.sv:70217:3
	reg dma_read_fsm_state;
	reg dma_read_fsm_n_state;
	// Trace: design.sv:70223:3
	reg dma_write_fsm_state;
	reg dma_write_fsm_n_state;
	// Trace: design.sv:70229:3
	assign dma_master0_ch0_req_o[69] = data_in_req;
	// Trace: design.sv:70230:3
	assign dma_master0_ch0_req_o[68] = data_in_we;
	// Trace: design.sv:70231:3
	assign dma_master0_ch0_req_o[67-:4] = data_in_be;
	// Trace: design.sv:70232:3
	assign dma_master0_ch0_req_o[63-:32] = data_in_addr;
	// Trace: design.sv:70233:3
	assign dma_master0_ch0_req_o[31-:32] = 32'h00000000;
	// Trace: design.sv:70235:3
	assign data_in_gnt = dma_master0_ch0_resp_i[33];
	// Trace: design.sv:70236:3
	assign data_in_rvalid = dma_master0_ch0_resp_i[32];
	// Trace: design.sv:70237:3
	assign data_in_rdata = dma_master0_ch0_resp_i[31-:32];
	// Trace: design.sv:70239:3
	assign dma_master1_ch0_req_o[69] = data_out_req;
	// Trace: design.sv:70240:3
	assign dma_master1_ch0_req_o[68] = data_out_we;
	// Trace: design.sv:70241:3
	assign dma_master1_ch0_req_o[67-:4] = data_out_be;
	// Trace: design.sv:70242:3
	assign dma_master1_ch0_req_o[63-:32] = data_out_addr;
	// Trace: design.sv:70243:3
	assign dma_master1_ch0_req_o[31-:32] = data_out_wdata;
	// Trace: design.sv:70245:3
	assign data_out_gnt = dma_master1_ch0_resp_i[33];
	// Trace: design.sv:70246:3
	assign data_out_rvalid = dma_master1_ch0_resp_i[32];
	// Trace: design.sv:70247:3
	assign data_out_rdata = dma_master1_ch0_resp_i[31-:32];
	// Trace: design.sv:70249:3
	assign dma_intr_o = dma_done;
	// Trace: design.sv:70250:3
	assign spi_dma_mode = reg2hw[4-:3];
	// Trace: design.sv:70251:3
	assign data_type = reg2hw[1-:2];
	// Trace: design.sv:70253:3
	assign hw2reg[0] = dma_done | dma_start;
	// Trace: design.sv:70254:3
	assign hw2reg[32-:32] = (dma_done == 1'b1 ? 1'b1 : 1'b0);
	// Trace: design.sv:70256:3
	assign hw2reg[33] = dma_start;
	// Trace: design.sv:70257:3
	assign hw2reg[65-:32] = 32'h00000000;
	// Trace: design.sv:70259:3
	assign wait_for_rx_spi = ((spi_dma_mode == 3'h1) && ~spi_rx_valid_i) || ((spi_dma_mode == 3'h3) && ~spi_flash_rx_valid_i);
	// Trace: design.sv:70260:3
	assign wait_for_tx_spi = ((spi_dma_mode == 3'h2) && ~spi_tx_ready_i) || ((spi_dma_mode == 3'h4) && ~spi_flash_tx_ready_i);
	// Trace: design.sv:70262:3
	assign fifo_alm_full = fifo_usage == LastFifoUsage[Addr_Fifo_Depth - 1:0];
	// Trace: design.sv:70265:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_dma_start
		// Trace: design.sv:70266:5
		if (~rst_ni)
			// Trace: design.sv:70267:7
			dma_start <= 1'b0;
		else
			// Trace: design.sv:70269:7
			if (dma_start == 1'b1)
				// Trace: design.sv:70270:9
				dma_start <= 1'b0;
			else
				// Trace: design.sv:70272:9
				dma_start <= |reg2hw[100-:32];
	end
	// Trace: design.sv:70278:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_ptr_in_reg
		// Trace: design.sv:70279:5
		if (~rst_ni)
			// Trace: design.sv:70280:7
			read_ptr_reg <= 1'sb0;
		else
			// Trace: design.sv:70282:7
			if (dma_start == 1'b1)
				// Trace: design.sv:70283:9
				read_ptr_reg <= reg2hw[164-:32];
			else if (data_in_gnt == 1'b1)
				// Trace: design.sv:70285:9
				read_ptr_reg <= read_ptr_reg + reg2hw[68-:32];
	end
	// Trace: design.sv:70291:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_ptr_valid_in_reg
		// Trace: design.sv:70292:5
		if (~rst_ni)
			// Trace: design.sv:70293:7
			read_ptr_valid_reg <= 1'sb0;
		else
			// Trace: design.sv:70295:7
			if (dma_start == 1'b1)
				// Trace: design.sv:70296:9
				read_ptr_valid_reg <= reg2hw[164-:32];
			else if (data_in_rvalid == 1'b1)
				// Trace: design.sv:70298:9
				read_ptr_valid_reg <= read_ptr_valid_reg + reg2hw[68-:32];
	end
	// Trace: design.sv:70304:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_ptr_out_reg
		// Trace: design.sv:70305:5
		if (~rst_ni)
			// Trace: design.sv:70306:7
			write_ptr_reg <= 1'sb0;
		else
			// Trace: design.sv:70308:7
			if (dma_start == 1'b1)
				// Trace: design.sv:70309:9
				write_ptr_reg <= reg2hw[132-:32];
			else if (data_out_gnt == 1'b1)
				// Trace: design.sv:70311:9
				write_ptr_reg <= write_ptr_reg + reg2hw[36-:32];
	end
	// Trace: design.sv:70317:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_dma_cnt_reg
		// Trace: design.sv:70318:5
		if (~rst_ni)
			// Trace: design.sv:70319:7
			dma_cnt <= 1'sb0;
		else
			// Trace: design.sv:70321:7
			if (dma_start == 1'b1)
				// Trace: design.sv:70322:9
				dma_cnt <= reg2hw[100-:32];
			else if (data_in_gnt == 1'b1)
				// Trace: design.sv:70324:9
				dma_cnt <= dma_cnt - dma_cnt_dec;
	end
	// Trace: design.sv:70329:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:70330:5
		case (data_type)
			2'b00:
				// Trace: design.sv:70331:14
				dma_cnt_dec = 32'h00000004;
			2'b01:
				// Trace: design.sv:70332:14
				dma_cnt_dec = 32'h00000002;
			2'b10, 2'b11:
				// Trace: design.sv:70333:21
				dma_cnt_dec = 32'h00000001;
		endcase
	end
	// Trace: design.sv:70337:3
	always @(*) begin : proc_byte_enable_out
		if (_sv2v_0)
			;
		// Trace: design.sv:70338:5
		case (data_type)
			2'b00:
				// Trace: design.sv:70339:14
				byte_enable_out = 4'b1111;
			2'b01:
				// Trace: design.sv:70342:9
				case (write_ptr_reg[1])
					1'b0:
						// Trace: design.sv:70343:17
						byte_enable_out = 4'b0011;
					1'b1:
						// Trace: design.sv:70344:17
						byte_enable_out = 4'b1100;
				endcase
			2'b10, 2'b11:
				// Trace: design.sv:70350:9
				case (write_ptr_reg[1:0])
					2'b00:
						// Trace: design.sv:70351:18
						byte_enable_out = 4'b0001;
					2'b01:
						// Trace: design.sv:70352:18
						byte_enable_out = 4'b0010;
					2'b10:
						// Trace: design.sv:70353:18
						byte_enable_out = 4'b0100;
					2'b11:
						// Trace: design.sv:70354:18
						byte_enable_out = 4'b1000;
				endcase
		endcase
	end
	// Trace: design.sv:70363:3
	always @(*) begin : proc_output_data
		if (_sv2v_0)
			;
		// Trace: design.sv:70365:5
		data_out_wdata[7:0] = fifo_output[7:0];
		// Trace: design.sv:70366:5
		data_out_wdata[15:8] = fifo_output[15:8];
		// Trace: design.sv:70367:5
		data_out_wdata[23:16] = fifo_output[23:16];
		// Trace: design.sv:70368:5
		data_out_wdata[31:24] = fifo_output[31:24];
		// Trace: design.sv:70370:5
		case (write_ptr_reg[1:0])
			2'b00:
				;
			2'b01:
				// Trace: design.sv:70373:14
				data_out_wdata[15:8] = fifo_output[7:0];
			2'b10: begin
				// Trace: design.sv:70376:9
				data_out_wdata[23:16] = fifo_output[7:0];
				// Trace: design.sv:70377:9
				data_out_wdata[31:24] = fifo_output[15:8];
			end
			2'b11:
				// Trace: design.sv:70380:14
				data_out_wdata[31:24] = fifo_output[7:0];
		endcase
	end
	// Trace: design.sv:70385:3
	always @(*) begin : proc_input_data
		if (_sv2v_0)
			;
		// Trace: design.sv:70387:5
		fifo_input[7:0] = data_in_rdata[7:0];
		// Trace: design.sv:70388:5
		fifo_input[15:8] = data_in_rdata[15:8];
		// Trace: design.sv:70389:5
		fifo_input[23:16] = data_in_rdata[23:16];
		// Trace: design.sv:70390:5
		fifo_input[31:24] = data_in_rdata[31:24];
		// Trace: design.sv:70392:5
		case (read_ptr_valid_reg[1:0])
			2'b00:
				;
			2'b01:
				// Trace: design.sv:70395:14
				fifo_input[7:0] = data_in_rdata[15:8];
			2'b10: begin
				// Trace: design.sv:70398:9
				fifo_input[7:0] = data_in_rdata[23:16];
				// Trace: design.sv:70399:9
				fifo_input[15:8] = data_in_rdata[31:24];
			end
			2'b11:
				// Trace: design.sv:70402:14
				fifo_input[7:0] = data_in_rdata[31:24];
		endcase
	end
	// Trace: design.sv:70407:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_fsm_state
		// Trace: design.sv:70408:5
		if (~rst_ni) begin
			// Trace: design.sv:70409:7
			dma_read_fsm_state <= 1'd0;
			// Trace: design.sv:70410:7
			dma_write_fsm_state <= 1'd0;
		end
		else begin
			// Trace: design.sv:70412:7
			dma_read_fsm_state <= dma_read_fsm_n_state;
			// Trace: design.sv:70413:7
			dma_write_fsm_state <= dma_write_fsm_n_state;
		end
	end
	// Trace: design.sv:70418:3
	always @(*) begin : proc_dma_read_fsm_logic
		if (_sv2v_0)
			;
		// Trace: design.sv:70420:5
		dma_read_fsm_n_state = 1'd0;
		// Trace: design.sv:70422:5
		data_in_req = 1'sb0;
		// Trace: design.sv:70423:5
		data_in_we = 1'sb0;
		// Trace: design.sv:70424:5
		data_in_be = 1'sb0;
		// Trace: design.sv:70425:5
		data_in_addr = 1'sb0;
		// Trace: design.sv:70427:5
		fifo_flush = 1'b0;
		// Trace: design.sv:70429:5
		(* full_case, parallel_case *)
		case (dma_read_fsm_state)
			1'd0:
				// Trace: design.sv:70433:9
				if (dma_start == 1'b1) begin
					// Trace: design.sv:70434:11
					dma_read_fsm_n_state = 1'd1;
					// Trace: design.sv:70435:11
					fifo_flush = 1'b1;
				end
				else
					// Trace: design.sv:70437:11
					dma_read_fsm_n_state = 1'd0;
			1'd1:
				// Trace: design.sv:70443:9
				if (|dma_cnt == 1'b0)
					// Trace: design.sv:70444:11
					dma_read_fsm_n_state = 1'd0;
				else begin
					// Trace: design.sv:70446:11
					dma_read_fsm_n_state = 1'd1;
					// Trace: design.sv:70448:11
					if (((fifo_full == 1'b0) && (fifo_alm_full == 1'b0)) && (wait_for_rx_spi == 1'b0)) begin
						// Trace: design.sv:70449:13
						data_in_req = 1'b1;
						// Trace: design.sv:70450:13
						data_in_we = 1'b0;
						// Trace: design.sv:70451:13
						data_in_be = 4'b1111;
						// Trace: design.sv:70452:13
						data_in_addr = read_ptr_reg;
					end
				end
		endcase
	end
	// Trace: design.sv:70460:3
	always @(*) begin : proc_dma_write_fsm_logic
		if (_sv2v_0)
			;
		// Trace: design.sv:70462:5
		dma_write_fsm_n_state = 1'd0;
		// Trace: design.sv:70463:5
		dma_done = 1'b0;
		// Trace: design.sv:70465:5
		data_out_req = 1'sb0;
		// Trace: design.sv:70466:5
		data_out_we = 1'sb0;
		// Trace: design.sv:70467:5
		data_out_be = 1'sb0;
		// Trace: design.sv:70468:5
		data_out_addr = 1'sb0;
		// Trace: design.sv:70470:5
		(* full_case, parallel_case *)
		case (dma_write_fsm_state)
			1'd0:
				// Trace: design.sv:70474:9
				if (dma_start == 1'b1)
					// Trace: design.sv:70475:11
					dma_write_fsm_n_state = 1'd1;
				else
					// Trace: design.sv:70477:11
					dma_write_fsm_n_state = 1'd0;
			1'd1:
				// Trace: design.sv:70483:9
				if ((fifo_empty == 1'b1) && (dma_read_fsm_state == 1'd0)) begin
					// Trace: design.sv:70484:11
					dma_write_fsm_n_state = 1'd0;
					// Trace: design.sv:70485:11
					dma_done = 1'b1;
				end
				else begin
					// Trace: design.sv:70487:11
					dma_write_fsm_n_state = 1'd1;
					// Trace: design.sv:70489:11
					if ((fifo_empty == 1'b0) && (wait_for_tx_spi == 1'b0)) begin
						// Trace: design.sv:70490:13
						data_out_req = 1'b1;
						// Trace: design.sv:70491:13
						data_out_we = 1'b1;
						// Trace: design.sv:70492:13
						data_out_be = byte_enable_out;
						// Trace: design.sv:70493:13
						data_out_addr = write_ptr_reg;
					end
				end
		endcase
	end
	// Trace: design.sv:70500:3
	fifo_v3 #(.DEPTH(FIFO_DEPTH)) dma_fifo_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(fifo_flush),
		.testmode_i(1'b0),
		.full_o(fifo_full),
		.empty_o(fifo_empty),
		.usage_o(fifo_usage),
		.data_i(fifo_input),
		.push_i(data_in_rvalid),
		.data_o(fifo_output),
		.pop_i(data_out_gnt)
	);
	// Trace: design.sv:70519:3
	dma_reg_top_A4ADD dma_reg_top_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(reg_req_i),
		.reg_rsp_o(reg_rsp_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.devmode_i(1'b1)
	);
	initial _sv2v_0 = 0;
endmodule
// removed package "obi_spimemio_reg_pkg"
module obi_spimemio_reg_top_73C2E (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	reg2hw,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:70583:20
	// removed localparam type reg_req_t
	// Trace: design.sv:70584:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:70585:15
	parameter signed [31:0] AW = 3;
	// Trace: design.sv:70587:5
	input clk_i;
	// Trace: design.sv:70588:5
	input rst_ni;
	// Trace: design.sv:70589:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:70590:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:70592:5
	// removed localparam type obi_spimemio_reg_pkg_obi_spimemio_reg2hw_start_spimem_reg_t
	// removed localparam type obi_spimemio_reg_pkg_obi_spimemio_reg2hw_t
	output wire [0:0] reg2hw;
	// Trace: design.sv:70596:5
	input devmode_i;
	// Trace: design.sv:70599:3
	// removed import obi_spimemio_reg_pkg::*;
	// Trace: design.sv:70601:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:70602:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:70605:3
	wire reg_we;
	// Trace: design.sv:70606:3
	wire reg_re;
	// Trace: design.sv:70607:3
	wire [AW - 1:0] reg_addr;
	// Trace: design.sv:70608:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:70609:3
	wire [3:0] reg_be;
	// Trace: design.sv:70610:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:70611:3
	wire reg_error;
	// Trace: design.sv:70613:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:70615:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:70618:3
	wire [69:0] reg_intf_req;
	// Trace: design.sv:70619:3
	wire [33:0] reg_intf_rsp;
	// Trace: design.sv:70622:3
	assign reg_intf_req = reg_req_i;
	// Trace: design.sv:70623:3
	assign reg_rsp_o = reg_intf_rsp;
	// Trace: design.sv:70626:3
	assign reg_we = reg_intf_req[69] & reg_intf_req[68];
	// Trace: design.sv:70627:3
	assign reg_re = reg_intf_req[69] & ~reg_intf_req[68];
	// Trace: design.sv:70628:3
	assign reg_addr = reg_intf_req[63-:32];
	// Trace: design.sv:70629:3
	assign reg_wdata = reg_intf_req[31-:32];
	// Trace: design.sv:70630:3
	assign reg_be = reg_intf_req[67-:4];
	// Trace: design.sv:70631:3
	assign reg_intf_rsp[31-:32] = reg_rdata;
	// Trace: design.sv:70632:3
	assign reg_intf_rsp[33] = reg_error;
	// Trace: design.sv:70633:3
	assign reg_intf_rsp[32] = 1'b1;
	// Trace: design.sv:70635:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:70636:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:70642:3
	wire start_spimem_qs;
	// Trace: design.sv:70643:3
	wire start_spimem_wd;
	// Trace: design.sv:70644:3
	wire start_spimem_we;
	// Trace: design.sv:70649:3
	localparam signed [31:0] sv2v_uu_u_start_spimem_DW = 1;
	// removed localparam type sv2v_uu_u_start_spimem_d
	localparam [0:0] sv2v_uu_u_start_spimem_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_start_spimem(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(start_spimem_we),
		.wd(start_spimem_wd),
		.de(1'b0),
		.d(sv2v_uu_u_start_spimem_ext_d_0),
		.qe(),
		.q(reg2hw[-0]),
		.qs(start_spimem_qs)
	);
	// Trace: design.sv:70676:3
	localparam signed [31:0] sv2v_uu_u_cfg_spimem_DW = 32;
	// removed localparam type sv2v_uu_u_cfg_spimem_wd
	localparam [31:0] sv2v_uu_u_cfg_spimem_ext_wd_0 = 1'sb0;
	// removed localparam type sv2v_uu_u_cfg_spimem_d
	localparam [31:0] sv2v_uu_u_cfg_spimem_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("NONE"),
		.RESVAL(32'h00000000)
	) u_cfg_spimem(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_cfg_spimem_ext_wd_0),
		.de(1'b0),
		.d(sv2v_uu_u_cfg_spimem_ext_d_0),
		.qe(),
		.q(),
		.qs()
	);
	// Trace: design.sv:70701:3
	reg [1:0] addr_hit;
	// Trace: design.sv:70702:3
	localparam signed [31:0] obi_spimemio_reg_pkg_BlockAw = 3;
	localparam [2:0] obi_spimemio_reg_pkg_OBI_SPIMEMIO_CFG_SPIMEM_OFFSET = 3'h4;
	localparam [2:0] obi_spimemio_reg_pkg_OBI_SPIMEMIO_START_SPIMEM_OFFSET = 3'h0;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:70703:5
		addr_hit = 1'sb0;
		// Trace: design.sv:70704:5
		addr_hit[0] = reg_addr == obi_spimemio_reg_pkg_OBI_SPIMEMIO_START_SPIMEM_OFFSET;
		// Trace: design.sv:70705:5
		addr_hit[1] = reg_addr == obi_spimemio_reg_pkg_OBI_SPIMEMIO_CFG_SPIMEM_OFFSET;
	end
	// Trace: design.sv:70708:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:70711:3
	localparam [7:0] obi_spimemio_reg_pkg_OBI_SPIMEMIO_PERMIT = 8'b00011111;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:70712:5
		wr_err = reg_we & ((addr_hit[0] & |(obi_spimemio_reg_pkg_OBI_SPIMEMIO_PERMIT[4+:4] & ~reg_be)) | (addr_hit[1] & |(obi_spimemio_reg_pkg_OBI_SPIMEMIO_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:70717:3
	assign start_spimem_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:70718:3
	assign start_spimem_wd = reg_wdata[0];
	// Trace: design.sv:70721:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:70722:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:70723:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]:
				// Trace: design.sv:70725:9
				reg_rdata_next[0] = start_spimem_qs;
			addr_hit[1]:
				// Trace: design.sv:70729:9
				reg_rdata_next[31:0] = 1'sb0;
			default:
				// Trace: design.sv:70733:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:70742:3
	wire unused_wdata;
	// Trace: design.sv:70743:3
	wire unused_be;
	// Trace: design.sv:70744:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:70745:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
// removed package "picorv32_pkg"
module obi_to_picorv32 (
	clk_i,
	rst_ni,
	obi_req_i,
	obi_resp_o,
	picorv32_req_o,
	picorv32_resp_i
);
	reg _sv2v_0;
	// removed import obi_pkg::*;
	// removed import picorv32_pkg::*;
	// Trace: design.sv:70783:5
	input wire clk_i;
	// Trace: design.sv:70784:5
	input wire rst_ni;
	// Trace: design.sv:70786:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [69:0] obi_req_i;
	// Trace: design.sv:70787:5
	// removed localparam type obi_pkg_obi_resp_t
	output reg [33:0] obi_resp_o;
	// Trace: design.sv:70789:5
	// removed localparam type picorv32_pkg_picorv32_req_t
	output reg [68:0] picorv32_req_o;
	// Trace: design.sv:70790:5
	// removed localparam type picorv32_pkg_picorv32_resp_t
	input wire [32:0] picorv32_resp_i;
	// Trace: design.sv:70793:3
	// removed localparam type picorv_request_e
	// Trace: design.sv:70804:3
	reg [1:0] state;
	reg [1:0] state_next;
	// Trace: design.sv:70813:3
	reg [31:0] addr_buf;
	reg [31:0] addr_buf_next;
	reg [31:0] rdata_buf;
	reg [31:0] rdata_buf_next;
	// Trace: design.sv:70816:3
	always @(posedge clk_i or negedge rst_ni) begin : ram_valid_q
		// Trace: design.sv:70817:5
		if (!rst_ni) begin
			// Trace: design.sv:70818:7
			state <= 2'd0;
			// Trace: design.sv:70819:7
			addr_buf <= 1'sb0;
			// Trace: design.sv:70820:7
			rdata_buf <= 1'sb0;
		end
		else begin
			// Trace: design.sv:70822:7
			state <= state_next;
			// Trace: design.sv:70823:7
			addr_buf <= addr_buf_next;
			// Trace: design.sv:70824:7
			rdata_buf <= rdata_buf_next;
		end
	end
	// Trace: design.sv:70829:3
	always @(*) begin : fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:70831:5
		addr_buf_next = addr_buf;
		// Trace: design.sv:70832:5
		state_next = state;
		// Trace: design.sv:70833:5
		picorv32_req_o[68] = 1'b0;
		// Trace: design.sv:70834:5
		picorv32_req_o[63-:32] = 1'sb0;
		// Trace: design.sv:70835:5
		picorv32_req_o[31-:32] = 1'sb0;
		// Trace: design.sv:70836:5
		picorv32_req_o[67-:4] = 4'b0000;
		// Trace: design.sv:70837:5
		obi_resp_o[33] = 1'b0;
		// Trace: design.sv:70838:5
		obi_resp_o[32] = 1'b0;
		// Trace: design.sv:70839:5
		obi_resp_o[31-:32] = rdata_buf;
		// Trace: design.sv:70840:5
		rdata_buf_next = picorv32_resp_i[31-:32];
		// Trace: design.sv:70842:5
		case (state)
			2'd0:
				// Trace: design.sv:70844:9
				if (obi_req_i[69]) begin
					begin
						// Trace: design.sv:70845:11
						if (obi_req_i[68] == 1'b1) begin
							// Trace: design.sv:70846:13
							state_next = 2'd2;
							// Trace: design.sv:70847:13
							obi_resp_o[33] = 1'b1;
						end
						else begin
							// Trace: design.sv:70849:13
							state_next = 2'd1;
							// Trace: design.sv:70850:13
							addr_buf_next = obi_req_i[63-:32];
							// Trace: design.sv:70851:13
							obi_resp_o[33] = 1'b1;
						end
					end
				end
			2'd1: begin
				// Trace: design.sv:70856:9
				picorv32_req_o[63-:32] = addr_buf;
				// Trace: design.sv:70857:9
				picorv32_req_o[68] = 1'b1;
				// Trace: design.sv:70858:9
				if (picorv32_resp_i[32])
					// Trace: design.sv:70859:11
					state_next = 2'd3;
			end
			2'd2: begin
				// Trace: design.sv:70864:9
				state_next = 2'd0;
				// Trace: design.sv:70865:9
				obi_resp_o[32] = 1'b1;
			end
			2'd3: begin
				// Trace: design.sv:70869:9
				state_next = 2'd0;
				// Trace: design.sv:70870:9
				obi_resp_o[32] = 1'b1;
			end
			default:
				// Trace: design.sv:70874:9
				state_next = 2'd0;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module obi_spimemio (
	clk_i,
	rst_ni,
	flash_csb_o,
	flash_clk_o,
	flash_io0_oe_o,
	flash_io1_oe_o,
	flash_io2_oe_o,
	flash_io3_oe_o,
	flash_io0_do_o,
	flash_io1_do_o,
	flash_io2_do_o,
	flash_io3_do_o,
	flash_io0_di_i,
	flash_io1_di_i,
	flash_io2_di_i,
	flash_io3_di_i,
	reg_req_i,
	reg_rsp_o,
	spimemio_req_i,
	spimemio_resp_o
);
	reg _sv2v_0;
	// removed import obi_pkg::*;
	// removed import reg_pkg::*;
	// Trace: design.sv:70892:5
	input wire clk_i;
	// Trace: design.sv:70893:5
	input wire rst_ni;
	// Trace: design.sv:70894:5
	output wire flash_csb_o;
	// Trace: design.sv:70895:5
	output wire flash_clk_o;
	// Trace: design.sv:70897:5
	output wire flash_io0_oe_o;
	// Trace: design.sv:70898:5
	output wire flash_io1_oe_o;
	// Trace: design.sv:70899:5
	output wire flash_io2_oe_o;
	// Trace: design.sv:70900:5
	output wire flash_io3_oe_o;
	// Trace: design.sv:70902:5
	output wire flash_io0_do_o;
	// Trace: design.sv:70903:5
	output wire flash_io1_do_o;
	// Trace: design.sv:70904:5
	output wire flash_io2_do_o;
	// Trace: design.sv:70905:5
	output wire flash_io3_do_o;
	// Trace: design.sv:70907:5
	input wire flash_io0_di_i;
	// Trace: design.sv:70908:5
	input wire flash_io1_di_i;
	// Trace: design.sv:70909:5
	input wire flash_io2_di_i;
	// Trace: design.sv:70910:5
	input wire flash_io3_di_i;
	// Trace: design.sv:70912:5
	// removed localparam type reg_pkg_reg_req_t
	input wire [69:0] reg_req_i;
	// Trace: design.sv:70913:5
	// removed localparam type reg_pkg_reg_rsp_t
	output reg [33:0] reg_rsp_o;
	// Trace: design.sv:70915:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [69:0] spimemio_req_i;
	// Trace: design.sv:70916:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [33:0] spimemio_resp_o;
	// Trace: design.sv:70919:3
	// removed import picorv32_pkg::*;
	// Trace: design.sv:70920:3
	// removed import obi_spimemio_reg_pkg::*;
	// Trace: design.sv:70922:3
	// removed localparam type picorv32_pkg_picorv32_req_t
	wire [68:0] picorv32_req;
	// Trace: design.sv:70923:3
	// removed localparam type picorv32_pkg_picorv32_resp_t
	wire [32:0] picorv32_resp;
	// Trace: design.sv:70925:3
	wire [33:0] reg_rsp_reg;
	reg [33:0] reg_rsp_spimem;
	// Trace: design.sv:70927:3
	wire [31:0] cfgreg_do;
	// Trace: design.sv:70928:3
	wire cfgreg_we;
	wire cfgreg_rd;
	// Trace: design.sv:70930:3
	// removed localparam type obi_spimemio_reg_pkg_obi_spimemio_reg2hw_start_spimem_reg_t
	// removed localparam type obi_spimemio_reg_pkg_obi_spimemio_reg2hw_t
	wire [0:0] reg2hw;
	// Trace: design.sv:70932:3
	obi_to_picorv32 obi_to_picorv32_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.picorv32_req_o(picorv32_req),
		.picorv32_resp_i(picorv32_resp),
		.obi_req_i(spimemio_req_i),
		.obi_resp_o(spimemio_resp_o)
	);
	// Trace: design.sv:70941:3
	obi_spimemio_reg_top_73C2E obi_spimemio_reg_top_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(reg_req_i),
		.reg_rsp_o(reg_rsp_reg),
		.reg2hw(reg2hw),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:70953:3
	localparam signed [31:0] obi_spimemio_reg_pkg_BlockAw = 3;
	localparam [2:0] obi_spimemio_reg_pkg_OBI_SPIMEMIO_CFG_SPIMEM_OFFSET = 3'h4;
	assign cfgreg_we = (reg_req_i[69] & reg_req_i[68]) && (reg_req_i[34:32] == obi_spimemio_reg_pkg_OBI_SPIMEMIO_CFG_SPIMEM_OFFSET);
	// Trace: design.sv:70954:3
	assign cfgreg_rd = (reg_req_i[69] & ~reg_req_i[68]) && (reg_req_i[34:32] == obi_spimemio_reg_pkg_OBI_SPIMEMIO_CFG_SPIMEM_OFFSET);
	// Trace: design.sv:70956:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:70957:5
		reg_rsp_spimem[31-:32] = cfgreg_do;
		// Trace: design.sv:70958:5
		reg_rsp_spimem[33] = 1'b0;
		// Trace: design.sv:70959:5
		reg_rsp_spimem[32] = 1'b1;
		// Trace: design.sv:70961:5
		if (cfgreg_rd)
			// Trace: design.sv:70962:7
			reg_rsp_o = reg_rsp_spimem;
		else
			// Trace: design.sv:70964:7
			reg_rsp_o = reg_rsp_reg;
	end
	// Trace: design.sv:70968:3
	spimemio spimemio_i(
		.clk(clk_i),
		.resetn(rst_ni),
		.start_spi_i(reg2hw[-0]),
		.valid(picorv32_req[68]),
		.ready(picorv32_resp[32]),
		.addr({picorv32_req[55:34], 2'b00}),
		.rdata(picorv32_resp[31-:32]),
		.flash_csb(flash_csb_o),
		.flash_clk(flash_clk_o),
		.flash_io0_oe(flash_io0_oe_o),
		.flash_io1_oe(flash_io1_oe_o),
		.flash_io2_oe(flash_io2_oe_o),
		.flash_io3_oe(flash_io3_oe_o),
		.flash_io0_do(flash_io0_do_o),
		.flash_io1_do(flash_io1_do_o),
		.flash_io2_do(flash_io2_do_o),
		.flash_io3_do(flash_io3_do_o),
		.flash_io0_di(flash_io0_di_i),
		.flash_io1_di(flash_io1_di_i),
		.flash_io2_di(flash_io2_di_i),
		.flash_io3_di(flash_io3_di_i),
		.cfgreg_we({4 {cfgreg_we}}),
		.cfgreg_di(reg_req_i[31-:32]),
		.cfgreg_do(cfgreg_do)
	);
	initial _sv2v_0 = 0;
endmodule
module prim_buf (
	in_i,
	out_o
);
	// Trace: design.sv:71017:13
	parameter signed [31:0] Width = 1;
	// Trace: design.sv:71020:3
	input [Width - 1:0] in_i;
	// Trace: design.sv:71021:3
	output wire [Width - 1:0] out_o;
	// Trace: design.sv:71024:3
	generate
		if (1) begin : gen_generic
			// Trace: design.sv:71025:5
			prim_generic_buf #(.Width(Width)) u_impl_generic(
				.in_i(in_i),
				.out_o(out_o)
			);
		end
	endgenerate
endmodule
module prim_clock_mux2 (
	clk0_i,
	clk1_i,
	sel_i,
	clk_o
);
	// Trace: design.sv:71051:13
	parameter [0:0] NoFpgaBufG = 1'b0;
	// Trace: design.sv:71054:3
	input clk0_i;
	// Trace: design.sv:71055:3
	input clk1_i;
	// Trace: design.sv:71056:3
	input sel_i;
	// Trace: design.sv:71057:3
	output wire clk_o;
	// Trace: design.sv:71060:3
	generate
		if (1) begin : gen_generic
			// Trace: design.sv:71061:5
			prim_generic_clock_mux2 #(.NoFpgaBufG(NoFpgaBufG)) u_impl_generic(
				.clk0_i(clk0_i),
				.clk1_i(clk1_i),
				.sel_i(sel_i),
				.clk_o(clk_o)
			);
		end
	endgenerate
endmodule
module prim_flop (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	// Trace: design.sv:71087:13
	parameter signed [31:0] Width = 1;
	// Trace: design.sv:71088:13
	parameter [Width - 1:0] ResetValue = 0;
	// Trace: design.sv:71091:3
	input clk_i;
	// Trace: design.sv:71092:3
	input rst_ni;
	// Trace: design.sv:71093:3
	input [Width - 1:0] d_i;
	// Trace: design.sv:71094:3
	output wire [Width - 1:0] q_o;
	// Trace: design.sv:71097:3
	generate
		if (1) begin : gen_generic
			// Trace: design.sv:71098:5
			prim_generic_flop #(
				.Width(Width),
				.ResetValue(ResetValue)
			) u_impl_generic(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(d_i),
				.q_o(q_o)
			);
		end
	endgenerate
endmodule
module prim_flop_2sync (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	// Trace: design.sv:71125:13
	parameter signed [31:0] Width = 16;
	// Trace: design.sv:71126:13
	parameter [Width - 1:0] ResetValue = 1'sb0;
	// Trace: design.sv:71129:3
	input clk_i;
	// Trace: design.sv:71130:3
	input rst_ni;
	// Trace: design.sv:71131:3
	input [Width - 1:0] d_i;
	// Trace: design.sv:71132:3
	output wire [Width - 1:0] q_o;
	// Trace: design.sv:71135:3
	generate
		if (1) begin : gen_generic
			// Trace: design.sv:71136:5
			prim_generic_flop_2sync #(
				.Width(Width),
				.ResetValue(ResetValue)
			) u_impl_generic(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(d_i),
				.q_o(q_o)
			);
		end
	endgenerate
endmodule
module prim_flop_en (
	clk_i,
	rst_ni,
	en_i,
	d_i,
	q_o
);
	// Trace: design.sv:71163:13
	parameter signed [31:0] Width = 1;
	// Trace: design.sv:71164:13
	parameter [Width - 1:0] ResetValue = 0;
	// Trace: design.sv:71167:3
	input clk_i;
	// Trace: design.sv:71168:3
	input rst_ni;
	// Trace: design.sv:71169:3
	input en_i;
	// Trace: design.sv:71170:3
	input [Width - 1:0] d_i;
	// Trace: design.sv:71171:3
	output wire [Width - 1:0] q_o;
	// Trace: design.sv:71174:3
	generate
		if (1) begin : gen_generic
			// Trace: design.sv:71175:5
			prim_generic_flop_en #(
				.ResetValue(ResetValue),
				.Width(Width)
			) u_impl_generic(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.en_i(en_i),
				.d_i(d_i),
				.q_o(q_o)
			);
		end
	endgenerate
endmodule
module prim_xor2 (
	in0_i,
	in1_i,
	out_o
);
	// Trace: design.sv:71202:13
	parameter signed [31:0] Width = 1;
	// Trace: design.sv:71205:3
	input [Width - 1:0] in0_i;
	// Trace: design.sv:71206:3
	input [Width - 1:0] in1_i;
	// Trace: design.sv:71207:3
	output wire [Width - 1:0] out_o;
	// Trace: design.sv:71210:3
	generate
		if (1) begin : gen_generic
			// Trace: design.sv:71211:5
			prim_generic_xor2 #(.Width(Width)) u_impl_generic(
				.in0_i(in0_i),
				.in1_i(in1_i),
				.out_o(out_o)
			);
		end
	endgenerate
endmodule
// removed package "prim_alert_pkg"
module prim_alert_receiver (
	clk_i,
	rst_ni,
	ping_req_i,
	ping_ok_o,
	integ_fail_o,
	alert_o,
	alert_rx_o,
	alert_tx_i
);
	reg _sv2v_0;
	// removed import prim_alert_pkg::*;
	// Trace: design.sv:71283:13
	parameter [0:0] AsyncOn = 1'b0;
	// Trace: design.sv:71285:3
	input clk_i;
	// Trace: design.sv:71286:3
	input rst_ni;
	// Trace: design.sv:71289:3
	input ping_req_i;
	// Trace: design.sv:71290:3
	output reg ping_ok_o;
	// Trace: design.sv:71292:3
	output reg integ_fail_o;
	// Trace: design.sv:71295:3
	output reg alert_o;
	// Trace: design.sv:71297:3
	// removed localparam type prim_alert_pkg_alert_rx_t
	output wire [3:0] alert_rx_o;
	// Trace: design.sv:71299:3
	// removed localparam type prim_alert_pkg_alert_tx_t
	input wire [1:0] alert_tx_i;
	// Trace: design.sv:71306:3
	wire alert_level;
	wire alert_sigint;
	// Trace: design.sv:71308:3
	prim_diff_decode #(.AsyncOn(AsyncOn)) i_decode_alert(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(alert_tx_i[1]),
		.diff_ni(alert_tx_i[0]),
		.level_o(alert_level),
		.rise_o(),
		.fall_o(),
		.event_o(),
		.sigint_o(alert_sigint)
	);
	// Trace: design.sv:71325:3
	// removed localparam type state_e
	// Trace: design.sv:71326:3
	reg [1:0] state_d;
	reg [1:0] state_q;
	// Trace: design.sv:71327:3
	wire ping_rise;
	// Trace: design.sv:71328:3
	wire ping_tog;
	wire ping_tog_dp;
	reg ping_tog_qp;
	wire ping_tog_dn;
	reg ping_tog_qn;
	// Trace: design.sv:71329:3
	reg ack;
	wire ack_dp;
	reg ack_qp;
	wire ack_dn;
	reg ack_qn;
	// Trace: design.sv:71330:3
	wire ping_req_d;
	reg ping_req_q;
	// Trace: design.sv:71331:3
	wire ping_pending_d;
	reg ping_pending_q;
	// Trace: design.sv:71335:3
	assign ping_req_d = ping_req_i;
	// Trace: design.sv:71336:3
	assign ping_rise = ping_req_i && !ping_req_q;
	// Trace: design.sv:71337:3
	assign ping_tog = (ping_rise ? ~ping_tog_qp : ping_tog_qp);
	// Trace: design.sv:71340:3
	prim_buf u_prim_buf_ack_p(
		.in_i(ack),
		.out_o(ack_dp)
	);
	// Trace: design.sv:71344:3
	prim_buf u_prim_buf_ack_n(
		.in_i(~ack),
		.out_o(ack_dn)
	);
	// Trace: design.sv:71348:3
	prim_buf u_prim_buf_ping_p(
		.in_i(ping_tog),
		.out_o(ping_tog_dp)
	);
	// Trace: design.sv:71352:3
	prim_buf u_prim_buf_ping_n(
		.in_i(~ping_tog),
		.out_o(ping_tog_dn)
	);
	// Trace: design.sv:71362:3
	assign ping_pending_d = ping_rise | ((~ping_ok_o & ping_req_i) & ping_pending_q);
	// Trace: design.sv:71365:3
	assign alert_rx_o[1] = ack_qp;
	// Trace: design.sv:71366:3
	assign alert_rx_o[0] = ack_qn;
	// Trace: design.sv:71368:3
	assign alert_rx_o[3] = ping_tog_qp;
	// Trace: design.sv:71369:3
	assign alert_rx_o[2] = ping_tog_qn;
	// Trace: design.sv:71375:3
	always @(*) begin : p_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:71377:5
		state_d = state_q;
		// Trace: design.sv:71378:5
		ack = 1'b0;
		// Trace: design.sv:71379:5
		ping_ok_o = 1'b0;
		// Trace: design.sv:71380:5
		integ_fail_o = 1'b0;
		// Trace: design.sv:71381:5
		alert_o = 1'b0;
		// Trace: design.sv:71383:5
		(* full_case, parallel_case *)
		case (state_q)
			2'd0:
				// Trace: design.sv:71386:9
				if (alert_level) begin
					// Trace: design.sv:71387:11
					state_d = 2'd1;
					// Trace: design.sv:71388:11
					ack = 1'b1;
					// Trace: design.sv:71390:11
					if (ping_pending_q)
						// Trace: design.sv:71391:13
						ping_ok_o = 1'b1;
					else
						// Trace: design.sv:71393:13
						alert_o = 1'b1;
				end
			2'd1:
				// Trace: design.sv:71399:9
				if (!alert_level)
					// Trace: design.sv:71400:11
					state_d = 2'd2;
				else
					// Trace: design.sv:71402:11
					ack = 1'b1;
			2'd2:
				// Trace: design.sv:71406:15
				state_d = 2'd3;
			2'd3:
				// Trace: design.sv:71407:15
				state_d = 2'd0;
			default:
				;
		endcase
		if (alert_sigint) begin
			// Trace: design.sv:71413:7
			state_d = 2'd0;
			// Trace: design.sv:71414:7
			ack = 1'b0;
			// Trace: design.sv:71415:7
			ping_ok_o = 1'b0;
			// Trace: design.sv:71416:7
			integ_fail_o = 1'b1;
			// Trace: design.sv:71417:7
			alert_o = 1'b0;
		end
	end
	// Trace: design.sv:71421:3
	always @(posedge clk_i or negedge rst_ni) begin : p_reg
		// Trace: design.sv:71422:5
		if (!rst_ni) begin
			// Trace: design.sv:71423:7
			state_q <= 2'd0;
			// Trace: design.sv:71424:7
			ack_qp <= 1'b0;
			// Trace: design.sv:71425:7
			ack_qn <= 1'b1;
			// Trace: design.sv:71426:7
			ping_tog_qp <= 1'b0;
			// Trace: design.sv:71427:7
			ping_tog_qn <= 1'b1;
			// Trace: design.sv:71428:7
			ping_req_q <= 1'b0;
			// Trace: design.sv:71429:7
			ping_pending_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:71431:7
			state_q <= state_d;
			// Trace: design.sv:71432:7
			ack_qp <= ack_dp;
			// Trace: design.sv:71433:7
			ack_qn <= ack_dn;
			// Trace: design.sv:71434:7
			ping_tog_qp <= ping_tog_dp;
			// Trace: design.sv:71435:7
			ping_tog_qn <= ping_tog_dn;
			// Trace: design.sv:71436:7
			ping_req_q <= ping_req_d;
			// Trace: design.sv:71437:7
			ping_pending_q <= ping_pending_d;
		end
	end
	// Trace: design.sv:71462:3
	initial _sv2v_0 = 0;
endmodule
module prim_alert_sender (
	clk_i,
	rst_ni,
	alert_test_i,
	alert_req_i,
	alert_ack_o,
	alert_state_o,
	alert_rx_i,
	alert_tx_o
);
	reg _sv2v_0;
	// removed import prim_alert_pkg::*;
	// Trace: design.sv:71533:13
	parameter [0:0] AsyncOn = 1'b1;
	// Trace: design.sv:71536:13
	parameter [0:0] IsFatal = 1'b0;
	// Trace: design.sv:71538:3
	input clk_i;
	// Trace: design.sv:71539:3
	input rst_ni;
	// Trace: design.sv:71541:3
	input alert_test_i;
	// Trace: design.sv:71543:3
	input alert_req_i;
	// Trace: design.sv:71544:3
	output wire alert_ack_o;
	// Trace: design.sv:71546:3
	output wire alert_state_o;
	// Trace: design.sv:71548:3
	// removed localparam type prim_alert_pkg_alert_rx_t
	input wire [3:0] alert_rx_i;
	// Trace: design.sv:71550:3
	// removed localparam type prim_alert_pkg_alert_tx_t
	output wire [1:0] alert_tx_o;
	// Trace: design.sv:71557:3
	wire ping_sigint;
	wire ping_event;
	// Trace: design.sv:71559:3
	prim_diff_decode #(.AsyncOn(AsyncOn)) i_decode_ping(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(alert_rx_i[3]),
		.diff_ni(alert_rx_i[2]),
		.level_o(),
		.rise_o(),
		.fall_o(),
		.event_o(ping_event),
		.sigint_o(ping_sigint)
	);
	// Trace: design.sv:71573:3
	wire ack_sigint;
	wire ack_level;
	// Trace: design.sv:71575:3
	prim_diff_decode #(.AsyncOn(AsyncOn)) i_decode_ack(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(alert_rx_i[1]),
		.diff_ni(alert_rx_i[0]),
		.level_o(ack_level),
		.rise_o(),
		.fall_o(),
		.event_o(),
		.sigint_o(ack_sigint)
	);
	// Trace: design.sv:71593:3
	// removed localparam type state_e
	// Trace: design.sv:71603:3
	reg [2:0] state_d;
	reg [2:0] state_q;
	// Trace: design.sv:71604:3
	reg alert_p;
	reg alert_n;
	reg alert_pq;
	reg alert_nq;
	wire alert_pd;
	wire alert_nd;
	// Trace: design.sv:71605:3
	wire sigint_detected;
	// Trace: design.sv:71607:3
	assign sigint_detected = ack_sigint | ping_sigint;
	// Trace: design.sv:71611:3
	assign alert_tx_o[1] = alert_pq;
	// Trace: design.sv:71612:3
	assign alert_tx_o[0] = alert_nq;
	// Trace: design.sv:71615:3
	wire alert_set_d;
	reg alert_set_q;
	reg alert_clr;
	// Trace: design.sv:71616:3
	wire alert_test_set_d;
	reg alert_test_set_q;
	// Trace: design.sv:71617:3
	wire ping_set_d;
	reg ping_set_q;
	reg ping_clr;
	// Trace: design.sv:71618:3
	wire alert_req_trigger;
	wire alert_test_trigger;
	wire ping_trigger;
	// Trace: design.sv:71621:3
	assign alert_req_trigger = alert_req_i | alert_set_q;
	// Trace: design.sv:71622:3
	generate
		if (IsFatal) begin : gen_fatal
			// Trace: design.sv:71623:5
			assign alert_set_d = alert_req_trigger;
		end
		else begin : gen_recov
			// Trace: design.sv:71625:5
			assign alert_set_d = (alert_clr ? 1'b0 : alert_req_trigger);
		end
	endgenerate
	// Trace: design.sv:71629:3
	assign alert_test_trigger = alert_test_i | alert_test_set_q;
	// Trace: design.sv:71630:3
	assign alert_test_set_d = (alert_clr ? 1'b0 : alert_test_trigger);
	// Trace: design.sv:71632:3
	wire alert_trigger;
	// Trace: design.sv:71633:3
	assign alert_trigger = alert_req_trigger | alert_test_trigger;
	// Trace: design.sv:71635:3
	assign ping_trigger = ping_set_q | ping_event;
	// Trace: design.sv:71636:3
	assign ping_set_d = (ping_clr ? 1'b0 : ping_trigger);
	// Trace: design.sv:71640:3
	assign alert_ack_o = alert_clr & alert_set_q;
	// Trace: design.sv:71641:3
	assign alert_state_o = alert_set_q;
	// Trace: design.sv:71649:3
	always @(*) begin : p_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:71651:5
		state_d = state_q;
		// Trace: design.sv:71652:5
		alert_p = 1'b0;
		// Trace: design.sv:71653:5
		alert_n = 1'b1;
		// Trace: design.sv:71654:5
		ping_clr = 1'b0;
		// Trace: design.sv:71655:5
		alert_clr = 1'b0;
		// Trace: design.sv:71657:5
		(* full_case, parallel_case *)
		case (state_q)
			3'd0:
				// Trace: design.sv:71660:9
				if (alert_trigger || ping_trigger) begin
					// Trace: design.sv:71661:11
					state_d = (alert_trigger ? 3'd1 : 3'd3);
					// Trace: design.sv:71662:11
					alert_p = 1'b1;
					// Trace: design.sv:71663:11
					alert_n = 1'b0;
				end
			3'd1:
				// Trace: design.sv:71668:9
				if (ack_level)
					// Trace: design.sv:71669:11
					state_d = 3'd2;
				else begin
					// Trace: design.sv:71671:11
					alert_p = 1'b1;
					// Trace: design.sv:71672:11
					alert_n = 1'b0;
				end
			3'd2:
				// Trace: design.sv:71677:9
				if (!ack_level) begin
					// Trace: design.sv:71678:11
					state_d = 3'd6;
					// Trace: design.sv:71679:11
					alert_clr = 1'b1;
				end
			3'd3:
				// Trace: design.sv:71684:9
				if (ack_level)
					// Trace: design.sv:71685:11
					state_d = 3'd4;
				else begin
					// Trace: design.sv:71687:11
					alert_p = 1'b1;
					// Trace: design.sv:71688:11
					alert_n = 1'b0;
				end
			3'd4:
				// Trace: design.sv:71693:9
				if (!ack_level) begin
					// Trace: design.sv:71694:11
					ping_clr = 1'b1;
					// Trace: design.sv:71695:11
					state_d = 3'd6;
				end
			3'd6:
				// Trace: design.sv:71700:9
				state_d = 3'd7;
			3'd7:
				// Trace: design.sv:71705:9
				state_d = 3'd0;
			3'd5: begin
				// Trace: design.sv:71714:9
				state_d = 3'd0;
				// Trace: design.sv:71715:9
				if (sigint_detected) begin
					// Trace: design.sv:71716:11
					state_d = 3'd5;
					// Trace: design.sv:71717:11
					alert_p = ~alert_pq;
					// Trace: design.sv:71718:11
					alert_n = ~alert_pq;
				end
			end
			default:
				// Trace: design.sv:71722:17
				state_d = 3'd0;
		endcase
		if (sigint_detected && (state_q != 3'd5)) begin
			// Trace: design.sv:71726:7
			state_d = 3'd5;
			// Trace: design.sv:71727:7
			alert_p = 1'b0;
			// Trace: design.sv:71728:7
			alert_n = 1'b0;
			// Trace: design.sv:71729:7
			ping_clr = 1'b0;
			// Trace: design.sv:71730:7
			alert_clr = 1'b0;
		end
	end
	// Trace: design.sv:71735:3
	prim_buf u_prim_buf_p(
		.in_i(alert_p),
		.out_o(alert_pd)
	);
	// Trace: design.sv:71739:3
	prim_buf u_prim_buf_n(
		.in_i(alert_n),
		.out_o(alert_nd)
	);
	// Trace: design.sv:71744:3
	always @(posedge clk_i or negedge rst_ni) begin : p_reg
		// Trace: design.sv:71745:5
		if (!rst_ni) begin
			// Trace: design.sv:71746:7
			state_q <= 3'd0;
			// Trace: design.sv:71747:7
			alert_pq <= 1'b0;
			// Trace: design.sv:71748:7
			alert_nq <= 1'b1;
			// Trace: design.sv:71749:7
			alert_set_q <= 1'b0;
			// Trace: design.sv:71750:7
			alert_test_set_q <= 1'b0;
			// Trace: design.sv:71751:7
			ping_set_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:71753:7
			state_q <= state_d;
			// Trace: design.sv:71754:7
			alert_pq <= alert_pd;
			// Trace: design.sv:71755:7
			alert_nq <= alert_nd;
			// Trace: design.sv:71756:7
			alert_set_q <= alert_set_d;
			// Trace: design.sv:71757:7
			alert_test_set_q <= alert_test_set_d;
			// Trace: design.sv:71758:7
			ping_set_q <= ping_set_d;
		end
	end
	// Trace: design.sv:71770:3
	// Trace: design.sv:71807:3
	initial _sv2v_0 = 0;
endmodule
module prim_fifo_async (
	clk_wr_i,
	rst_wr_ni,
	wvalid_i,
	wready_o,
	wdata_i,
	wdepth_o,
	clk_rd_i,
	rst_rd_ni,
	rvalid_o,
	rready_i,
	rdata_o,
	rdepth_o
);
	// Trace: design.sv:71837:14
	parameter [31:0] Width = 16;
	// Trace: design.sv:71838:14
	parameter [31:0] Depth = 4;
	// Trace: design.sv:71839:14
	parameter [0:0] OutputZeroIfEmpty = 1'b0;
	// Trace: design.sv:71840:14
	localparam [31:0] DepthW = $clog2(Depth + 1);
	// Trace: design.sv:71843:3
	input wire clk_wr_i;
	// Trace: design.sv:71844:3
	input wire rst_wr_ni;
	// Trace: design.sv:71845:3
	input wire wvalid_i;
	// Trace: design.sv:71846:3
	output wire wready_o;
	// Trace: design.sv:71847:3
	input wire [Width - 1:0] wdata_i;
	// Trace: design.sv:71848:3
	output wire [DepthW - 1:0] wdepth_o;
	// Trace: design.sv:71851:3
	input wire clk_rd_i;
	// Trace: design.sv:71852:3
	input wire rst_rd_ni;
	// Trace: design.sv:71853:3
	output wire rvalid_o;
	// Trace: design.sv:71854:3
	input wire rready_i;
	// Trace: design.sv:71855:3
	output wire [Width - 1:0] rdata_o;
	// Trace: design.sv:71856:3
	output wire [DepthW - 1:0] rdepth_o;
	// Trace: design.sv:71862:3
	localparam [31:0] PTRV_W = (Depth == 1 ? 1 : $clog2(Depth));
	// Trace: design.sv:71863:3
	localparam [31:0] PTR_WIDTH = (Depth == 1 ? 1 : PTRV_W + 1);
	// Trace: design.sv:71865:3
	reg [PTR_WIDTH - 1:0] fifo_wptr_q;
	wire [PTR_WIDTH - 1:0] fifo_wptr_d;
	// Trace: design.sv:71866:3
	reg [PTR_WIDTH - 1:0] fifo_rptr_q;
	wire [PTR_WIDTH - 1:0] fifo_rptr_d;
	// Trace: design.sv:71867:3
	wire [PTR_WIDTH - 1:0] fifo_wptr_sync_combi;
	wire [PTR_WIDTH - 1:0] fifo_rptr_sync_combi;
	// Trace: design.sv:71868:3
	wire [PTR_WIDTH - 1:0] fifo_wptr_gray_sync;
	wire [PTR_WIDTH - 1:0] fifo_rptr_gray_sync;
	reg [PTR_WIDTH - 1:0] fifo_rptr_sync_q;
	// Trace: design.sv:71869:3
	reg [PTR_WIDTH - 1:0] fifo_wptr_gray_q;
	wire [PTR_WIDTH - 1:0] fifo_wptr_gray_d;
	// Trace: design.sv:71870:3
	reg [PTR_WIDTH - 1:0] fifo_rptr_gray_q;
	wire [PTR_WIDTH - 1:0] fifo_rptr_gray_d;
	// Trace: design.sv:71871:3
	wire fifo_incr_wptr;
	wire fifo_incr_rptr;
	// Trace: design.sv:71872:3
	wire full_wclk;
	wire full_rclk;
	wire empty_rclk;
	// Trace: design.sv:71873:3
	reg [Width - 1:0] storage [0:Depth - 1];
	// Trace: design.sv:71879:3
	assign fifo_incr_wptr = wvalid_i & wready_o;
	// Trace: design.sv:71882:3
	function automatic signed [PTR_WIDTH - 1:0] sv2v_cast_62A53_signed;
		input reg signed [PTR_WIDTH - 1:0] inp;
		sv2v_cast_62A53_signed = inp;
	endfunction
	assign fifo_wptr_d = fifo_wptr_q + sv2v_cast_62A53_signed(1);
	// Trace: design.sv:71884:3
	always @(posedge clk_wr_i or negedge rst_wr_ni)
		// Trace: design.sv:71885:5
		if (!rst_wr_ni)
			// Trace: design.sv:71886:7
			fifo_wptr_q <= 1'sb0;
		else if (fifo_incr_wptr)
			// Trace: design.sv:71888:7
			fifo_wptr_q <= fifo_wptr_d;
	// Trace: design.sv:71893:3
	always @(posedge clk_wr_i or negedge rst_wr_ni)
		// Trace: design.sv:71894:5
		if (!rst_wr_ni)
			// Trace: design.sv:71895:7
			fifo_wptr_gray_q <= 1'sb0;
		else if (fifo_incr_wptr)
			// Trace: design.sv:71897:7
			fifo_wptr_gray_q <= fifo_wptr_gray_d;
	// Trace: design.sv:71902:3
	prim_flop_2sync #(.Width(PTR_WIDTH)) sync_wptr(
		.clk_i(clk_rd_i),
		.rst_ni(rst_rd_ni),
		.d_i(fifo_wptr_gray_q),
		.q_o(fifo_wptr_gray_sync)
	);
	// Trace: design.sv:71912:3
	assign fifo_incr_rptr = rvalid_o & rready_i;
	// Trace: design.sv:71915:3
	assign fifo_rptr_d = fifo_rptr_q + sv2v_cast_62A53_signed(1);
	// Trace: design.sv:71917:3
	always @(posedge clk_rd_i or negedge rst_rd_ni)
		// Trace: design.sv:71918:5
		if (!rst_rd_ni)
			// Trace: design.sv:71919:7
			fifo_rptr_q <= 1'sb0;
		else if (fifo_incr_rptr)
			// Trace: design.sv:71921:7
			fifo_rptr_q <= fifo_rptr_d;
	// Trace: design.sv:71926:3
	always @(posedge clk_rd_i or negedge rst_rd_ni)
		// Trace: design.sv:71927:5
		if (!rst_rd_ni)
			// Trace: design.sv:71928:7
			fifo_rptr_gray_q <= 1'sb0;
		else if (fifo_incr_rptr)
			// Trace: design.sv:71930:7
			fifo_rptr_gray_q <= fifo_rptr_gray_d;
	// Trace: design.sv:71935:3
	prim_flop_2sync #(.Width(PTR_WIDTH)) sync_rptr(
		.clk_i(clk_wr_i),
		.rst_ni(rst_wr_ni),
		.d_i(fifo_rptr_gray_q),
		.q_o(fifo_rptr_gray_sync)
	);
	// Trace: design.sv:71942:3
	always @(posedge clk_wr_i or negedge rst_wr_ni)
		// Trace: design.sv:71943:5
		if (!rst_wr_ni)
			// Trace: design.sv:71944:7
			fifo_rptr_sync_q <= 1'sb0;
		else
			// Trace: design.sv:71946:7
			fifo_rptr_sync_q <= fifo_rptr_sync_combi;
	// Trace: design.sv:71954:3
	assign full_wclk = fifo_wptr_q == (fifo_rptr_sync_q ^ {1'b1, {PTR_WIDTH - 1 {1'b0}}});
	// Trace: design.sv:71955:3
	assign full_rclk = fifo_wptr_sync_combi == (fifo_rptr_q ^ {1'b1, {PTR_WIDTH - 1 {1'b0}}});
	// Trace: design.sv:71956:3
	assign empty_rclk = fifo_wptr_sync_combi == fifo_rptr_q;
	// Trace: design.sv:71958:3
	function automatic [DepthW - 1:0] sv2v_cast_2DA09;
		input reg [DepthW - 1:0] inp;
		sv2v_cast_2DA09 = inp;
	endfunction
	generate
		if (Depth > 1) begin : g_depth_calc
			// Trace: design.sv:71961:5
			wire wptr_msb;
			// Trace: design.sv:71962:5
			wire rptr_sync_msb;
			// Trace: design.sv:71963:5
			wire [PTRV_W - 1:0] wptr_value;
			// Trace: design.sv:71964:5
			wire [PTRV_W - 1:0] rptr_sync_value;
			// Trace: design.sv:71966:5
			assign wptr_msb = fifo_wptr_q[PTR_WIDTH - 1];
			// Trace: design.sv:71967:5
			assign rptr_sync_msb = fifo_rptr_sync_q[PTR_WIDTH - 1];
			// Trace: design.sv:71968:5
			assign wptr_value = fifo_wptr_q[0+:PTRV_W];
			// Trace: design.sv:71969:5
			assign rptr_sync_value = fifo_rptr_sync_q[0+:PTRV_W];
			// Trace: design.sv:71970:5
			assign wdepth_o = (full_wclk ? sv2v_cast_2DA09(Depth) : (wptr_msb == rptr_sync_msb ? sv2v_cast_2DA09(wptr_value) - sv2v_cast_2DA09(rptr_sync_value) : (sv2v_cast_2DA09(Depth) - sv2v_cast_2DA09(rptr_sync_value)) + sv2v_cast_2DA09(wptr_value)));
			// Trace: design.sv:71975:5
			wire rptr_msb;
			// Trace: design.sv:71976:5
			wire wptr_sync_msb;
			// Trace: design.sv:71977:5
			wire [PTRV_W - 1:0] rptr_value;
			// Trace: design.sv:71978:5
			wire [PTRV_W - 1:0] wptr_sync_value;
			// Trace: design.sv:71980:5
			assign wptr_sync_msb = fifo_wptr_sync_combi[PTR_WIDTH - 1];
			// Trace: design.sv:71981:5
			assign rptr_msb = fifo_rptr_q[PTR_WIDTH - 1];
			// Trace: design.sv:71982:5
			assign wptr_sync_value = fifo_wptr_sync_combi[0+:PTRV_W];
			// Trace: design.sv:71983:5
			assign rptr_value = fifo_rptr_q[0+:PTRV_W];
			// Trace: design.sv:71984:5
			assign rdepth_o = (full_rclk ? sv2v_cast_2DA09(Depth) : (wptr_sync_msb == rptr_msb ? sv2v_cast_2DA09(wptr_sync_value) - sv2v_cast_2DA09(rptr_value) : (sv2v_cast_2DA09(Depth) - sv2v_cast_2DA09(rptr_value)) + sv2v_cast_2DA09(wptr_sync_value)));
		end
		else begin : g_no_depth_calc
			// Trace: design.sv:71990:5
			assign rdepth_o = full_rclk;
			// Trace: design.sv:71991:5
			assign wdepth_o = full_wclk;
		end
	endgenerate
	// Trace: design.sv:71995:3
	assign wready_o = !full_wclk;
	// Trace: design.sv:71996:3
	assign rvalid_o = !empty_rclk;
	// Trace: design.sv:72002:3
	wire [Width - 1:0] rdata_int;
	// Trace: design.sv:72003:3
	generate
		if (Depth > 1) begin : g_storage_mux
			// Trace: design.sv:72005:5
			always @(posedge clk_wr_i)
				// Trace: design.sv:72006:7
				if (fifo_incr_wptr)
					// Trace: design.sv:72007:9
					storage[fifo_wptr_q[PTRV_W - 1:0]] <= wdata_i;
			// Trace: design.sv:72011:5
			assign rdata_int = storage[fifo_rptr_q[PTRV_W - 1:0]];
		end
		else begin : g_storage_simple
			// Trace: design.sv:72015:5
			always @(posedge clk_wr_i)
				// Trace: design.sv:72016:7
				if (fifo_incr_wptr)
					// Trace: design.sv:72017:9
					storage[0] <= wdata_i;
			// Trace: design.sv:72021:5
			assign rdata_int = storage[0];
		end
	endgenerate
	// Trace: design.sv:72025:3
	generate
		if (OutputZeroIfEmpty == 1'b1) begin : gen_output_zero
			// Trace: design.sv:72026:5
			assign rdata_o = (empty_rclk ? {Width {1'sb0}} : rdata_int);
		end
		else begin : gen_no_output_zero
			// Trace: design.sv:72028:5
			assign rdata_o = rdata_int;
		end
	endgenerate
	// Trace: design.sv:72036:3
	function automatic [PTR_WIDTH - 1:0] sv2v_cast_62A53;
		input reg [PTR_WIDTH - 1:0] inp;
		sv2v_cast_62A53 = inp;
	endfunction
	function automatic [((PTR_WIDTH - 2) >= 0 ? PTR_WIDTH - 1 : 3 - PTR_WIDTH) - 1:0] sv2v_cast_0A027;
		input reg [((PTR_WIDTH - 2) >= 0 ? PTR_WIDTH - 1 : 3 - PTR_WIDTH) - 1:0] inp;
		sv2v_cast_0A027 = inp;
	endfunction
	generate
		if (Depth > 2) begin : g_full_gray_conversion
			// Trace: design.sv:72038:5
			function automatic [PTR_WIDTH - 1:0] dec2gray;
				// Trace: design.sv:72038:49
				input reg [PTR_WIDTH - 1:0] decval;
				// Trace: design.sv:72039:7
				reg [PTR_WIDTH - 1:0] decval_sub;
				// Trace: design.sv:72040:7
				reg [PTR_WIDTH - 2:0] decval_in;
				// Trace: design.sv:72041:7
				reg unused_decval_msb;
				begin
					// Trace: design.sv:72043:7
					decval_sub = (sv2v_cast_62A53(Depth) - {1'b0, decval[PTR_WIDTH - 2:0]}) - 1'b1;
					// Trace: design.sv:72045:7
					{unused_decval_msb, decval_in} = (decval[PTR_WIDTH - 1] ? decval_sub : decval);
					// Trace: design.sv:72048:7
					dec2gray = {decval[PTR_WIDTH - 1], {1'b0, decval_in[PTR_WIDTH - 2:1]} ^ decval_in[PTR_WIDTH - 2:0]};
				end
			endfunction
			// Trace: design.sv:72053:5
			function automatic [PTR_WIDTH - 1:0] gray2dec;
				// Trace: design.sv:72053:49
				input reg [PTR_WIDTH - 1:0] grayval;
				// Trace: design.sv:72054:7
				reg [PTR_WIDTH - 2:0] dec_tmp;
				reg [PTR_WIDTH - 2:0] dec_tmp_sub;
				// Trace: design.sv:72055:7
				reg unused_decsub_msb;
				begin
					// Trace: design.sv:72057:7
					dec_tmp[PTR_WIDTH - 2] = grayval[PTR_WIDTH - 2];
					// Trace: design.sv:72058:7
					begin : sv2v_autoblock_1
						// Trace: design.sv:72058:12
						reg signed [31:0] i;
						// Trace: design.sv:72058:12
						for (i = PTR_WIDTH - 3; i >= 0; i = i - 1)
							begin
								// Trace: design.sv:72059:9
								dec_tmp[i] = dec_tmp[i + 1] ^ grayval[i];
							end
					end
					// Trace: design.sv:72061:7
					{unused_decsub_msb, dec_tmp_sub} = (sv2v_cast_0A027(Depth) - {1'b0, dec_tmp}) - 1'b1;
					if (grayval[PTR_WIDTH - 1])
						// Trace: design.sv:72063:9
						gray2dec = {1'b1, dec_tmp_sub};
					else
						// Trace: design.sv:72065:9
						gray2dec = {1'b0, dec_tmp};
				end
			endfunction
			// Trace: design.sv:72070:5
			assign fifo_rptr_sync_combi = gray2dec(fifo_rptr_gray_sync);
			// Trace: design.sv:72072:5
			assign fifo_wptr_sync_combi = gray2dec(fifo_wptr_gray_sync);
			// Trace: design.sv:72074:5
			assign fifo_rptr_gray_d = dec2gray(fifo_rptr_d);
			// Trace: design.sv:72075:5
			assign fifo_wptr_gray_d = dec2gray(fifo_wptr_d);
		end
		else if (Depth == 2) begin : g_simple_gray_conversion
			// Trace: design.sv:72079:5
			assign fifo_rptr_sync_combi = {fifo_rptr_gray_sync[PTR_WIDTH - 1], ^fifo_rptr_gray_sync};
			// Trace: design.sv:72080:5
			assign fifo_wptr_sync_combi = {fifo_wptr_gray_sync[PTR_WIDTH - 1], ^fifo_rptr_gray_sync};
			// Trace: design.sv:72082:5
			assign fifo_rptr_gray_d = {fifo_rptr_d[PTR_WIDTH - 1], ^fifo_rptr_d};
			// Trace: design.sv:72083:5
			assign fifo_wptr_gray_d = {fifo_wptr_d[PTR_WIDTH - 1], ^fifo_rptr_d};
		end
		else begin : g_no_gray_conversion
			// Trace: design.sv:72087:5
			assign fifo_rptr_sync_combi = fifo_rptr_gray_sync;
			// Trace: design.sv:72088:5
			assign fifo_wptr_sync_combi = fifo_wptr_gray_sync;
			// Trace: design.sv:72090:5
			assign fifo_rptr_gray_d = fifo_rptr_d;
			// Trace: design.sv:72091:5
			assign fifo_wptr_gray_d = fifo_rptr_d;
		end
	endgenerate
endmodule
module prim_fifo_sync (
	clk_i,
	rst_ni,
	clr_i,
	wvalid_i,
	wready_o,
	wdata_i,
	rvalid_o,
	rready_i,
	rdata_o,
	full_o,
	depth_o
);
	// Trace: design.sv:72111:13
	parameter [31:0] Width = 16;
	// Trace: design.sv:72112:13
	parameter [0:0] Pass = 1'b1;
	// Trace: design.sv:72113:13
	parameter [31:0] Depth = 4;
	// Trace: design.sv:72114:13
	parameter [0:0] OutputZeroIfEmpty = 1'b1;
	// Trace: design.sv:72116:14
	function automatic integer prim_util_pkg_vbits;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:74:36
		input integer value;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:85:5
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] DepthW = prim_util_pkg_vbits(Depth + 1);
	// Trace: design.sv:72118:3
	input clk_i;
	// Trace: design.sv:72119:3
	input rst_ni;
	// Trace: design.sv:72121:3
	input clr_i;
	// Trace: design.sv:72123:3
	input wvalid_i;
	// Trace: design.sv:72124:3
	output wire wready_o;
	// Trace: design.sv:72125:3
	input [Width - 1:0] wdata_i;
	// Trace: design.sv:72127:3
	output wire rvalid_o;
	// Trace: design.sv:72128:3
	input rready_i;
	// Trace: design.sv:72129:3
	output wire [Width - 1:0] rdata_o;
	// Trace: design.sv:72131:3
	output wire full_o;
	// Trace: design.sv:72132:3
	output wire [DepthW - 1:0] depth_o;
	// Trace: design.sv:72137:3
	function automatic [DepthW - 1:0] sv2v_cast_2DA09;
		input reg [DepthW - 1:0] inp;
		sv2v_cast_2DA09 = inp;
	endfunction
	generate
		if (Depth == 0) begin : gen_passthru_fifo
			// Trace: design.sv:72140:5
			assign depth_o = 1'b0;
			// Trace: design.sv:72143:5
			assign rvalid_o = wvalid_i;
			// Trace: design.sv:72144:5
			assign rdata_o = wdata_i;
			// Trace: design.sv:72147:5
			assign wready_o = rready_i;
			// Trace: design.sv:72148:5
			assign full_o = rready_i;
			// Trace: design.sv:72151:5
			wire unused_clr;
			// Trace: design.sv:72152:5
			assign unused_clr = clr_i;
		end
		else begin : gen_normal_fifo
			// Trace: design.sv:72157:5
			localparam [31:0] PTRV_W = prim_util_pkg_vbits(Depth);
			// Trace: design.sv:72158:5
			localparam [31:0] PTR_WIDTH = PTRV_W + 1;
			// Trace: design.sv:72160:5
			reg [PTR_WIDTH - 1:0] fifo_wptr;
			reg [PTR_WIDTH - 1:0] fifo_rptr;
			// Trace: design.sv:72161:5
			wire fifo_incr_wptr;
			wire fifo_incr_rptr;
			wire fifo_empty;
			// Trace: design.sv:72164:5
			reg under_rst;
			// Trace: design.sv:72165:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:72166:7
				if (!rst_ni)
					// Trace: design.sv:72167:9
					under_rst <= 1'b1;
				else if (under_rst)
					// Trace: design.sv:72169:9
					under_rst <= ~under_rst;
			// Trace: design.sv:72174:5
			wire full;
			wire empty;
			// Trace: design.sv:72175:5
			wire wptr_msb;
			// Trace: design.sv:72176:5
			wire rptr_msb;
			// Trace: design.sv:72177:5
			wire [PTRV_W - 1:0] wptr_value;
			// Trace: design.sv:72178:5
			wire [PTRV_W - 1:0] rptr_value;
			// Trace: design.sv:72180:5
			assign wptr_msb = fifo_wptr[PTR_WIDTH - 1];
			// Trace: design.sv:72181:5
			assign rptr_msb = fifo_rptr[PTR_WIDTH - 1];
			// Trace: design.sv:72182:5
			assign wptr_value = fifo_wptr[0+:PTRV_W];
			// Trace: design.sv:72183:5
			assign rptr_value = fifo_rptr[0+:PTRV_W];
			// Trace: design.sv:72184:5
			assign depth_o = (full ? sv2v_cast_2DA09(Depth) : (wptr_msb == rptr_msb ? sv2v_cast_2DA09(wptr_value) - sv2v_cast_2DA09(rptr_value) : (sv2v_cast_2DA09(Depth) - sv2v_cast_2DA09(rptr_value)) + sv2v_cast_2DA09(wptr_value)));
			// Trace: design.sv:72188:5
			assign fifo_incr_wptr = (wvalid_i & wready_o) & ~under_rst;
			// Trace: design.sv:72189:5
			assign fifo_incr_rptr = (rvalid_o & rready_i) & ~under_rst;
			// Trace: design.sv:72194:5
			assign wready_o = ~full & ~under_rst;
			// Trace: design.sv:72195:5
			assign full_o = full;
			// Trace: design.sv:72196:5
			assign rvalid_o = ~empty & ~under_rst;
			// Trace: design.sv:72198:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:72199:7
				if (!rst_ni)
					// Trace: design.sv:72200:9
					fifo_wptr <= {PTR_WIDTH {1'b0}};
				else if (clr_i)
					// Trace: design.sv:72202:9
					fifo_wptr <= {PTR_WIDTH {1'b0}};
				else if (fifo_incr_wptr)
					// Trace: design.sv:72204:9
					begin : sv2v_autoblock_1
						reg [((PTR_WIDTH - 2) >= 0 ? PTR_WIDTH - 1 : 3 - PTR_WIDTH) - 1:0] sv2v_tmp_cast;
						sv2v_tmp_cast = Depth - 1;
						if (fifo_wptr[PTR_WIDTH - 2:0] == sv2v_tmp_cast)
							// Trace: design.sv:72205:11
							fifo_wptr <= {~fifo_wptr[PTR_WIDTH - 1], {PTR_WIDTH - 1 {1'b0}}};
						else
							// Trace: design.sv:72207:11
							fifo_wptr <= fifo_wptr + {{PTR_WIDTH - 1 {1'b0}}, 1'b1};
					end
			// Trace: design.sv:72212:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:72213:7
				if (!rst_ni)
					// Trace: design.sv:72214:9
					fifo_rptr <= {PTR_WIDTH {1'b0}};
				else if (clr_i)
					// Trace: design.sv:72216:9
					fifo_rptr <= {PTR_WIDTH {1'b0}};
				else if (fifo_incr_rptr)
					// Trace: design.sv:72218:9
					begin : sv2v_autoblock_2
						reg [((PTR_WIDTH - 2) >= 0 ? PTR_WIDTH - 1 : 3 - PTR_WIDTH) - 1:0] sv2v_tmp_cast;
						sv2v_tmp_cast = Depth - 1;
						if (fifo_rptr[PTR_WIDTH - 2:0] == sv2v_tmp_cast)
							// Trace: design.sv:72219:11
							fifo_rptr <= {~fifo_rptr[PTR_WIDTH - 1], {PTR_WIDTH - 1 {1'b0}}};
						else
							// Trace: design.sv:72221:11
							fifo_rptr <= fifo_rptr + {{PTR_WIDTH - 1 {1'b0}}, 1'b1};
					end
			// Trace: design.sv:72226:5
			assign full = fifo_wptr == (fifo_rptr ^ {1'b1, {PTR_WIDTH - 1 {1'b0}}});
			// Trace: design.sv:72227:5
			assign fifo_empty = fifo_wptr == fifo_rptr;
			// Trace: design.sv:72232:5
			reg [(Depth * Width) - 1:0] storage;
			// Trace: design.sv:72233:5
			wire [Width - 1:0] storage_rdata;
			if (Depth == 1) begin : gen_depth_eq1
				// Trace: design.sv:72235:7
				assign storage_rdata = storage[0+:Width];
				// Trace: design.sv:72237:7
				always @(posedge clk_i)
					if (fifo_incr_wptr)
						// Trace: design.sv:72239:11
						storage[0+:Width] <= wdata_i;
			end
			else begin : gen_depth_gt1
				// Trace: design.sv:72243:7
				assign storage_rdata = storage[fifo_rptr[PTR_WIDTH - 2:0] * Width+:Width];
				// Trace: design.sv:72245:7
				always @(posedge clk_i)
					if (fifo_incr_wptr)
						// Trace: design.sv:72247:11
						storage[fifo_wptr[PTR_WIDTH - 2:0] * Width+:Width] <= wdata_i;
			end
			// Trace: design.sv:72251:5
			wire [Width - 1:0] rdata_int;
			if (Pass == 1'b1) begin : gen_pass
				// Trace: design.sv:72253:7
				assign rdata_int = (fifo_empty && wvalid_i ? wdata_i : storage_rdata);
				// Trace: design.sv:72254:7
				assign empty = fifo_empty & ~wvalid_i;
			end
			else begin : gen_nopass
				// Trace: design.sv:72256:7
				assign rdata_int = storage_rdata;
				// Trace: design.sv:72257:7
				assign empty = fifo_empty;
			end
			if (OutputZeroIfEmpty == 1'b1) begin : gen_output_zero
				// Trace: design.sv:72261:7
				assign rdata_o = (empty ? 'b0 : rdata_int);
			end
			else begin : gen_no_output_zero
				// Trace: design.sv:72263:7
				assign rdata_o = rdata_int;
			end
		end
	endgenerate
endmodule
module prim_clock_gating_sync (
	clk_i,
	rst_ni,
	test_en_i,
	async_en_i,
	en_o,
	clk_o
);
	// Trace: design.sv:72287:3
	input clk_i;
	// Trace: design.sv:72288:3
	input rst_ni;
	// Trace: design.sv:72289:3
	input test_en_i;
	// Trace: design.sv:72290:3
	input async_en_i;
	// Trace: design.sv:72291:3
	output wire en_o;
	// Trace: design.sv:72292:3
	output wire clk_o;
	// Trace: design.sv:72296:3
	prim_flop_2sync #(.Width(1)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(async_en_i),
		.q_o(en_o)
	);
	// Trace: design.sv:72305:3
	prim_clock_gating i_cg(
		.clk_i(clk_i),
		.en_i(en_o),
		.test_en_i(test_en_i),
		.clk_o(clk_o)
	);
endmodule
// removed package "prim_esc_pkg"
module prim_esc_receiver (
	clk_i,
	rst_ni,
	esc_en_o,
	esc_rx_o,
	esc_tx_i
);
	reg _sv2v_0;
	// removed import prim_esc_pkg::*;
	// Trace: design.sv:72360:3
	input clk_i;
	// Trace: design.sv:72361:3
	input rst_ni;
	// Trace: design.sv:72363:3
	output reg esc_en_o;
	// Trace: design.sv:72365:3
	// removed localparam type prim_esc_pkg_esc_rx_t
	output wire [1:0] esc_rx_o;
	// Trace: design.sv:72367:3
	// removed localparam type prim_esc_pkg_esc_tx_t
	input wire [1:0] esc_tx_i;
	// Trace: design.sv:72374:3
	wire esc_level;
	wire sigint_detected;
	// Trace: design.sv:72376:3
	prim_diff_decode #(.AsyncOn(1'b0)) i_decode_esc(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(esc_tx_i[1]),
		.diff_ni(esc_tx_i[0]),
		.level_o(esc_level),
		.rise_o(),
		.fall_o(),
		.event_o(),
		.sigint_o(sigint_detected)
	);
	// Trace: design.sv:72394:3
	// removed localparam type state_e
	// Trace: design.sv:72395:3
	reg [2:0] state_d;
	reg [2:0] state_q;
	// Trace: design.sv:72396:3
	reg resp_p;
	wire resp_pd;
	reg resp_pq;
	// Trace: design.sv:72397:3
	reg resp_n;
	wire resp_nd;
	reg resp_nq;
	// Trace: design.sv:72400:3
	prim_buf u_prim_buf_p(
		.in_i(resp_p),
		.out_o(resp_pd)
	);
	// Trace: design.sv:72404:3
	prim_buf u_prim_buf_n(
		.in_i(resp_n),
		.out_o(resp_nd)
	);
	// Trace: design.sv:72409:3
	assign esc_rx_o[1] = resp_pq;
	// Trace: design.sv:72410:3
	assign esc_rx_o[0] = resp_nq;
	// Trace: design.sv:72412:3
	always @(*) begin : p_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:72414:5
		state_d = state_q;
		// Trace: design.sv:72415:5
		resp_p = 1'b0;
		// Trace: design.sv:72416:5
		resp_n = 1'b1;
		// Trace: design.sv:72417:5
		esc_en_o = 1'b0;
		// Trace: design.sv:72419:5
		(* full_case, parallel_case *)
		case (state_q)
			3'd0:
				// Trace: design.sv:72422:9
				if (esc_level) begin
					// Trace: design.sv:72423:11
					state_d = 3'd1;
					// Trace: design.sv:72424:11
					resp_p = 1'b1;
					// Trace: design.sv:72425:11
					resp_n = 1'b0;
				end
			3'd1: begin
				// Trace: design.sv:72431:9
				state_d = 3'd2;
				// Trace: design.sv:72432:9
				if (esc_level) begin
					// Trace: design.sv:72433:11
					state_d = 3'd3;
					// Trace: design.sv:72434:11
					esc_en_o = 1'b1;
				end
			end
			3'd2: begin
				// Trace: design.sv:72440:9
				state_d = 3'd0;
				// Trace: design.sv:72441:9
				resp_p = 1'b1;
				// Trace: design.sv:72442:9
				resp_n = 1'b0;
				// Trace: design.sv:72443:9
				if (esc_level) begin
					// Trace: design.sv:72444:11
					state_d = 3'd3;
					// Trace: design.sv:72445:11
					esc_en_o = 1'b1;
				end
			end
			3'd3: begin
				// Trace: design.sv:72451:9
				state_d = 3'd0;
				// Trace: design.sv:72452:9
				if (esc_level) begin
					// Trace: design.sv:72453:11
					state_d = 3'd3;
					// Trace: design.sv:72454:11
					resp_p = ~resp_pq;
					// Trace: design.sv:72455:11
					resp_n = resp_pq;
					// Trace: design.sv:72456:11
					esc_en_o = 1'b1;
				end
			end
			3'd4: begin
				// Trace: design.sv:72465:9
				state_d = 3'd0;
				// Trace: design.sv:72466:9
				if (sigint_detected) begin
					// Trace: design.sv:72467:11
					state_d = 3'd4;
					// Trace: design.sv:72468:11
					resp_p = ~resp_pq;
					// Trace: design.sv:72469:11
					resp_n = ~resp_pq;
				end
			end
			default:
				// Trace: design.sv:72472:17
				state_d = 3'd0;
		endcase
		if (sigint_detected && (state_q != 3'd4)) begin
			// Trace: design.sv:72477:7
			state_d = 3'd4;
			// Trace: design.sv:72478:7
			resp_p = 1'b0;
			// Trace: design.sv:72479:7
			resp_n = 1'b0;
		end
	end
	// Trace: design.sv:72488:3
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:72489:5
		if (!rst_ni) begin
			// Trace: design.sv:72490:7
			state_q <= 3'd0;
			// Trace: design.sv:72491:7
			resp_pq <= 1'b0;
			// Trace: design.sv:72492:7
			resp_nq <= 1'b1;
		end
		else begin
			// Trace: design.sv:72494:7
			state_q <= state_d;
			// Trace: design.sv:72495:7
			resp_pq <= resp_pd;
			// Trace: design.sv:72496:7
			resp_nq <= resp_nd;
		end
	end
	initial _sv2v_0 = 0;
endmodule
module prim_esc_sender (
	clk_i,
	rst_ni,
	ping_req_i,
	ping_ok_o,
	integ_fail_o,
	esc_req_i,
	esc_rx_i,
	esc_tx_o
);
	reg _sv2v_0;
	// removed import prim_esc_pkg::*;
	// Trace: design.sv:72553:3
	input clk_i;
	// Trace: design.sv:72554:3
	input rst_ni;
	// Trace: design.sv:72556:3
	input ping_req_i;
	// Trace: design.sv:72557:3
	output reg ping_ok_o;
	// Trace: design.sv:72559:3
	output reg integ_fail_o;
	// Trace: design.sv:72561:3
	input esc_req_i;
	// Trace: design.sv:72563:3
	// removed localparam type prim_esc_pkg_esc_rx_t
	input wire [1:0] esc_rx_i;
	// Trace: design.sv:72565:3
	// removed localparam type prim_esc_pkg_esc_tx_t
	output wire [1:0] esc_tx_o;
	// Trace: design.sv:72572:3
	wire resp;
	wire sigint_detected;
	// Trace: design.sv:72574:3
	prim_diff_decode #(.AsyncOn(1'b0)) i_decode_resp(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(esc_rx_i[1]),
		.diff_ni(esc_rx_i[0]),
		.level_o(resp),
		.rise_o(),
		.fall_o(),
		.event_o(),
		.sigint_o(sigint_detected)
	);
	// Trace: design.sv:72592:3
	wire ping_req_d;
	reg ping_req_q;
	// Trace: design.sv:72593:3
	wire esc_req_d;
	reg esc_req_q;
	reg esc_req_q1;
	// Trace: design.sv:72595:3
	assign ping_req_d = ping_req_i;
	// Trace: design.sv:72596:3
	assign esc_req_d = esc_req_i;
	// Trace: design.sv:72600:3
	wire esc_p;
	// Trace: design.sv:72601:3
	assign esc_p = (esc_req_i | esc_req_q) | (ping_req_d & ~ping_req_q);
	// Trace: design.sv:72604:3
	prim_buf u_prim_buf_p(
		.in_i(esc_p),
		.out_o(esc_tx_o[1])
	);
	// Trace: design.sv:72608:3
	prim_buf u_prim_buf_n(
		.in_i(~esc_p),
		.out_o(esc_tx_o[0])
	);
	// Trace: design.sv:72617:3
	// removed localparam type fsm_e
	// Trace: design.sv:72620:3
	reg [2:0] state_d;
	reg [2:0] state_q;
	// Trace: design.sv:72622:3
	always @(*) begin : p_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:72624:5
		state_d = state_q;
		// Trace: design.sv:72625:5
		ping_ok_o = 1'b0;
		// Trace: design.sv:72626:5
		integ_fail_o = sigint_detected;
		// Trace: design.sv:72628:5
		(* full_case, parallel_case *)
		case (state_q)
			3'd0: begin
				// Trace: design.sv:72631:9
				if (esc_req_i)
					// Trace: design.sv:72632:11
					state_d = 3'd2;
				else if (ping_req_i)
					// Trace: design.sv:72634:11
					state_d = 3'd3;
				if (resp)
					// Trace: design.sv:72639:11
					integ_fail_o = 1'b1;
			end
			3'd1: begin
				// Trace: design.sv:72644:9
				state_d = 3'd2;
				// Trace: design.sv:72645:9
				if (!esc_tx_o[1] || resp) begin
					// Trace: design.sv:72646:11
					state_d = 3'd0;
					// Trace: design.sv:72647:11
					integ_fail_o = sigint_detected | resp;
				end
			end
			3'd2: begin
				// Trace: design.sv:72652:9
				state_d = 3'd1;
				// Trace: design.sv:72653:9
				if (!esc_tx_o[1] || !resp) begin
					// Trace: design.sv:72654:11
					state_d = 3'd0;
					// Trace: design.sv:72655:11
					integ_fail_o = sigint_detected | ~resp;
				end
			end
			3'd3: begin
				// Trace: design.sv:72661:9
				state_d = 3'd4;
				// Trace: design.sv:72664:9
				if (esc_req_i)
					// Trace: design.sv:72665:11
					state_d = 3'd1;
				else if (!resp) begin
					// Trace: design.sv:72668:11
					state_d = 3'd0;
					// Trace: design.sv:72669:11
					integ_fail_o = 1'b1;
				end
			end
			3'd4: begin
				// Trace: design.sv:72673:9
				state_d = 3'd5;
				// Trace: design.sv:72676:9
				if (esc_req_i)
					// Trace: design.sv:72677:11
					state_d = 3'd2;
				else if (resp) begin
					// Trace: design.sv:72680:11
					state_d = 3'd0;
					// Trace: design.sv:72681:11
					integ_fail_o = 1'b1;
				end
			end
			3'd5: begin
				// Trace: design.sv:72685:9
				state_d = 3'd6;
				// Trace: design.sv:72688:9
				if (esc_req_i)
					// Trace: design.sv:72689:11
					state_d = 3'd1;
				else if (!resp) begin
					// Trace: design.sv:72692:11
					state_d = 3'd0;
					// Trace: design.sv:72693:11
					integ_fail_o = 1'b1;
				end
			end
			3'd6: begin
				// Trace: design.sv:72697:9
				state_d = 3'd0;
				// Trace: design.sv:72700:9
				if (esc_req_i)
					// Trace: design.sv:72701:11
					state_d = 3'd2;
				else if (resp)
					// Trace: design.sv:72704:11
					integ_fail_o = 1'b1;
				else
					// Trace: design.sv:72706:11
					ping_ok_o = ping_req_i;
			end
			default:
				// Trace: design.sv:72709:17
				state_d = 3'd0;
		endcase
		if (sigint_detected) begin
			// Trace: design.sv:72716:7
			ping_ok_o = 1'b0;
			// Trace: design.sv:72717:7
			state_d = 3'd0;
		end
		if (((esc_req_i || esc_req_q) || esc_req_q1) && ping_req_i)
			// Trace: design.sv:72723:7
			ping_ok_o = 1'b1;
	end
	// Trace: design.sv:72731:3
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:72732:5
		if (!rst_ni) begin
			// Trace: design.sv:72733:7
			state_q <= 3'd0;
			// Trace: design.sv:72734:7
			esc_req_q <= 1'b0;
			// Trace: design.sv:72735:7
			esc_req_q1 <= 1'b0;
			// Trace: design.sv:72736:7
			ping_req_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:72738:7
			state_q <= state_d;
			// Trace: design.sv:72739:7
			esc_req_q <= esc_req_d;
			// Trace: design.sv:72740:7
			esc_req_q1 <= esc_req_q;
			// Trace: design.sv:72741:7
			ping_req_q <= ping_req_d;
		end
	end
	initial _sv2v_0 = 0;
endmodule
module prim_sram_arbiter (
	clk_i,
	rst_ni,
	req_i,
	req_addr_i,
	req_write_i,
	req_wdata_i,
	gnt_o,
	rsp_rvalid_o,
	rsp_rdata_o,
	rsp_error_o,
	sram_req_o,
	sram_addr_o,
	sram_write_o,
	sram_wdata_o,
	sram_rvalid_i,
	sram_rdata_i,
	sram_rerror_i
);
	// Trace: design.sv:72803:13
	parameter signed [31:0] N = 4;
	// Trace: design.sv:72804:13
	parameter signed [31:0] SramDw = 32;
	// Trace: design.sv:72805:13
	parameter signed [31:0] SramAw = 12;
	// Trace: design.sv:72806:13
	parameter ArbiterImpl = "PPC";
	// Trace: design.sv:72808:3
	input clk_i;
	// Trace: design.sv:72809:3
	input rst_ni;
	// Trace: design.sv:72811:3
	input [N - 1:0] req_i;
	// Trace: design.sv:72812:3
	input [(N * SramAw) - 1:0] req_addr_i;
	// Trace: design.sv:72813:3
	input [0:N - 1] req_write_i;
	// Trace: design.sv:72814:3
	input [(N * SramDw) - 1:0] req_wdata_i;
	// Trace: design.sv:72815:3
	output wire [N - 1:0] gnt_o;
	// Trace: design.sv:72817:3
	output wire [N - 1:0] rsp_rvalid_o;
	// Trace: design.sv:72818:3
	output wire [(N * SramDw) - 1:0] rsp_rdata_o;
	// Trace: design.sv:72819:3
	output wire [(N * 2) - 1:0] rsp_error_o;
	// Trace: design.sv:72822:3
	output wire sram_req_o;
	// Trace: design.sv:72823:3
	output wire [SramAw - 1:0] sram_addr_o;
	// Trace: design.sv:72824:3
	output wire sram_write_o;
	// Trace: design.sv:72825:3
	output wire [SramDw - 1:0] sram_wdata_o;
	// Trace: design.sv:72826:3
	input sram_rvalid_i;
	// Trace: design.sv:72827:3
	input [SramDw - 1:0] sram_rdata_i;
	// Trace: design.sv:72828:3
	input [1:0] sram_rerror_i;
	// Trace: design.sv:72832:3
	// removed localparam type req_t
	// Trace: design.sv:72838:3
	localparam signed [31:0] ARB_DW = (1 + SramAw) + SramDw;
	// Trace: design.sv:72840:3
	wire [(N * ((1 + SramAw) + SramDw)) - 1:0] req_packed;
	// Trace: design.sv:72842:3
	genvar _gv_i_83;
	generate
		for (_gv_i_83 = 0; _gv_i_83 < N; _gv_i_83 = _gv_i_83 + 1) begin : gen_reqs
			localparam i = _gv_i_83;
			// Trace: design.sv:72843:5
			assign req_packed[((N - 1) - i) * ((1 + SramAw) + SramDw)+:(1 + SramAw) + SramDw] = {req_write_i[i], req_addr_i[((N - 1) - i) * SramAw+:SramAw], req_wdata_i[((N - 1) - i) * SramDw+:SramDw]};
		end
	endgenerate
	// Trace: design.sv:72846:3
	wire [((1 + SramAw) + SramDw) - 1:0] sram_packed;
	// Trace: design.sv:72847:3
	assign sram_write_o = sram_packed[1 + (SramAw + (SramDw - 1))];
	// Trace: design.sv:72848:3
	assign sram_addr_o = sram_packed[SramAw + (SramDw - 1)-:((SramAw + (SramDw - 1)) >= (SramDw + 0) ? ((SramAw + (SramDw - 1)) - (SramDw + 0)) + 1 : ((SramDw + 0) - (SramAw + (SramDw - 1))) + 1)];
	// Trace: design.sv:72849:3
	assign sram_wdata_o = sram_packed[SramDw - 1-:SramDw];
	// Trace: design.sv:72851:3
	generate
		if (ArbiterImpl == "PPC") begin : gen_arb_ppc
			// Trace: design.sv:72852:5
			prim_arbiter_ppc #(
				.N(N),
				.DW(ARB_DW)
			) u_reqarb(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(req_i),
				.data_i(req_packed),
				.gnt_o(gnt_o),
				.idx_o(),
				.valid_o(sram_req_o),
				.data_o(sram_packed),
				.ready_i(1'b1)
			);
		end
		else if (ArbiterImpl == "BINTREE") begin : gen_tree_arb
			// Trace: design.sv:72867:5
			prim_arbiter_tree #(
				.N(N),
				.DW(ARB_DW)
			) u_reqarb(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(req_i),
				.data_i(req_packed),
				.gnt_o(gnt_o),
				.idx_o(),
				.valid_o(sram_req_o),
				.data_o(sram_packed),
				.ready_i(1'b1)
			);
		end
	endgenerate
	// Trace: design.sv:72886:3
	wire [N - 1:0] steer;
	// Trace: design.sv:72887:3
	wire sram_ack;
	// Trace: design.sv:72889:3
	assign sram_ack = sram_rvalid_i & |steer;
	// Trace: design.sv:72892:3
	prim_fifo_sync #(
		.Width(N),
		.Pass(1'b0),
		.Depth(4)
	) u_req_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(sram_req_o & ~sram_write_o),
		.wready_o(),
		.wdata_i(gnt_o),
		.rvalid_o(),
		.rready_i(sram_ack),
		.rdata_o(steer),
		.full_o(),
		.depth_o()
	);
	// Trace: design.sv:72910:3
	assign rsp_rvalid_o = steer & {N {sram_rvalid_i}};
	// Trace: design.sv:72912:3
	genvar _gv_i_84;
	generate
		for (_gv_i_84 = 0; _gv_i_84 < N; _gv_i_84 = _gv_i_84 + 1) begin : gen_rsp
			localparam i = _gv_i_84;
			// Trace: design.sv:72913:5
			assign rsp_rdata_o[((N - 1) - i) * SramDw+:SramDw] = sram_rdata_i;
			// Trace: design.sv:72914:5
			assign rsp_error_o[((N - 1) - i) * 2+:2] = sram_rerror_i;
		end
	endgenerate
endmodule
module prim_slicer (
	sel_i,
	data_i,
	data_o
);
	// Trace: design.sv:72928:13
	parameter signed [31:0] InW = 64;
	// Trace: design.sv:72929:13
	parameter signed [31:0] OutW = 8;
	// Trace: design.sv:72931:13
	parameter signed [31:0] IndexW = 4;
	// Trace: design.sv:72933:3
	input [IndexW - 1:0] sel_i;
	// Trace: design.sv:72934:3
	input [InW - 1:0] data_i;
	// Trace: design.sv:72935:3
	output wire [OutW - 1:0] data_o;
	// Trace: design.sv:72938:3
	localparam signed [31:0] UnrollW = OutW * (2 ** IndexW);
	// Trace: design.sv:72940:3
	wire [UnrollW - 1:0] unrolled_data;
	// Trace: design.sv:72942:3
	function automatic [UnrollW - 1:0] sv2v_cast_13D93;
		input reg [UnrollW - 1:0] inp;
		sv2v_cast_13D93 = inp;
	endfunction
	assign unrolled_data = sv2v_cast_13D93(data_i);
	// Trace: design.sv:72944:3
	assign data_o = unrolled_data[sel_i * OutW+:OutW];
endmodule
module prim_sync_reqack (
	clk_src_i,
	rst_src_ni,
	clk_dst_i,
	rst_dst_ni,
	src_req_i,
	src_ack_o,
	dst_req_o,
	dst_ack_i
);
	reg _sv2v_0;
	// Trace: design.sv:72977:13
	parameter [0:0] EnReqStabA = 1;
	// Trace: design.sv:72979:3
	input clk_src_i;
	// Trace: design.sv:72980:3
	input rst_src_ni;
	// Trace: design.sv:72981:3
	input clk_dst_i;
	// Trace: design.sv:72982:3
	input rst_dst_ni;
	// Trace: design.sv:72984:3
	input wire src_req_i;
	// Trace: design.sv:72985:3
	output reg src_ack_o;
	// Trace: design.sv:72986:3
	output reg dst_req_o;
	// Trace: design.sv:72987:3
	input wire dst_ack_i;
	// Trace: design.sv:72991:3
	// removed localparam type sync_reqack_fsm_e
	// Trace: design.sv:72996:3
	reg src_fsm_ns;
	reg src_fsm_cs;
	// Trace: design.sv:72997:3
	reg dst_fsm_ns;
	reg dst_fsm_cs;
	// Trace: design.sv:72998:3
	reg src_req_d;
	reg src_req_q;
	wire src_ack;
	// Trace: design.sv:72999:3
	reg dst_ack_d;
	reg dst_ack_q;
	wire dst_req;
	// Trace: design.sv:73000:3
	wire src_handshake;
	wire dst_handshake;
	// Trace: design.sv:73002:3
	assign src_handshake = src_req_i & src_ack_o;
	// Trace: design.sv:73003:3
	assign dst_handshake = dst_req_o & dst_ack_i;
	// Trace: design.sv:73006:3
	prim_flop_2sync #(.Width(1)) req_sync(
		.clk_i(clk_dst_i),
		.rst_ni(rst_dst_ni),
		.d_i(src_req_q),
		.q_o(dst_req)
	);
	// Trace: design.sv:73016:3
	prim_flop_2sync #(.Width(1)) ack_sync(
		.clk_i(clk_src_i),
		.rst_ni(rst_src_ni),
		.d_i(dst_ack_q),
		.q_o(src_ack)
	);
	// Trace: design.sv:73026:3
	always @(*) begin : src_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:73027:5
		src_fsm_ns = src_fsm_cs;
		// Trace: design.sv:73030:5
		src_req_d = src_req_q;
		// Trace: design.sv:73031:5
		src_ack_o = 1'b0;
		// Trace: design.sv:73033:5
		(* full_case, parallel_case *)
		case (src_fsm_cs)
			1'd0: begin
				// Trace: design.sv:73037:9
				src_req_d = src_req_i;
				// Trace: design.sv:73038:9
				src_ack_o = src_ack;
				// Trace: design.sv:73041:9
				if (src_handshake)
					// Trace: design.sv:73042:11
					src_fsm_ns = 1'd1;
			end
			1'd1: begin
				// Trace: design.sv:73049:9
				src_req_d = ~src_req_i;
				// Trace: design.sv:73050:9
				src_ack_o = ~src_ack;
				// Trace: design.sv:73053:9
				if (src_handshake)
					// Trace: design.sv:73054:11
					src_fsm_ns = 1'd0;
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:73063:3
	always @(*) begin : dst_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:73064:5
		dst_fsm_ns = dst_fsm_cs;
		// Trace: design.sv:73067:5
		dst_req_o = 1'b0;
		// Trace: design.sv:73068:5
		dst_ack_d = dst_ack_q;
		// Trace: design.sv:73070:5
		(* full_case, parallel_case *)
		case (dst_fsm_cs)
			1'd0: begin
				// Trace: design.sv:73074:9
				dst_req_o = dst_req;
				// Trace: design.sv:73075:9
				dst_ack_d = dst_ack_i;
				// Trace: design.sv:73078:9
				if (dst_handshake)
					// Trace: design.sv:73079:11
					dst_fsm_ns = 1'd1;
			end
			1'd1: begin
				// Trace: design.sv:73086:9
				dst_req_o = ~dst_req;
				// Trace: design.sv:73087:9
				dst_ack_d = ~dst_ack_i;
				// Trace: design.sv:73090:9
				if (dst_handshake)
					// Trace: design.sv:73091:11
					dst_fsm_ns = 1'd0;
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:73100:3
	always @(posedge clk_src_i or negedge rst_src_ni)
		// Trace: design.sv:73101:5
		if (!rst_src_ni) begin
			// Trace: design.sv:73102:7
			src_fsm_cs <= 1'd0;
			// Trace: design.sv:73103:7
			src_req_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:73105:7
			src_fsm_cs <= src_fsm_ns;
			// Trace: design.sv:73106:7
			src_req_q <= src_req_d;
		end
	// Trace: design.sv:73109:3
	always @(posedge clk_dst_i or negedge rst_dst_ni)
		// Trace: design.sv:73110:5
		if (!rst_dst_ni) begin
			// Trace: design.sv:73111:7
			dst_fsm_cs <= 1'd0;
			// Trace: design.sv:73112:7
			dst_ack_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:73114:7
			dst_fsm_cs <= dst_fsm_ns;
			// Trace: design.sv:73115:7
			dst_ack_q <= dst_ack_d;
		end
	// Trace: design.sv:73119:3
	initial _sv2v_0 = 0;
endmodule
module prim_sync_reqack_data (
	clk_src_i,
	rst_src_ni,
	clk_dst_i,
	rst_dst_ni,
	src_req_i,
	src_ack_o,
	dst_req_o,
	dst_ack_i,
	data_i,
	data_o
);
	// Trace: design.sv:73147:13
	parameter [31:0] Width = 1;
	// Trace: design.sv:73148:13
	parameter [0:0] DataSrc2Dst = 1'b1;
	// Trace: design.sv:73150:13
	parameter [0:0] DataReg = 1'b0;
	// Trace: design.sv:73152:13
	parameter [0:0] EnReqStabA = 1;
	// Trace: design.sv:73154:3
	input clk_src_i;
	// Trace: design.sv:73155:3
	input rst_src_ni;
	// Trace: design.sv:73156:3
	input clk_dst_i;
	// Trace: design.sv:73157:3
	input rst_dst_ni;
	// Trace: design.sv:73159:3
	input wire src_req_i;
	// Trace: design.sv:73160:3
	output wire src_ack_o;
	// Trace: design.sv:73161:3
	output wire dst_req_o;
	// Trace: design.sv:73162:3
	input wire dst_ack_i;
	// Trace: design.sv:73164:3
	input wire [Width - 1:0] data_i;
	// Trace: design.sv:73165:3
	output wire [Width - 1:0] data_o;
	// Trace: design.sv:73171:3
	prim_sync_reqack #(.EnReqStabA(EnReqStabA)) u_prim_sync_reqack(
		.clk_src_i(clk_src_i),
		.rst_src_ni(rst_src_ni),
		.clk_dst_i(clk_dst_i),
		.rst_dst_ni(rst_dst_ni),
		.src_req_i(src_req_i),
		.src_ack_o(src_ack_o),
		.dst_req_o(dst_req_o),
		.dst_ack_i(dst_ack_i)
	);
	// Trace: design.sv:73193:3
	generate
		if ((DataSrc2Dst == 1'b0) && (DataReg == 1'b1)) begin : gen_data_reg
			// Trace: design.sv:73194:5
			wire data_we;
			// Trace: design.sv:73195:5
			wire [Width - 1:0] data_d;
			reg [Width - 1:0] data_q;
			// Trace: design.sv:73198:5
			assign data_we = dst_req_o & dst_ack_i;
			// Trace: design.sv:73199:5
			assign data_d = data_i;
			// Trace: design.sv:73200:5
			always @(posedge clk_dst_i or negedge rst_dst_ni)
				// Trace: design.sv:73201:7
				if (!rst_dst_ni)
					// Trace: design.sv:73202:9
					data_q <= 1'sb0;
				else if (data_we)
					// Trace: design.sv:73204:9
					data_q <= data_d;
			// Trace: design.sv:73207:5
			assign data_o = data_q;
		end
		else begin : gen_no_data_reg
			// Trace: design.sv:73211:5
			assign data_o = data_i;
		end
	endgenerate
	// Trace: design.sv:73217:3
endmodule
module prim_sync_slow_fast (
	clk_slow_i,
	clk_fast_i,
	rst_fast_ni,
	wdata_i,
	rdata_o
);
	// Trace: design.sv:73252:13
	parameter [31:0] Width = 32;
	// Trace: design.sv:73254:3
	input wire clk_slow_i;
	// Trace: design.sv:73255:3
	input wire clk_fast_i;
	// Trace: design.sv:73256:3
	input wire rst_fast_ni;
	// Trace: design.sv:73257:3
	input wire [Width - 1:0] wdata_i;
	// Trace: design.sv:73258:3
	output wire [Width - 1:0] rdata_o;
	// Trace: design.sv:73261:3
	wire sync_clk_slow;
	reg sync_clk_slow_q;
	// Trace: design.sv:73262:3
	wire wdata_en;
	// Trace: design.sv:73263:3
	reg [Width - 1:0] wdata_q;
	// Trace: design.sv:73266:3
	prim_flop_2sync #(.Width(1)) sync_slow_clk(
		.clk_i(clk_fast_i),
		.rst_ni(rst_fast_ni),
		.d_i(clk_slow_i),
		.q_o(sync_clk_slow)
	);
	// Trace: design.sv:73273:3
	always @(posedge clk_fast_i or negedge rst_fast_ni)
		// Trace: design.sv:73274:5
		if (!rst_fast_ni)
			// Trace: design.sv:73275:7
			sync_clk_slow_q <= 1'b0;
		else
			// Trace: design.sv:73277:7
			sync_clk_slow_q <= sync_clk_slow;
	// Trace: design.sv:73282:3
	assign wdata_en = sync_clk_slow_q & !sync_clk_slow;
	// Trace: design.sv:73285:3
	always @(posedge clk_fast_i or negedge rst_fast_ni)
		// Trace: design.sv:73286:5
		if (!rst_fast_ni)
			// Trace: design.sv:73287:7
			wdata_q <= 1'sb0;
		else if (wdata_en)
			// Trace: design.sv:73289:7
			wdata_q <= wdata_i;
	// Trace: design.sv:73293:3
	assign rdata_o = wdata_q;
endmodule
module prim_keccak (
	rnd_i,
	s_i,
	s_o
);
	// Trace: design.sv:73303:13
	parameter signed [31:0] Width = 1600;
	// Trace: design.sv:73306:14
	localparam signed [31:0] W = Width / 25;
	// Trace: design.sv:73307:14
	localparam signed [31:0] L = $clog2(W);
	// Trace: design.sv:73308:14
	localparam signed [31:0] MaxRound = 12 + (2 * L);
	// Trace: design.sv:73309:14
	localparam signed [31:0] RndW = $clog2(MaxRound + 1);
	// Trace: design.sv:73311:3
	input [RndW - 1:0] rnd_i;
	// Trace: design.sv:73312:3
	input [Width - 1:0] s_i;
	// Trace: design.sv:73313:3
	output wire [Width - 1:0] s_o;
	// Trace: design.sv:73319:3
	// removed localparam type box_t
	// Trace: design.sv:73320:3
	// removed localparam type lane_t
	// Trace: design.sv:73321:3
	// removed localparam type plane_t
	// Trace: design.sv:73322:3
	// removed localparam type slice_t
	// Trace: design.sv:73323:3
	// removed localparam type sheet_t
	// Trace: design.sv:73324:3
	// removed localparam type row_t
	// Trace: design.sv:73325:3
	// removed localparam type col_t
	// Trace: design.sv:73330:3
	wire [(25 * W) - 1:0] state_in;
	wire [(25 * W) - 1:0] keccak_f;
	// Trace: design.sv:73331:3
	wire [(25 * W) - 1:0] theta_data;
	wire [(25 * W) - 1:0] rho_data;
	wire [(25 * W) - 1:0] pi_data;
	wire [(25 * W) - 1:0] chi_data;
	wire [(25 * W) - 1:0] iota_data;
	// Trace: design.sv:73332:3
	function automatic [(25 * W) - 1:0] bitarray_to_box;
		// Trace: design.sv:73384:44
		input reg [Width - 1:0] s_in;
		// Trace: design.sv:73385:5
		reg [(25 * W) - 1:0] box;
		begin
			// Trace: design.sv:73386:5
			begin : sv2v_autoblock_1
				// Trace: design.sv:73386:10
				reg signed [31:0] y;
				// Trace: design.sv:73386:10
				for (y = 0; y < 5; y = y + 1)
					begin
						// Trace: design.sv:73387:7
						begin : sv2v_autoblock_2
							// Trace: design.sv:73387:12
							reg signed [31:0] x;
							// Trace: design.sv:73387:12
							for (x = 0; x < 5; x = x + 1)
								begin
									// Trace: design.sv:73388:9
									begin : sv2v_autoblock_3
										// Trace: design.sv:73388:14
										reg signed [31:0] z;
										// Trace: design.sv:73388:14
										for (z = 0; z < W; z = z + 1)
											begin
												// Trace: design.sv:73389:11
												box[(((x * 5) + y) * W) + z] = s_in[(W * ((5 * y) + x)) + z];
											end
									end
								end
						end
					end
			end
			bitarray_to_box = box;
		end
	endfunction
	assign state_in = bitarray_to_box(s_i);
	// Trace: design.sv:73333:3
	function automatic [(25 * W) - 1:0] theta;
		// Trace: design.sv:73415:34
		input reg [(25 * W) - 1:0] state;
		// Trace: design.sv:73416:5
		reg [(5 * W) - 1:0] c;
		// Trace: design.sv:73417:5
		reg [(5 * W) - 1:0] d;
		// Trace: design.sv:73418:5
		reg [(25 * W) - 1:0] result;
		begin
			// Trace: design.sv:73419:5
			begin : sv2v_autoblock_4
				// Trace: design.sv:73419:10
				reg signed [31:0] x;
				// Trace: design.sv:73419:10
				for (x = 0; x < 5; x = x + 1)
					begin
						// Trace: design.sv:73420:7
						begin : sv2v_autoblock_5
							// Trace: design.sv:73420:12
							reg signed [31:0] z;
							// Trace: design.sv:73420:12
							for (z = 0; z < W; z = z + 1)
								begin
									// Trace: design.sv:73421:9
									c[(x * W) + z] = (((state[((x * 5) * W) + z] ^ state[(((x * 5) + 1) * W) + z]) ^ state[(((x * 5) + 2) * W) + z]) ^ state[(((x * 5) + 3) * W) + z]) ^ state[(((x * 5) + 4) * W) + z];
								end
						end
					end
			end
			begin : sv2v_autoblock_6
				// Trace: design.sv:73425:10
				reg signed [31:0] x;
				// Trace: design.sv:73425:10
				for (x = 0; x < 5; x = x + 1)
					begin : sv2v_autoblock_7
						// Trace: design.sv:73426:7
						reg signed [31:0] index_x1;
						reg signed [31:0] index_x2;
						// Trace: design.sv:73427:7
						index_x1 = (x == 0 ? 4 : x - 1);
						// Trace: design.sv:73428:7
						index_x2 = (x == 4 ? 0 : x + 1);
						// Trace: design.sv:73429:7
						begin : sv2v_autoblock_8
							// Trace: design.sv:73429:12
							reg signed [31:0] z;
							// Trace: design.sv:73429:12
							for (z = 0; z < W; z = z + 1)
								begin : sv2v_autoblock_9
									// Trace: design.sv:73430:9
									reg signed [31:0] index_z;
									// Trace: design.sv:73431:9
									index_z = (z == 0 ? W - 1 : z - 1);
									// Trace: design.sv:73432:9
									d[(x * W) + z] = c[(index_x1 * W) + z] ^ c[(index_x2 * W) + index_z];
								end
						end
					end
			end
			begin : sv2v_autoblock_10
				// Trace: design.sv:73435:10
				reg signed [31:0] x;
				// Trace: design.sv:73435:10
				for (x = 0; x < 5; x = x + 1)
					begin
						// Trace: design.sv:73436:7
						begin : sv2v_autoblock_11
							// Trace: design.sv:73436:12
							reg signed [31:0] y;
							// Trace: design.sv:73436:12
							for (y = 0; y < 5; y = y + 1)
								begin
									// Trace: design.sv:73437:9
									begin : sv2v_autoblock_12
										// Trace: design.sv:73437:14
										reg signed [31:0] z;
										// Trace: design.sv:73437:14
										for (z = 0; z < W; z = z + 1)
											begin
												// Trace: design.sv:73438:11
												result[(((x * 5) + y) * W) + z] = state[(((x * 5) + y) * W) + z] ^ d[(x * W) + z];
											end
									end
								end
						end
					end
			end
			theta = result;
		end
	endfunction
	assign theta_data = theta(state_in);
	// Trace: design.sv:73336:3
	localparam signed [799:0] PiRotate = 800'h30000000100000004000000020000000100000004000000020000000000000003000000020000000000000003000000010000000400000003000000010000000400000002000000000000000400000002000000000000000300000001;
	function automatic [(25 * W) - 1:0] pi;
		// Trace: design.sv:73494:31
		input reg [(25 * W) - 1:0] state;
		// Trace: design.sv:73495:5
		reg [(25 * W) - 1:0] result;
		begin
			// Trace: design.sv:73496:5
			begin : sv2v_autoblock_13
				// Trace: design.sv:73496:10
				reg signed [31:0] x;
				// Trace: design.sv:73496:10
				for (x = 0; x < 5; x = x + 1)
					begin
						// Trace: design.sv:73497:7
						begin : sv2v_autoblock_14
							// Trace: design.sv:73497:12
							reg signed [31:0] y;
							// Trace: design.sv:73497:12
							for (y = 0; y < 5; y = y + 1)
								begin : sv2v_autoblock_15
									// Trace: design.sv:73498:9
									reg signed [31:0] index_x;
									// Trace: design.sv:73499:9
									result[(((x * 5) + y) * W) + (W - 1)-:W] = state[(((PiRotate[(((4 - x) * 5) + (4 - y)) * 32+:32] * 5) + x) * W) + (W - 1)-:W];
								end
						end
					end
			end
			pi = result;
		end
	endfunction
	assign pi_data = pi(rho_data);
	// Trace: design.sv:73337:3
	function automatic [(25 * W) - 1:0] chi;
		// Trace: design.sv:73507:32
		input reg [(25 * W) - 1:0] state;
		// Trace: design.sv:73508:5
		reg [(25 * W) - 1:0] result;
		begin
			// Trace: design.sv:73509:5
			begin : sv2v_autoblock_16
				// Trace: design.sv:73509:10
				reg signed [31:0] x;
				// Trace: design.sv:73509:10
				for (x = 0; x < 5; x = x + 1)
					begin : sv2v_autoblock_17
						// Trace: design.sv:73510:7
						reg signed [31:0] index_x1;
						reg signed [31:0] index_x2;
						// Trace: design.sv:73511:7
						index_x1 = (x == 4 ? 0 : x + 1);
						// Trace: design.sv:73512:7
						index_x2 = (x >= 3 ? x - 3 : x + 2);
						// Trace: design.sv:73513:7
						begin : sv2v_autoblock_18
							// Trace: design.sv:73513:12
							reg signed [31:0] y;
							// Trace: design.sv:73513:12
							for (y = 0; y < 5; y = y + 1)
								begin
									// Trace: design.sv:73514:9
									begin : sv2v_autoblock_19
										// Trace: design.sv:73514:14
										reg signed [31:0] z;
										// Trace: design.sv:73514:14
										for (z = 0; z < W; z = z + 1)
											begin
												// Trace: design.sv:73515:11
												result[(((x * 5) + y) * W) + z] = state[(((x * 5) + y) * W) + z] ^ (~state[(((index_x1 * 5) + y) * W) + z] & state[(((index_x2 * 5) + y) * W) + z]);
											end
									end
								end
						end
					end
			end
			chi = result;
		end
	endfunction
	assign chi_data = chi(pi_data);
	// Trace: design.sv:73338:3
	localparam [1535:0] RC = 1536'h10000000000008082800000000000808a8000000080008000000000000000808b000000008000000180000000800080818000000000008009000000000000008a00000000000000880000000080008009000000008000000a000000008000808b800000000000008b8000000000008089800000000000800380000000000080028000000000000080000000000000800a800000008000000a8000000080008081800000000000808000000000800000018000000080008008;
	function automatic [(25 * W) - 1:0] iota;
		// Trace: design.sv:73571:33
		input reg [(25 * W) - 1:0] state;
		// Trace: design.sv:73571:46
		input reg [RndW - 1:0] rnd;
		// Trace: design.sv:73572:5
		reg [(25 * W) - 1:0] result;
		begin
			// Trace: design.sv:73573:5
			result = state;
			// Trace: design.sv:73574:5
			result[W - 1-:W] = state[W - 1-:W] ^ RC[((23 - rnd) * 64) + (W - 1)-:W];
			// Trace: design.sv:73576:5
			iota = result;
		end
	endfunction
	assign iota_data = iota(chi_data, rnd_i);
	// Trace: design.sv:73339:3
	assign keccak_f = iota_data;
	// Trace: design.sv:73340:3
	function automatic [Width - 1:0] box_to_bitarray;
		// Trace: design.sv:73397:56
		input reg [(25 * W) - 1:0] state;
		// Trace: design.sv:73398:5
		reg [Width - 1:0] bitarray;
		begin
			// Trace: design.sv:73399:5
			begin : sv2v_autoblock_20
				// Trace: design.sv:73399:10
				reg signed [31:0] y;
				// Trace: design.sv:73399:10
				for (y = 0; y < 5; y = y + 1)
					begin
						// Trace: design.sv:73400:7
						begin : sv2v_autoblock_21
							// Trace: design.sv:73400:12
							reg signed [31:0] x;
							// Trace: design.sv:73400:12
							for (x = 0; x < 5; x = x + 1)
								begin
									// Trace: design.sv:73401:9
									begin : sv2v_autoblock_22
										// Trace: design.sv:73401:14
										reg signed [31:0] z;
										// Trace: design.sv:73401:14
										for (z = 0; z < W; z = z + 1)
											begin
												// Trace: design.sv:73402:11
												bitarray[(W * ((5 * y) + x)) + z] = state[(((x * 5) + y) * W) + z];
											end
									end
								end
						end
					end
			end
			box_to_bitarray = bitarray;
		end
	endfunction
	assign s_o = box_to_bitarray(keccak_f);
	// Trace: design.sv:73345:3
	localparam signed [799:0] RhoOffset = 800'h240000000300000069000000d2000000010000012c0000000a0000002d00000042000000be00000006000000ab0000000f000000fd0000001c000000370000009900000015000000780000005b00000114000000e7000000880000004e;
	// Trace: design.sv:73353:3
	genvar _gv_x_1;
	generate
		for (_gv_x_1 = 0; _gv_x_1 < 5; _gv_x_1 = _gv_x_1 + 1) begin : gen_rho_x
			localparam x = _gv_x_1;
			genvar _gv_y_1;
			for (_gv_y_1 = 0; _gv_y_1 < 5; _gv_y_1 = _gv_y_1 + 1) begin : gen_rho_y
				localparam y = _gv_y_1;
				// Trace: design.sv:73355:7
				localparam signed [31:0] Offset = RhoOffset[(((4 - x) * 5) + (4 - y)) * 32+:32] % W;
				// Trace: design.sv:73356:7
				localparam signed [31:0] ShiftAmt = W - Offset;
				if (Offset == 0) begin : gen_offset0
					// Trace: design.sv:73358:9
					assign rho_data[(((x * 5) + y) * W) + (W - 1)-:W] = theta_data[(((x * 5) + y) * W) + (W - 1)-:W];
				end
				else begin : gen_others
					// Trace: design.sv:73360:9
					assign rho_data[(((x * 5) + y) * W) + (W - 1)-:W] = {theta_data[((x * 5) + y) * W+:ShiftAmt], theta_data[(((x * 5) + y) * W) + ShiftAmt+:Offset]};
				end
			end
		end
	endgenerate
	// Trace: design.sv:73384:3
	// Trace: design.sv:73397:3
	// Trace: design.sv:73415:3
	// Trace: design.sv:73486:3
	// Trace: design.sv:73494:3
	// Trace: design.sv:73507:3
	// Trace: design.sv:73543:3
	// Trace: design.sv:73571:3
endmodule
module prim_packer (
	clk_i,
	rst_ni,
	valid_i,
	data_i,
	mask_i,
	ready_o,
	valid_o,
	data_o,
	mask_o,
	ready_i,
	flush_i,
	flush_done_o
);
	reg _sv2v_0;
	// Trace: design.sv:73600:13
	parameter signed [31:0] InW = 32;
	// Trace: design.sv:73601:13
	parameter signed [31:0] OutW = 32;
	// Trace: design.sv:73602:13
	parameter signed [31:0] HintByteData = 0;
	// Trace: design.sv:73604:3
	input clk_i;
	// Trace: design.sv:73605:3
	input rst_ni;
	// Trace: design.sv:73607:3
	input valid_i;
	// Trace: design.sv:73608:3
	input [InW - 1:0] data_i;
	// Trace: design.sv:73609:3
	input [InW - 1:0] mask_i;
	// Trace: design.sv:73610:3
	output wire ready_o;
	// Trace: design.sv:73612:3
	output wire valid_o;
	// Trace: design.sv:73613:3
	output wire [OutW - 1:0] data_o;
	// Trace: design.sv:73614:3
	output wire [OutW - 1:0] mask_o;
	// Trace: design.sv:73615:3
	input ready_i;
	// Trace: design.sv:73617:3
	input flush_i;
	// Trace: design.sv:73618:3
	output wire flush_done_o;
	// Trace: design.sv:73621:3
	localparam signed [31:0] Width = InW + OutW;
	// Trace: design.sv:73622:3
	localparam signed [31:0] ConcatW = Width + InW;
	// Trace: design.sv:73623:3
	localparam signed [31:0] PtrW = $clog2(ConcatW + 1);
	// Trace: design.sv:73624:3
	localparam signed [31:0] IdxW = $clog2(InW) + ~|$clog2(InW);
	// Trace: design.sv:73626:3
	wire valid_next;
	wire ready_next;
	// Trace: design.sv:73627:3
	reg [Width - 1:0] stored_data;
	reg [Width - 1:0] stored_mask;
	// Trace: design.sv:73628:3
	wire [ConcatW - 1:0] concat_data;
	wire [ConcatW - 1:0] concat_mask;
	// Trace: design.sv:73629:3
	wire [ConcatW - 1:0] shiftl_data;
	wire [ConcatW - 1:0] shiftl_mask;
	// Trace: design.sv:73631:3
	reg [PtrW - 1:0] pos;
	reg [PtrW - 1:0] pos_next;
	// Trace: design.sv:73632:3
	reg [IdxW - 1:0] lod_idx;
	// Trace: design.sv:73633:3
	reg [$clog2(InW + 1) - 1:0] inmask_ones;
	// Trace: design.sv:73635:3
	wire ack_in;
	wire ack_out;
	// Trace: design.sv:73637:3
	reg flush_valid;
	// Trace: design.sv:73638:3
	reg flush_done;
	// Trace: design.sv:73641:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:73643:5
		inmask_ones = 1'sb0;
		// Trace: design.sv:73644:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:73644:10
			reg signed [31:0] i;
			// Trace: design.sv:73644:10
			for (i = 0; i < InW; i = i + 1)
				begin
					// Trace: design.sv:73645:7
					inmask_ones = inmask_ones + mask_i[i];
				end
		end
	end
	// Trace: design.sv:73649:3
	reg [PtrW - 1:0] pos_with_input;
	// Trace: design.sv:73651:3
	function automatic [PtrW - 1:0] sv2v_cast_09B00;
		input reg [PtrW - 1:0] inp;
		sv2v_cast_09B00 = inp;
	endfunction
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:73652:5
		pos_next = pos;
		// Trace: design.sv:73653:5
		pos_with_input = pos + sv2v_cast_09B00(inmask_ones);
		// Trace: design.sv:73655:5
		(* full_case, parallel_case *)
		case ({ack_in, ack_out})
			2'b00:
				// Trace: design.sv:73656:14
				pos_next = pos;
			2'b01:
				// Trace: design.sv:73657:14
				pos_next = (pos <= OutW ? {PtrW {1'sb0}} : pos - OutW);
			2'b10:
				// Trace: design.sv:73658:14
				pos_next = pos_with_input;
			2'b11:
				// Trace: design.sv:73659:14
				pos_next = (pos_with_input <= OutW ? {PtrW {1'sb0}} : pos_with_input - OutW);
			default:
				// Trace: design.sv:73660:16
				pos_next = pos;
		endcase
	end
	// Trace: design.sv:73664:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:73665:5
		if (!rst_ni)
			// Trace: design.sv:73666:7
			pos <= 1'sb0;
		else if (flush_done)
			// Trace: design.sv:73668:7
			pos <= 1'sb0;
		else
			// Trace: design.sv:73670:7
			pos <= pos_next;
	// Trace: design.sv:73676:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:73677:5
		lod_idx = 0;
		// Trace: design.sv:73678:5
		begin : sv2v_autoblock_2
			// Trace: design.sv:73678:10
			reg signed [31:0] i;
			// Trace: design.sv:73678:10
			for (i = InW - 1; i >= 0; i = i - 1)
				begin
					// Trace: design.sv:73679:7
					if (mask_i[i] == 1'b1)
						// Trace: design.sv:73680:9
						lod_idx = $unsigned(i);
				end
		end
	end
	// Trace: design.sv:73685:3
	assign ack_in = valid_i & ready_o;
	// Trace: design.sv:73686:3
	assign ack_out = valid_o & ready_i;
	// Trace: design.sv:73690:3
	function automatic [Width - 1:0] sv2v_cast_62596;
		input reg [Width - 1:0] inp;
		sv2v_cast_62596 = inp;
	endfunction
	assign shiftl_data = (valid_i ? sv2v_cast_62596(data_i >> lod_idx) << pos : {ConcatW {1'sb0}});
	// Trace: design.sv:73691:3
	assign shiftl_mask = (valid_i ? sv2v_cast_62596(mask_i >> lod_idx) << pos : {ConcatW {1'sb0}});
	// Trace: design.sv:73694:3
	assign concat_data = {{InW {1'b0}}, stored_data & stored_mask} | (shiftl_data & shiftl_mask);
	// Trace: design.sv:73696:3
	assign concat_mask = {{InW {1'b0}}, stored_mask} | shiftl_mask;
	// Trace: design.sv:73698:3
	reg [Width - 1:0] stored_data_next;
	reg [Width - 1:0] stored_mask_next;
	// Trace: design.sv:73700:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:73701:5
		(* full_case, parallel_case *)
		case ({ack_in, ack_out})
			2'b00: begin
				// Trace: design.sv:73703:9
				stored_data_next = stored_data;
				// Trace: design.sv:73704:9
				stored_mask_next = stored_mask;
			end
			2'b01: begin
				// Trace: design.sv:73708:9
				stored_data_next = {{OutW {1'b0}}, stored_data[Width - 1:OutW]};
				// Trace: design.sv:73709:9
				stored_mask_next = {{OutW {1'b0}}, stored_mask[Width - 1:OutW]};
			end
			2'b10: begin
				// Trace: design.sv:73713:9
				stored_data_next = concat_data[0+:Width];
				// Trace: design.sv:73714:9
				stored_mask_next = concat_mask[0+:Width];
			end
			2'b11: begin
				// Trace: design.sv:73718:9
				stored_data_next = concat_data[ConcatW - 1:OutW];
				// Trace: design.sv:73719:9
				stored_mask_next = concat_mask[ConcatW - 1:OutW];
			end
			default: begin
				// Trace: design.sv:73722:9
				stored_data_next = stored_data;
				// Trace: design.sv:73723:9
				stored_mask_next = stored_mask;
			end
		endcase
	end
	// Trace: design.sv:73729:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:73730:5
		if (!rst_ni) begin
			// Trace: design.sv:73731:7
			stored_data <= 1'sb0;
			// Trace: design.sv:73732:7
			stored_mask <= 1'sb0;
		end
		else if (flush_done) begin
			// Trace: design.sv:73734:7
			stored_data <= 1'sb0;
			// Trace: design.sv:73735:7
			stored_mask <= 1'sb0;
		end
		else begin
			// Trace: design.sv:73737:7
			stored_data <= stored_data_next;
			// Trace: design.sv:73738:7
			stored_mask <= stored_mask_next;
		end
	// Trace: design.sv:73744:3
	// removed localparam type flush_st_e
	// Trace: design.sv:73748:3
	reg flush_st;
	reg flush_st_next;
	// Trace: design.sv:73750:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:73751:5
		if (!rst_ni)
			// Trace: design.sv:73752:7
			flush_st <= 1'd0;
		else
			// Trace: design.sv:73754:7
			flush_st <= flush_st_next;
	// Trace: design.sv:73758:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:73759:5
		flush_st_next = 1'd0;
		// Trace: design.sv:73761:5
		flush_valid = 1'b0;
		// Trace: design.sv:73762:5
		flush_done = 1'b0;
		// Trace: design.sv:73764:5
		(* full_case, parallel_case *)
		case (flush_st)
			1'd0:
				// Trace: design.sv:73766:9
				if (flush_i)
					// Trace: design.sv:73767:11
					flush_st_next = 1'd1;
				else
					// Trace: design.sv:73769:11
					flush_st_next = 1'd0;
			1'd1:
				// Trace: design.sv:73774:9
				if (pos == {PtrW {1'sb0}}) begin
					// Trace: design.sv:73775:11
					flush_st_next = 1'd0;
					// Trace: design.sv:73777:11
					flush_valid = 1'b0;
					// Trace: design.sv:73778:11
					flush_done = 1'b1;
				end
				else begin
					// Trace: design.sv:73780:11
					flush_st_next = 1'd1;
					// Trace: design.sv:73782:11
					flush_valid = 1'b1;
					// Trace: design.sv:73783:11
					flush_done = 1'b0;
				end
			default: begin
				// Trace: design.sv:73787:9
				flush_st_next = 1'd0;
				// Trace: design.sv:73789:9
				flush_valid = 1'b0;
				// Trace: design.sv:73790:9
				flush_done = 1'b0;
			end
		endcase
	end
	// Trace: design.sv:73795:3
	assign flush_done_o = flush_done;
	// Trace: design.sv:73799:3
	assign valid_next = (pos >= OutW ? 1'b1 : flush_valid);
	// Trace: design.sv:73807:3
	assign ready_next = pos <= OutW;
	// Trace: design.sv:73810:3
	assign valid_o = valid_next;
	// Trace: design.sv:73811:3
	assign data_o = stored_data[OutW - 1:0];
	// Trace: design.sv:73812:3
	assign mask_o = stored_mask[OutW - 1:0];
	// Trace: design.sv:73815:3
	assign ready_o = ready_next;
	// Trace: design.sv:73824:3
	// Trace: design.sv:73871:3
	generate
		if (HintByteData != 0) begin : g_byte_assert
			genvar _gv_i_85;
			genvar _gv_i_86;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
module prim_packer_fifo (
	clk_i,
	rst_ni,
	clr_i,
	wvalid_i,
	wdata_i,
	wready_o,
	rvalid_o,
	rdata_o,
	rready_i,
	depth_o
);
	// Trace: design.sv:73932:13
	parameter signed [31:0] InW = 32;
	// Trace: design.sv:73933:13
	parameter signed [31:0] OutW = 8;
	// Trace: design.sv:73935:14
	localparam signed [31:0] MaxW = (InW > OutW ? InW : OutW);
	// Trace: design.sv:73936:14
	localparam signed [31:0] MinW = (InW < OutW ? InW : OutW);
	// Trace: design.sv:73937:14
	localparam signed [31:0] DepthW = $clog2(MaxW / MinW);
	// Trace: design.sv:73939:3
	input wire clk_i;
	// Trace: design.sv:73940:3
	input wire rst_ni;
	// Trace: design.sv:73942:3
	input wire clr_i;
	// Trace: design.sv:73943:3
	input wire wvalid_i;
	// Trace: design.sv:73944:3
	input wire [InW - 1:0] wdata_i;
	// Trace: design.sv:73945:3
	output wire wready_o;
	// Trace: design.sv:73947:3
	output wire rvalid_o;
	// Trace: design.sv:73948:3
	output wire [OutW - 1:0] rdata_o;
	// Trace: design.sv:73949:3
	input wire rready_i;
	// Trace: design.sv:73950:3
	output wire [DepthW:0] depth_o;
	// Trace: design.sv:73953:3
	localparam [31:0] WidthRatio = MaxW / MinW;
	// Trace: design.sv:73954:3
	localparam [DepthW:0] FullDepth = WidthRatio[DepthW:0];
	// Trace: design.sv:73957:3
	wire load_data;
	// Trace: design.sv:73958:3
	wire clear_data;
	// Trace: design.sv:73961:3
	reg [DepthW:0] depth_q;
	wire [DepthW:0] depth_d;
	// Trace: design.sv:73962:3
	reg [MaxW - 1:0] data_q;
	wire [MaxW - 1:0] data_d;
	// Trace: design.sv:73963:3
	reg clr_q;
	wire clr_d;
	// Trace: design.sv:73965:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:73966:5
		if (!rst_ni) begin
			// Trace: design.sv:73967:7
			depth_q <= 1'sb0;
			// Trace: design.sv:73968:7
			data_q <= 1'sb0;
			// Trace: design.sv:73969:7
			clr_q <= 1'b1;
		end
		else begin
			// Trace: design.sv:73971:7
			depth_q <= depth_d;
			// Trace: design.sv:73972:7
			data_q <= data_d;
			// Trace: design.sv:73973:7
			clr_q <= clr_d;
		end
	// Trace: design.sv:73978:3
	assign clr_d = clr_i;
	// Trace: design.sv:73980:3
	assign depth_o = depth_q;
	// Trace: design.sv:73982:3
	generate
		if (InW < OutW) begin : gen_pack_mode
			// Trace: design.sv:73983:5
			wire [MaxW - 1:0] wdata_shifted;
			// Trace: design.sv:73985:5
			assign wdata_shifted = {{OutW - InW {1'b0}}, wdata_i} << (depth_q * InW);
			// Trace: design.sv:73986:5
			assign clear_data = (rready_i && rvalid_o) || clr_q;
			// Trace: design.sv:73987:5
			assign load_data = wvalid_i && wready_o;
			// Trace: design.sv:73989:5
			assign depth_d = (clear_data ? {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}} : (load_data ? depth_q + 1 : depth_q));
			// Trace: design.sv:73993:5
			assign data_d = (clear_data ? {MaxW {1'sb0}} : (load_data ? data_q | wdata_shifted : data_q));
			// Trace: design.sv:73998:5
			assign wready_o = (depth_q != FullDepth) && !clr_q;
			// Trace: design.sv:73999:5
			assign rdata_o = data_q;
			// Trace: design.sv:74000:5
			assign rvalid_o = (depth_q == FullDepth) && !clr_q;
		end
		else begin : gen_unpack_mode
			// Trace: design.sv:74003:5
			wire [MaxW - 1:0] rdata_shifted;
			// Trace: design.sv:74004:5
			wire pull_data;
			// Trace: design.sv:74005:5
			reg [DepthW:0] ptr_q;
			wire [DepthW:0] ptr_d;
			// Trace: design.sv:74006:5
			wire [DepthW:0] lsb_is_one;
			// Trace: design.sv:74007:5
			wire [DepthW:0] max_value;
			// Trace: design.sv:74009:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:74010:7
				if (!rst_ni)
					// Trace: design.sv:74011:9
					ptr_q <= 1'sb0;
				else
					// Trace: design.sv:74013:9
					ptr_q <= ptr_d;
			// Trace: design.sv:74017:5
			assign lsb_is_one = {{DepthW {1'b0}}, 1'b1};
			// Trace: design.sv:74018:5
			assign max_value = FullDepth;
			// Trace: design.sv:74019:5
			assign rdata_shifted = data_q >> (ptr_q * OutW);
			// Trace: design.sv:74020:5
			assign clear_data = (rready_i && (depth_q == lsb_is_one)) || clr_q;
			// Trace: design.sv:74021:5
			assign load_data = wvalid_i && wready_o;
			// Trace: design.sv:74022:5
			assign pull_data = rvalid_o && rready_i;
			// Trace: design.sv:74024:5
			assign depth_d = (clear_data ? {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}} : (load_data ? max_value : (pull_data ? depth_q - 1 : depth_q)));
			// Trace: design.sv:74029:5
			assign ptr_d = (clear_data ? {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}} : (pull_data ? ptr_q + 1 : ptr_q));
			// Trace: design.sv:74033:5
			assign data_d = (clear_data ? {MaxW {1'sb0}} : (load_data ? wdata_i : data_q));
			// Trace: design.sv:74038:5
			assign wready_o = (depth_q == {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}}) && !clr_q;
			// Trace: design.sv:74039:5
			assign rdata_o = rdata_shifted[OutW - 1:0];
			// Trace: design.sv:74040:5
			assign rvalid_o = (depth_q != {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}}) && !clr_q;
			if (InW > OutW) begin : gen_unused
				// Trace: design.sv:74044:7
				wire [(MaxW - MinW) - 1:0] unused_rdata_shifted;
				// Trace: design.sv:74045:7
				assign unused_rdata_shifted = rdata_shifted[MaxW - 1:MinW];
			end
		end
	endgenerate
endmodule
module prim_gate_gen (
	clk_i,
	rst_ni,
	valid_i,
	data_i,
	data_o,
	valid_o
);
	// Trace: design.sv:74099:13
	parameter signed [31:0] DataWidth = 32;
	// Trace: design.sv:74100:13
	parameter signed [31:0] NumGates = 1000;
	// Trace: design.sv:74102:3
	input clk_i;
	// Trace: design.sv:74103:3
	input rst_ni;
	// Trace: design.sv:74105:3
	input valid_i;
	// Trace: design.sv:74106:3
	input [DataWidth - 1:0] data_i;
	// Trace: design.sv:74107:3
	output wire [DataWidth - 1:0] data_o;
	// Trace: design.sv:74108:3
	output wire valid_o;
	// Trace: design.sv:74117:3
	localparam signed [31:0] NumInnerRounds = 2;
	// Trace: design.sv:74118:3
	localparam signed [31:0] GatesPerRound = DataWidth * 14;
	// Trace: design.sv:74120:3
	localparam signed [31:0] NumOuterRounds = (NumGates + (GatesPerRound / 2)) / GatesPerRound;
	// Trace: design.sv:74130:3
	wire [(NumOuterRounds * DataWidth) - 1:0] regs_d;
	reg [(NumOuterRounds * DataWidth) - 1:0] regs_q;
	// Trace: design.sv:74131:3
	wire [NumOuterRounds - 1:0] valid_d;
	reg [NumOuterRounds - 1:0] valid_q;
	// Trace: design.sv:74133:3
	genvar _gv_k_14;
	localparam [63:0] prim_cipher_pkg_PRINCE_SBOX4 = 64'h4d5e087619ca23fb;
	function automatic [7:0] prim_cipher_pkg_sbox4_8bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:325:45
		input reg [7:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:325:67
		input reg [63:0] sbox4;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:326:5
		reg [7:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:5
			begin : sv2v_autoblock_1
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:328:10
				for (k = 0; k < 2; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:329:7
						state_out[k * 4+:4] = sbox4[state_in[k * 4+:4] * 4+:4];
					end
			end
			prim_cipher_pkg_sbox4_8bit = state_out;
		end
	endfunction
	function automatic [31:0] prim_cipher_pkg_sbox4_32bit;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:343:47
		input reg [31:0] state_in;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:343:70
		input reg [63:0] sbox4;
		// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:344:5
		reg [31:0] state_out;
		begin
			// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:5
			begin : sv2v_autoblock_2
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:10
				reg signed [31:0] k;
				// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:346:10
				for (k = 0; k < 4; k = k + 1)
					begin
						// Trace: ../src/lowrisc_prim_cipher_pkg_0.1/rtl/prim_cipher_pkg.sv:347:7
						state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
					end
			end
			prim_cipher_pkg_sbox4_32bit = state_out;
		end
	endfunction
	generate
		for (_gv_k_14 = 0; _gv_k_14 < NumOuterRounds; _gv_k_14 = _gv_k_14 + 1) begin : gen_outer_round
			localparam k = _gv_k_14;
			// Trace: design.sv:74135:5
			wire [(3 * DataWidth) - 1:0] inner_data;
			if (k == 0) begin : gen_first
				// Trace: design.sv:74138:7
				assign inner_data[0+:DataWidth] = data_i;
				// Trace: design.sv:74139:7
				assign valid_d[0] = valid_i;
			end
			else begin : gen_others
				// Trace: design.sv:74141:7
				assign inner_data[0+:DataWidth] = regs_q[(k - 1) * DataWidth+:DataWidth];
				// Trace: design.sv:74142:7
				assign valid_d[k] = valid_q[k - 1];
			end
			genvar _gv_l_7;
			for (_gv_l_7 = 0; _gv_l_7 < NumInnerRounds; _gv_l_7 = _gv_l_7 + 1) begin : gen_inner
				localparam l = _gv_l_7;
				// Trace: design.sv:74147:7
				assign inner_data[(l + 1) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_32bit({inner_data[(l * DataWidth) + 1-:2], inner_data[(l * DataWidth) + ((DataWidth - 1) >= 2 ? DataWidth - 1 : ((DataWidth - 1) + ((DataWidth - 1) >= 2 ? DataWidth - 2 : 4 - DataWidth)) - 1)-:((DataWidth - 1) >= 2 ? DataWidth - 2 : 4 - DataWidth)]}, prim_cipher_pkg_PRINCE_SBOX4);
			end
			// Trace: design.sv:74152:5
			assign regs_d[k * DataWidth+:DataWidth] = inner_data[NumInnerRounds * DataWidth+:DataWidth];
		end
	endgenerate
	// Trace: design.sv:74155:3
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: design.sv:74156:5
		if (!rst_ni) begin
			// Trace: design.sv:74157:7
			regs_q <= 1'sb0;
			// Trace: design.sv:74158:7
			valid_q <= 1'sb0;
		end
		else begin
			// Trace: design.sv:74160:7
			valid_q <= valid_d;
			// Trace: design.sv:74161:7
			begin : sv2v_autoblock_3
				// Trace: design.sv:74161:12
				reg signed [31:0] k;
				// Trace: design.sv:74161:12
				for (k = 0; k < NumOuterRounds; k = k + 1)
					begin
						// Trace: design.sv:74162:9
						if (valid_d[k])
							// Trace: design.sv:74163:11
							regs_q[k * DataWidth+:DataWidth] <= regs_d[k * DataWidth+:DataWidth];
					end
			end
		end
	end
	// Trace: design.sv:74169:3
	assign data_o = regs_q[(NumOuterRounds - 1) * DataWidth+:DataWidth];
	// Trace: design.sv:74170:3
	assign valid_o = valid_q[NumOuterRounds - 1];
endmodule
module prim_pulse_sync (
	clk_src_i,
	rst_src_ni,
	src_pulse_i,
	clk_dst_i,
	rst_dst_ni,
	dst_pulse_o
);
	// Trace: design.sv:74185:3
	input wire clk_src_i;
	// Trace: design.sv:74186:3
	input wire rst_src_ni;
	// Trace: design.sv:74187:3
	input wire src_pulse_i;
	// Trace: design.sv:74189:3
	input wire clk_dst_i;
	// Trace: design.sv:74190:3
	input wire rst_dst_ni;
	// Trace: design.sv:74191:3
	output wire dst_pulse_o;
	// Trace: design.sv:74197:3
	reg src_level;
	// Trace: design.sv:74199:3
	always @(posedge clk_src_i or negedge rst_src_ni)
		// Trace: design.sv:74200:5
		if (!rst_src_ni)
			// Trace: design.sv:74201:7
			src_level <= 1'b0;
		else
			// Trace: design.sv:74203:7
			src_level <= src_level ^ src_pulse_i;
	// Trace: design.sv:74210:3
	wire dst_level;
	// Trace: design.sv:74212:3
	prim_flop_2sync #(.Width(1)) prim_flop_2sync(
		.d_i(src_level),
		.clk_i(clk_dst_i),
		.rst_ni(rst_dst_ni),
		.q_o(dst_level)
	);
	// Trace: design.sv:74224:3
	reg dst_level_q;
	// Trace: design.sv:74227:3
	always @(posedge clk_dst_i or negedge rst_dst_ni)
		// Trace: design.sv:74228:5
		if (!rst_dst_ni)
			// Trace: design.sv:74229:7
			dst_level_q <= 1'b0;
		else
			// Trace: design.sv:74231:7
			dst_level_q <= dst_level;
	// Trace: design.sv:74236:3
	assign dst_pulse_o = dst_level_q ^ dst_level;
endmodule
module prim_filter (
	clk_i,
	rst_ni,
	enable_i,
	filter_i,
	filter_o
);
	// Trace: design.sv:74251:32
	parameter signed [31:0] Cycles = 4;
	// Trace: design.sv:74252:3
	input clk_i;
	// Trace: design.sv:74253:3
	input rst_ni;
	// Trace: design.sv:74254:3
	input enable_i;
	// Trace: design.sv:74255:3
	input filter_i;
	// Trace: design.sv:74256:3
	output wire filter_o;
	// Trace: design.sv:74259:3
	reg [Cycles - 1:0] stored_vector_q;
	wire [Cycles - 1:0] stored_vector_d;
	// Trace: design.sv:74260:3
	reg stored_value_q;
	wire update_stored_value;
	// Trace: design.sv:74261:3
	wire unused_stored_vector_q_msb;
	// Trace: design.sv:74263:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:74264:5
		if (!rst_ni)
			// Trace: design.sv:74265:7
			stored_value_q <= 1'b0;
		else if (update_stored_value)
			// Trace: design.sv:74267:7
			stored_value_q <= filter_i;
	// Trace: design.sv:74271:3
	assign stored_vector_d = {stored_vector_q[Cycles - 2:0], filter_i};
	// Trace: design.sv:74272:3
	assign unused_stored_vector_q_msb = stored_vector_q[Cycles - 1];
	// Trace: design.sv:74274:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:74275:5
		if (!rst_ni)
			// Trace: design.sv:74276:7
			stored_vector_q <= {Cycles {1'b0}};
		else
			// Trace: design.sv:74278:7
			stored_vector_q <= stored_vector_d;
	// Trace: design.sv:74282:3
	assign update_stored_value = (stored_vector_d == {Cycles {1'b0}}) | (stored_vector_d == {Cycles {1'b1}});
	// Trace: design.sv:74286:3
	assign filter_o = (enable_i ? stored_value_q : filter_i);
endmodule
module prim_filter_ctr (
	clk_i,
	rst_ni,
	enable_i,
	filter_i,
	filter_o
);
	// Trace: design.sv:74304:36
	parameter [31:0] Cycles = 4;
	// Trace: design.sv:74305:3
	input clk_i;
	// Trace: design.sv:74306:3
	input rst_ni;
	// Trace: design.sv:74307:3
	input enable_i;
	// Trace: design.sv:74308:3
	input filter_i;
	// Trace: design.sv:74309:3
	output wire filter_o;
	// Trace: design.sv:74312:3
	localparam [31:0] CTR_WIDTH = $clog2(Cycles);
	// Trace: design.sv:74313:3
	function automatic [CTR_WIDTH - 1:0] sv2v_cast_A7990;
		input reg [CTR_WIDTH - 1:0] inp;
		sv2v_cast_A7990 = inp;
	endfunction
	localparam [CTR_WIDTH - 1:0] CYCLESM1 = sv2v_cast_A7990(Cycles - 1);
	// Trace: design.sv:74315:3
	reg [CTR_WIDTH - 1:0] diff_ctr_q;
	wire [CTR_WIDTH - 1:0] diff_ctr_d;
	// Trace: design.sv:74316:3
	reg filter_q;
	reg stored_value_q;
	wire update_stored_value;
	// Trace: design.sv:74318:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:74319:5
		if (!rst_ni)
			// Trace: design.sv:74320:7
			filter_q <= 1'b0;
		else
			// Trace: design.sv:74322:7
			filter_q <= filter_i;
	// Trace: design.sv:74326:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:74327:5
		if (!rst_ni)
			// Trace: design.sv:74328:7
			stored_value_q <= 1'b0;
		else if (update_stored_value)
			// Trace: design.sv:74330:7
			stored_value_q <= filter_i;
	// Trace: design.sv:74334:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:74335:5
		if (!rst_ni)
			// Trace: design.sv:74336:7
			diff_ctr_q <= {CTR_WIDTH {1'b0}};
		else
			// Trace: design.sv:74338:7
			diff_ctr_q <= diff_ctr_d;
	// Trace: design.sv:74343:3
	assign diff_ctr_d = (filter_i != filter_q ? {CTR_WIDTH {1'sb0}} : (diff_ctr_q == CYCLESM1 ? CYCLESM1 : diff_ctr_q + 1'b1));
	// Trace: design.sv:74347:3
	assign update_stored_value = diff_ctr_d == CYCLESM1;
	// Trace: design.sv:74349:3
	assign filter_o = (enable_i ? stored_value_q : filter_i);
endmodule
module prim_intr_hw (
	clk_i,
	rst_ni,
	event_intr_i,
	reg2hw_intr_enable_q_i,
	reg2hw_intr_test_q_i,
	reg2hw_intr_test_qe_i,
	reg2hw_intr_state_q_i,
	hw2reg_intr_state_de_o,
	hw2reg_intr_state_d_o,
	intr_o
);
	// Trace: design.sv:74363:13
	parameter [31:0] Width = 1;
	// Trace: design.sv:74364:13
	parameter [0:0] FlopOutput = 1;
	// Trace: design.sv:74367:3
	input clk_i;
	// Trace: design.sv:74368:3
	input rst_ni;
	// Trace: design.sv:74369:3
	input [Width - 1:0] event_intr_i;
	// Trace: design.sv:74372:3
	input [Width - 1:0] reg2hw_intr_enable_q_i;
	// Trace: design.sv:74373:3
	input [Width - 1:0] reg2hw_intr_test_q_i;
	// Trace: design.sv:74374:3
	input reg2hw_intr_test_qe_i;
	// Trace: design.sv:74375:3
	input [Width - 1:0] reg2hw_intr_state_q_i;
	// Trace: design.sv:74376:3
	output wire hw2reg_intr_state_de_o;
	// Trace: design.sv:74377:3
	output wire [Width - 1:0] hw2reg_intr_state_d_o;
	// Trace: design.sv:74380:3
	output reg [Width - 1:0] intr_o;
	// Trace: design.sv:74383:3
	wire [Width - 1:0] new_event;
	// Trace: design.sv:74384:3
	assign new_event = ({Width {reg2hw_intr_test_qe_i}} & reg2hw_intr_test_q_i) | event_intr_i;
	// Trace: design.sv:74386:3
	assign hw2reg_intr_state_de_o = |new_event;
	// Trace: design.sv:74389:3
	assign hw2reg_intr_state_d_o = new_event | reg2hw_intr_state_q_i;
	// Trace: design.sv:74391:3
	generate
		if (FlopOutput == 1) begin : gen_flop_intr_output
			// Trace: design.sv:74393:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:74394:7
				if (!rst_ni)
					// Trace: design.sv:74395:9
					intr_o <= 1'sb0;
				else
					// Trace: design.sv:74397:9
					intr_o <= reg2hw_intr_state_q_i & reg2hw_intr_enable_q_i;
		end
		else begin : gen_intr_passthrough_output
			// Trace: design.sv:74402:5
			wire unused_clk;
			// Trace: design.sv:74403:5
			wire unused_rst_n;
			// Trace: design.sv:74404:5
			assign unused_clk = clk_i;
			// Trace: design.sv:74405:5
			assign unused_rst_n = rst_ni;
			// Trace: design.sv:74406:5
			wire [Width:1] sv2v_tmp_4934E;
			assign sv2v_tmp_4934E = reg2hw_intr_state_q_i & reg2hw_intr_enable_q_i;
			always @(*) intr_o = sv2v_tmp_4934E;
		end
	endgenerate
endmodule
module tlul_fifo_sync (
	clk_i,
	rst_ni,
	tl_h_i,
	tl_h_o,
	tl_d_o,
	tl_d_i,
	spare_req_i,
	spare_req_o,
	spare_rsp_i,
	spare_rsp_o
);
	// Trace: design.sv:74420:13
	parameter [0:0] ReqPass = 1'b1;
	// Trace: design.sv:74421:13
	parameter [0:0] RspPass = 1'b1;
	// Trace: design.sv:74422:13
	parameter [31:0] ReqDepth = 2;
	// Trace: design.sv:74423:13
	parameter [31:0] RspDepth = 2;
	// Trace: design.sv:74424:13
	parameter [31:0] SpareReqW = 1;
	// Trace: design.sv:74425:13
	parameter [31:0] SpareRspW = 1;
	// Trace: design.sv:74427:3
	input clk_i;
	// Trace: design.sv:74428:3
	input rst_ni;
	// Trace: design.sv:74429:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_h_i;
	// Trace: design.sv:74430:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o;
	// Trace: design.sv:74431:3
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_d_o;
	// Trace: design.sv:74432:3
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d_i;
	// Trace: design.sv:74433:3
	input [SpareReqW - 1:0] spare_req_i;
	// Trace: design.sv:74434:3
	output wire [SpareReqW - 1:0] spare_req_o;
	// Trace: design.sv:74435:3
	input [SpareRspW - 1:0] spare_rsp_i;
	// Trace: design.sv:74436:3
	output wire [SpareRspW - 1:0] spare_rsp_o;
	// Trace: design.sv:74440:3
	localparam [31:0] REQFIFO_WIDTH = ((1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)) - 2) + SpareReqW;
	// Trace: design.sv:74441:3
	wire [2:0] reqfifo_tl_d_a_opcode;
	// Trace: design.sv:74443:3
	assign tl_d_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] = reqfifo_tl_d_a_opcode;
	// Trace: design.sv:74445:3
	prim_fifo_sync #(
		.Width(REQFIFO_WIDTH),
		.Pass(ReqPass),
		.Depth(ReqDepth)
	) reqfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(tl_h_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))]),
		.wready_o(tl_h_o[0]),
		.wdata_i({tl_h_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)], tl_h_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)], tl_h_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)], tl_h_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)], tl_h_i[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)], tl_h_i[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))], tl_h_i[53-:32], tl_h_i[21-:21], spare_req_i}),
		.rvalid_o(tl_d_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))]),
		.rready_i(tl_d_i[0]),
		.rdata_o({reqfifo_tl_d_a_opcode, tl_d_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)], tl_d_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)], tl_d_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)], tl_d_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)], tl_d_o[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))], tl_d_o[53-:32], tl_d_o[21-:21], spare_req_o}),
		.full_o(),
		.depth_o()
	);
	// Trace: design.sv:74476:3
	localparam [31:0] RSPFIFO_WIDTH = ((1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 2) + SpareRspW;
	// Trace: design.sv:74477:3
	wire [2:0] rspfifo_tl_h_d_opcode;
	// Trace: design.sv:74479:3
	assign tl_h_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = rspfifo_tl_h_d_opcode;
	// Trace: design.sv:74481:3
	prim_fifo_sync #(
		.Width(RSPFIFO_WIDTH),
		.Pass(RspPass),
		.Depth(RspDepth)
	) rspfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(tl_d_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))]),
		.wready_o(tl_d_o[0]),
		.wdata_i({tl_d_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_d_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_d_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_d_i[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_d_i[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], (tl_d_i[6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) - (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))))) + 1 : ((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) - (6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))))) + 1)] == 3'h1 ? tl_d_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)] : {top_pkg_TL_DW {1'b0}}), tl_d_i[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))], tl_d_i[1], spare_rsp_i}),
		.rvalid_o(tl_h_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))]),
		.rready_i(tl_h_i[0]),
		.rdata_o({rspfifo_tl_h_d_opcode, tl_h_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_h_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_h_o[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_h_o[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], tl_h_o[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)], tl_h_o[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))], tl_h_o[1], spare_rsp_o}),
		.full_o(),
		.depth_o()
	);
endmodule
module tlul_fifo_async (
	clk_h_i,
	rst_h_ni,
	clk_d_i,
	rst_d_ni,
	tl_h_i,
	tl_h_o,
	tl_d_o,
	tl_d_i
);
	// Trace: design.sv:74523:13
	parameter [31:0] ReqDepth = 3;
	// Trace: design.sv:74524:13
	parameter [31:0] RspDepth = 3;
	// Trace: design.sv:74526:3
	input clk_h_i;
	// Trace: design.sv:74527:3
	input rst_h_ni;
	// Trace: design.sv:74528:3
	input clk_d_i;
	// Trace: design.sv:74529:3
	input rst_d_ni;
	// Trace: design.sv:74530:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_h_i;
	// Trace: design.sv:74531:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o;
	// Trace: design.sv:74532:3
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_d_o;
	// Trace: design.sv:74533:3
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d_i;
	// Trace: design.sv:74537:3
	localparam [31:0] REQFIFO_WIDTH = (1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)) - 2;
	// Trace: design.sv:74538:3
	wire [2:0] reqfifo_tl_d_a_opcode;
	// Trace: design.sv:74540:3
	assign tl_d_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] = reqfifo_tl_d_a_opcode;
	// Trace: design.sv:74542:3
	prim_fifo_async #(
		.Width(REQFIFO_WIDTH),
		.Depth(ReqDepth)
	) reqfifo(
		.clk_wr_i(clk_h_i),
		.rst_wr_ni(rst_h_ni),
		.clk_rd_i(clk_d_i),
		.rst_rd_ni(rst_d_ni),
		.wvalid_i(tl_h_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))]),
		.wready_o(tl_h_o[0]),
		.wdata_i({tl_h_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)], tl_h_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)], tl_h_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)], tl_h_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)], tl_h_i[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)], tl_h_i[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))], tl_h_i[53-:32], tl_h_i[21-:21]}),
		.rvalid_o(tl_d_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))]),
		.rready_i(tl_d_i[0]),
		.rdata_o({reqfifo_tl_d_a_opcode, tl_d_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)], tl_d_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)], tl_d_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)], tl_d_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)], tl_d_o[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))], tl_d_o[53-:32], tl_d_o[21-:21]}),
		.wdepth_o(),
		.rdepth_o()
	);
	// Trace: design.sv:74573:3
	localparam [31:0] RSPFIFO_WIDTH = (1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 2;
	// Trace: design.sv:74574:3
	wire [2:0] rspfifo_tl_h_d_opcode;
	// Trace: design.sv:74576:3
	assign tl_h_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = rspfifo_tl_h_d_opcode;
	// Trace: design.sv:74578:3
	prim_fifo_async #(
		.Width(RSPFIFO_WIDTH),
		.Depth(RspDepth)
	) rspfifo(
		.clk_wr_i(clk_d_i),
		.rst_wr_ni(rst_d_ni),
		.clk_rd_i(clk_h_i),
		.rst_rd_ni(rst_h_ni),
		.wvalid_i(tl_d_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))]),
		.wready_o(tl_d_o[0]),
		.wdata_i({tl_d_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_d_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_d_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_d_i[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_d_i[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], tl_d_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)], tl_d_i[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))], tl_d_i[1]}),
		.rvalid_o(tl_h_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))]),
		.rready_i(tl_h_i[0]),
		.rdata_o({rspfifo_tl_h_d_opcode, tl_h_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_h_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_h_o[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_h_o[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], tl_h_o[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)], tl_h_o[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))], tl_h_o[1]}),
		.wdepth_o(),
		.rdepth_o()
	);
endmodule
module tlul_assert (
	clk_i,
	rst_ni,
	h2d,
	d2h
);
	// Trace: design.sv:74623:13
	parameter EndpointType = "Device";
	// Trace: design.sv:74625:3
	input clk_i;
	// Trace: design.sv:74626:3
	input rst_ni;
	// Trace: design.sv:74629:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] h2d;
	// Trace: design.sv:74630:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] d2h;
endmodule
module tlul_err (
	clk_i,
	rst_ni,
	tl_i,
	err_o
);
	reg _sv2v_0;
	// removed import tlul_pkg::*;
	// Trace: design.sv:75004:3
	input clk_i;
	// Trace: design.sv:75005:3
	input rst_ni;
	// Trace: design.sv:75007:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:75009:3
	output wire err_o;
	// Trace: design.sv:75012:3
	localparam signed [31:0] IW = top_pkg_TL_AIW;
	// Trace: design.sv:75013:3
	localparam signed [31:0] SZW = top_pkg_TL_SZW;
	// Trace: design.sv:75014:3
	localparam signed [31:0] DW = top_pkg_TL_DW;
	// Trace: design.sv:75015:3
	localparam signed [31:0] MW = top_pkg_TL_DBW;
	// Trace: design.sv:75016:3
	localparam signed [31:0] SubAW = 2;
	// Trace: design.sv:75018:3
	wire opcode_allowed;
	wire a_config_allowed;
	// Trace: design.sv:75020:3
	wire op_full;
	wire op_partial;
	wire op_get;
	// Trace: design.sv:75021:3
	assign op_full = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h0;
	// Trace: design.sv:75022:3
	assign op_partial = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h1;
	// Trace: design.sv:75023:3
	assign op_get = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h4;
	// Trace: design.sv:75026:3
	wire instr_wr_err;
	// Trace: design.sv:75027:3
	assign instr_wr_err = (tl_i[16-:2] == 2'b01) & (op_full | op_partial);
	// Trace: design.sv:75031:3
	assign err_o = ~(opcode_allowed & a_config_allowed) | instr_wr_err;
	// Trace: design.sv:75034:3
	assign opcode_allowed = ((tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h0) | (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h1)) | (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h4);
	// Trace: design.sv:75039:3
	reg addr_sz_chk;
	// Trace: design.sv:75040:3
	reg mask_chk;
	// Trace: design.sv:75041:3
	reg fulldata_chk;
	// Trace: design.sv:75043:3
	wire [MW - 1:0] mask;
	// Trace: design.sv:75045:3
	assign mask = 1 << tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 30:(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 31];
	// Trace: design.sv:75047:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:75048:5
		addr_sz_chk = 1'b0;
		// Trace: design.sv:75049:5
		mask_chk = 1'b0;
		// Trace: design.sv:75050:5
		fulldata_chk = 1'b0;
		// Trace: design.sv:75052:5
		if (tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))])
			// Trace: design.sv:75053:7
			(* full_case, parallel_case *)
			case (tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)])
				'h0: begin
					// Trace: design.sv:75055:11
					addr_sz_chk = 1'b1;
					// Trace: design.sv:75056:11
					mask_chk = ~|(tl_i[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))] & ~mask);
					// Trace: design.sv:75057:11
					fulldata_chk = |(tl_i[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))] & mask);
				end
				'h1: begin
					// Trace: design.sv:75061:11
					addr_sz_chk = ~tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 31];
					// Trace: design.sv:75063:11
					mask_chk = (tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 30] ? ~|(tl_i[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))] & 4'b0011) : ~|(tl_i[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))] & 4'b1100));
					// Trace: design.sv:75065:11
					fulldata_chk = (tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 30] ? &tl_i[(top_pkg_TL_DBW + 53) - (top_pkg_TL_DBW - 4):(top_pkg_TL_DBW + 53) - (top_pkg_TL_DBW - 3)] : &tl_i[(top_pkg_TL_DBW + 53) - (top_pkg_TL_DBW - 2):(top_pkg_TL_DBW + 53) - (top_pkg_TL_DBW - 1)]);
				end
				'h2: begin
					// Trace: design.sv:75069:11
					addr_sz_chk = ~|tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 30:(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 31];
					// Trace: design.sv:75070:11
					mask_chk = 1'b1;
					// Trace: design.sv:75071:11
					fulldata_chk = &tl_i[(top_pkg_TL_DBW + 53) - (top_pkg_TL_DBW - 4):(top_pkg_TL_DBW + 53) - (top_pkg_TL_DBW - 1)];
				end
				default: begin
					// Trace: design.sv:75075:11
					addr_sz_chk = 1'b0;
					// Trace: design.sv:75076:11
					mask_chk = 1'b0;
					// Trace: design.sv:75077:11
					fulldata_chk = 1'b0;
				end
			endcase
		else begin
			// Trace: design.sv:75081:7
			addr_sz_chk = 1'b0;
			// Trace: design.sv:75082:7
			mask_chk = 1'b0;
			// Trace: design.sv:75083:7
			fulldata_chk = 1'b0;
		end
	end
	// Trace: design.sv:75087:3
	assign a_config_allowed = (addr_sz_chk & mask_chk) & ((op_get | op_partial) | fulldata_chk);
	initial _sv2v_0 = 0;
endmodule
module tlul_assert_multiple (
	clk_i,
	rst_ni,
	h2d,
	d2h
);
	// Trace: design.sv:75102:13
	parameter [31:0] N = 2;
	// Trace: design.sv:75103:13
	parameter EndpointType = "Device";
	// Trace: design.sv:75105:3
	input clk_i;
	// Trace: design.sv:75106:3
	input rst_ni;
	// Trace: design.sv:75109:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? (N * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)) - 1 : (N * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 20)):(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21)] h2d;
	// Trace: design.sv:75110:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	input wire [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (N * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 1 : (N * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 0)):((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)] d2h;
	// Trace: design.sv:75114:3
	genvar _gv_ii_1;
	generate
		for (_gv_ii_1 = 0; _gv_ii_1 < N; _gv_ii_1 = _gv_ii_1 + 1) begin : gen_assert
			localparam ii = _gv_ii_1;
			// Trace: design.sv:75115:5
			tlul_assert #(.EndpointType(EndpointType)) tlul_assert(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.h2d(h2d[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21) + (((N - 1) - ii) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21)))+:(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21))]),
				.d2h(d2h[((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1) + (((N - 1) - ii) * ((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)))+:((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))])
			);
		end
	endgenerate
endmodule
// removed package "spi_host_reg_pkg"
// removed package "spi_host_cmd_pkg"
module spi_host_shift_register (
	clk_i,
	rst_ni,
	wr_en_i,
	wr_ready_o,
	rd_en_i,
	rd_ready_o,
	speed_i,
	shift_en_i,
	sample_en_i,
	full_cyc_i,
	last_read_i,
	last_write_i,
	tx_data_i,
	tx_valid_i,
	tx_ready_o,
	tx_flush_o,
	rx_data_o,
	rx_valid_o,
	rx_ready_i,
	rx_last_o,
	sd_i,
	sd_o,
	sw_rst_i
);
	// Trace: design.sv:75559:3
	input clk_i;
	// Trace: design.sv:75560:3
	input rst_ni;
	// Trace: design.sv:75561:3
	input wr_en_i;
	// Trace: design.sv:75562:3
	output wire wr_ready_o;
	// Trace: design.sv:75563:3
	input rd_en_i;
	// Trace: design.sv:75564:3
	output wire rd_ready_o;
	// Trace: design.sv:75566:3
	input [1:0] speed_i;
	// Trace: design.sv:75567:3
	input shift_en_i;
	// Trace: design.sv:75568:3
	input sample_en_i;
	// Trace: design.sv:75569:3
	input full_cyc_i;
	// Trace: design.sv:75570:3
	input last_read_i;
	// Trace: design.sv:75571:3
	input last_write_i;
	// Trace: design.sv:75573:3
	input [7:0] tx_data_i;
	// Trace: design.sv:75574:3
	input tx_valid_i;
	// Trace: design.sv:75575:3
	output wire tx_ready_o;
	// Trace: design.sv:75576:3
	output wire tx_flush_o;
	// Trace: design.sv:75578:3
	output wire [7:0] rx_data_o;
	// Trace: design.sv:75579:3
	output wire rx_valid_o;
	// Trace: design.sv:75580:3
	input rx_ready_i;
	// Trace: design.sv:75581:3
	output wire rx_last_o;
	// Trace: design.sv:75583:3
	input [3:0] sd_i;
	// Trace: design.sv:75584:3
	output wire [3:0] sd_o;
	// Trace: design.sv:75586:3
	input sw_rst_i;
	// Trace: design.sv:75588:3
	// removed import spi_host_cmd_pkg::*;
	// Trace: design.sv:75590:3
	reg [7:0] sr_q;
	// Trace: design.sv:75591:3
	wire [7:0] sr_d;
	// Trace: design.sv:75592:3
	reg [3:0] sd_i_q;
	wire [3:0] sd_i_d;
	// Trace: design.sv:75593:3
	wire [3:0] next_bits;
	// Trace: design.sv:75594:3
	wire [7:0] sr_shifted;
	// Trace: design.sv:75599:3
	reg [8:0] rx_buf_q;
	// Trace: design.sv:75600:3
	wire [8:0] rx_buf_d;
	// Trace: design.sv:75601:3
	reg rx_buf_valid_q;
	// Trace: design.sv:75602:3
	wire rx_buf_valid_d;
	// Trace: design.sv:75606:3
	assign next_bits = (full_cyc_i ? sd_i : sd_i_q);
	// Trace: design.sv:75607:3
	// removed localparam type spi_host_cmd_pkg_speed_t
	assign sr_shifted = (speed_i == 2'b00 ? {sr_q[6:0], next_bits[1]} : (speed_i == 2'b01 ? {sr_q[5:0], next_bits[1:0]} : (speed_i == 2'b10 ? {sr_q[3:0], next_bits[3:0]} : 8'h00)));
	// Trace: design.sv:75612:3
	assign sd_o = (speed_i == 2'b00 ? {3'b000, sr_q[7]} : (speed_i == 2'b01 ? {2'b00, sr_q[7:6]} : (speed_i == 2'b10 ? {sr_q[7:4]} : 4'h0)));
	// Trace: design.sv:75619:3
	assign rd_ready_o = ~rx_buf_valid_q | (rx_valid_o & rx_ready_i);
	// Trace: design.sv:75620:3
	assign rx_valid_o = rx_buf_valid_q;
	// Trace: design.sv:75622:3
	assign rx_buf_d = (sw_rst_i ? 9'h000 : (rd_en_i && rd_ready_o ? {last_read_i, sr_shifted} : rx_buf_q));
	// Trace: design.sv:75626:3
	assign rx_buf_valid_d = (sw_rst_i ? 1'b0 : (rd_en_i && rd_ready_o ? 1'b1 : (rx_valid_o & rx_ready_i ? 1'b0 : rx_buf_valid_q)));
	// Trace: design.sv:75631:3
	assign sd_i_d = (sw_rst_i ? 4'b0000 : (sample_en_i ? sd_i : sd_i_q));
	// Trace: design.sv:75635:3
	assign {rx_last_o, rx_data_o} = rx_buf_q;
	// Trace: design.sv:75640:3
	assign wr_ready_o = tx_valid_i;
	// Trace: design.sv:75641:3
	assign tx_ready_o = wr_en_i;
	// Trace: design.sv:75642:3
	assign tx_flush_o = last_write_i;
	// Trace: design.sv:75644:3
	assign sr_d = (sw_rst_i ? 8'h00 : (wr_en_i & wr_ready_o ? tx_data_i : (shift_en_i ? sr_shifted : sr_q)));
	// Trace: design.sv:75649:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:75650:5
		if (!rst_ni) begin
			// Trace: design.sv:75651:7
			sd_i_q <= 4'h0;
			// Trace: design.sv:75652:7
			sr_q <= 8'h00;
			// Trace: design.sv:75653:7
			rx_buf_valid_q <= 1'b0;
			// Trace: design.sv:75654:7
			rx_buf_q <= 9'h000;
		end
		else begin
			// Trace: design.sv:75656:7
			sd_i_q <= sd_i_d;
			// Trace: design.sv:75657:7
			sr_q <= sr_d;
			// Trace: design.sv:75658:7
			rx_buf_valid_q <= rx_buf_valid_d;
			// Trace: design.sv:75659:7
			rx_buf_q <= rx_buf_d;
		end
endmodule
module spi_host_byte_select (
	clk_i,
	rst_ni,
	word_i,
	word_be_i,
	word_valid_i,
	word_ready_o,
	byte_o,
	byte_valid_o,
	byte_ready_i,
	flush_i,
	sw_rst_i
);
	// Trace: design.sv:75671:3
	input clk_i;
	// Trace: design.sv:75672:3
	input rst_ni;
	// Trace: design.sv:75673:3
	input [31:0] word_i;
	// Trace: design.sv:75674:3
	input [3:0] word_be_i;
	// Trace: design.sv:75675:3
	input word_valid_i;
	// Trace: design.sv:75676:3
	output wire word_ready_o;
	// Trace: design.sv:75677:3
	output wire [7:0] byte_o;
	// Trace: design.sv:75678:3
	output wire byte_valid_o;
	// Trace: design.sv:75679:3
	input byte_ready_i;
	// Trace: design.sv:75680:3
	input flush_i;
	// Trace: design.sv:75681:3
	input sw_rst_i;
	// Trace: design.sv:75684:3
	wire [35:0] wdata_be;
	// Trace: design.sv:75685:3
	wire do_drain;
	// Trace: design.sv:75686:3
	wire byte_en;
	// Trace: design.sv:75687:3
	wire byte_valid;
	// Trace: design.sv:75688:3
	wire byte_ready;
	// Trace: design.sv:75689:3
	wire clr;
	// Trace: design.sv:75691:3
	assign clr = flush_i | sw_rst_i;
	// Trace: design.sv:75692:3
	assign byte_valid_o = byte_valid & byte_en;
	// Trace: design.sv:75693:3
	assign do_drain = byte_valid & ~byte_en;
	// Trace: design.sv:75694:3
	assign byte_ready = byte_ready_i | do_drain;
	// Trace: design.sv:75696:3
	genvar _gv_ii_2;
	generate
		for (_gv_ii_2 = 0; _gv_ii_2 < 4; _gv_ii_2 = _gv_ii_2 + 1) begin : gen_map_data_be
			localparam ii = _gv_ii_2;
			// Trace: design.sv:75697:5
			assign wdata_be[9 * ii+:9] = {word_be_i[ii], word_i[8 * ii+:8]};
		end
	endgenerate
	// Trace: design.sv:75700:3
	prim_packer_fifo #(
		.InW(36),
		.OutW(9)
	) u_packer(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(clr),
		.wdata_i(wdata_be),
		.wvalid_i(word_valid_i),
		.wready_o(word_ready_o),
		.rdata_o({byte_en, byte_o}),
		.rvalid_o(byte_valid),
		.rready_i(byte_ready),
		.depth_o()
	);
endmodule
module spi_host_byte_merge (
	clk_i,
	rst_ni,
	byte_i,
	byte_last_i,
	byte_valid_i,
	byte_ready_o,
	word_o,
	word_valid_o,
	word_ready_i,
	sw_rst_i
);
	// Trace: design.sv:75725:3
	input clk_i;
	// Trace: design.sv:75726:3
	input rst_ni;
	// Trace: design.sv:75727:3
	input [7:0] byte_i;
	// Trace: design.sv:75728:3
	input byte_last_i;
	// Trace: design.sv:75729:3
	input byte_valid_i;
	// Trace: design.sv:75730:3
	output wire byte_ready_o;
	// Trace: design.sv:75731:3
	output wire [31:0] word_o;
	// Trace: design.sv:75732:3
	output wire word_valid_o;
	// Trace: design.sv:75733:3
	input word_ready_i;
	// Trace: design.sv:75734:3
	input sw_rst_i;
	// Trace: design.sv:75737:3
	wire clr;
	// Trace: design.sv:75738:3
	wire byte_valid;
	// Trace: design.sv:75739:3
	wire byte_ready;
	// Trace: design.sv:75740:3
	reg last_q;
	// Trace: design.sv:75741:3
	wire last_d;
	// Trace: design.sv:75742:3
	wire do_fill;
	// Trace: design.sv:75743:3
	wire byte_incoming;
	// Trace: design.sv:75746:3
	assign clr = sw_rst_i;
	// Trace: design.sv:75747:3
	assign byte_incoming = byte_valid_i & byte_ready_o;
	// Trace: design.sv:75749:3
	assign last_d = (sw_rst_i ? 1'b0 : (byte_incoming && byte_last_i ? 1'b1 : (word_valid_o ? 1'b0 : last_q)));
	// Trace: design.sv:75754:3
	assign do_fill = last_q & ~word_valid_o;
	// Trace: design.sv:75755:3
	assign byte_valid = do_fill | byte_valid_i;
	// Trace: design.sv:75756:3
	assign byte_ready_o = byte_ready & ~do_fill;
	// Trace: design.sv:75758:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:75759:5
		if (!rst_ni)
			// Trace: design.sv:75760:7
			last_q <= 1'b0;
		else
			// Trace: design.sv:75762:7
			last_q <= last_d;
	// Trace: design.sv:75766:3
	prim_packer_fifo #(
		.InW(8),
		.OutW(32)
	) u_packer(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(clr),
		.wdata_i((do_fill ? 8'h00 : byte_i)),
		.wvalid_i(byte_valid),
		.wready_o(byte_ready),
		.rdata_o(word_o),
		.rvalid_o(word_valid_o),
		.rready_i(word_ready_i),
		.depth_o()
	);
endmodule
module spi_host_fsm (
	clk_i,
	rst_ni,
	en_i,
	command_i,
	command_valid_i,
	command_ready_o,
	sck_o,
	csb_o,
	sd_en_o,
	last_read_o,
	last_write_o,
	wr_en_o,
	sr_wr_ready_i,
	rd_en_o,
	sr_rd_ready_i,
	sample_en_o,
	shift_en_o,
	speed_o,
	full_cyc_o,
	rx_stall_o,
	tx_stall_o,
	active_o,
	sw_rst_i
);
	reg _sv2v_0;
	// removed import spi_host_cmd_pkg::*;
	// Trace: design.sv:75795:14
	parameter signed [31:0] NumCS = 1;
	// Trace: design.sv:75797:3
	input clk_i;
	// Trace: design.sv:75798:3
	input rst_ni;
	// Trace: design.sv:75799:3
	input en_i;
	// Trace: design.sv:75800:3
	function automatic integer prim_util_pkg_vbits;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:74:36
		input integer value;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:85:5
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] spi_host_reg_pkg_NumCS = 2;
	localparam signed [31:0] spi_host_cmd_pkg_CSW = prim_util_pkg_vbits(spi_host_reg_pkg_NumCS);
	// removed localparam type spi_host_cmd_pkg_configopts_t
	// removed localparam type spi_host_cmd_pkg_segment_t
	// removed localparam type spi_host_cmd_pkg_command_t
	input wire [spi_host_cmd_pkg_CSW + 59:0] command_i;
	// Trace: design.sv:75801:3
	input command_valid_i;
	// Trace: design.sv:75802:3
	output wire command_ready_o;
	// Trace: design.sv:75803:3
	output wire sck_o;
	// Trace: design.sv:75804:3
	output wire [NumCS - 1:0] csb_o;
	// Trace: design.sv:75805:3
	output reg [3:0] sd_en_o;
	// Trace: design.sv:75806:3
	output wire last_read_o;
	// Trace: design.sv:75807:3
	output wire last_write_o;
	// Trace: design.sv:75808:3
	output wire wr_en_o;
	// Trace: design.sv:75809:3
	input sr_wr_ready_i;
	// Trace: design.sv:75810:3
	output wire rd_en_o;
	// Trace: design.sv:75811:3
	input sr_rd_ready_i;
	// Trace: design.sv:75812:3
	output wire sample_en_o;
	// Trace: design.sv:75813:3
	output wire shift_en_o;
	// Trace: design.sv:75814:3
	output wire [1:0] speed_o;
	// Trace: design.sv:75815:3
	output wire full_cyc_o;
	// Trace: design.sv:75816:3
	output wire rx_stall_o;
	// Trace: design.sv:75817:3
	output wire tx_stall_o;
	// Trace: design.sv:75818:3
	output wire active_o;
	// Trace: design.sv:75820:3
	input sw_rst_i;
	// Trace: design.sv:75823:3
	wire is_idle;
	// Trace: design.sv:75824:3
	reg [15:0] clkdiv;
	reg [15:0] clkdiv_q;
	// Trace: design.sv:75825:3
	reg [15:0] clk_cntr_q;
	wire [15:0] clk_cntr_d;
	// Trace: design.sv:75826:3
	wire clk_cntr_en;
	// Trace: design.sv:75828:3
	wire [1:0] speed_cpha0;
	reg [1:0] speed_cpha1;
	// Trace: design.sv:75830:3
	reg [spi_host_cmd_pkg_CSW - 1:0] csid;
	// Trace: design.sv:75831:3
	reg [spi_host_cmd_pkg_CSW - 1:0] csid_q;
	// Trace: design.sv:75833:3
	reg [3:0] csnidle;
	reg [3:0] csntrail;
	reg [3:0] csnlead;
	// Trace: design.sv:75834:3
	reg [3:0] csnidle_q;
	reg [3:0] csntrail_q;
	reg [3:0] csnlead_q;
	// Trace: design.sv:75835:3
	reg full_cyc;
	reg cpha;
	reg cpol;
	// Trace: design.sv:75836:3
	reg full_cyc_q;
	reg cpha_q;
	reg cpol_q;
	// Trace: design.sv:75848:3
	reg [1:0] cmd_speed_d;
	reg [1:0] cmd_speed_q;
	// Trace: design.sv:75849:3
	reg cmd_wr_en_d;
	reg cmd_wr_en_q;
	// Trace: design.sv:75850:3
	reg cmd_rd_en_d;
	reg cmd_rd_en_q;
	// Trace: design.sv:75851:3
	reg [23:0] cmd_len_d;
	reg [23:0] cmd_len_q;
	// Trace: design.sv:75852:3
	reg csaat;
	// Trace: design.sv:75853:3
	reg csaat_q;
	// Trace: design.sv:75855:3
	wire [2:0] bit_cntr_d;
	reg [2:0] bit_cntr_q;
	// Trace: design.sv:75856:3
	wire [23:0] byte_cntr_cpha0_d;
	wire [23:0] byte_cntr_cpha1_d;
	reg [23:0] byte_cntr_cpha0_q;
	reg [23:0] byte_cntr_cpha1_q;
	// Trace: design.sv:75857:3
	wire [23:0] byte_cntr_early;
	wire [23:0] byte_cntr_late;
	// Trace: design.sv:75858:3
	reg [3:0] wait_cntr_d;
	reg [3:0] wait_cntr_q;
	// Trace: design.sv:75859:3
	wire last_bit;
	wire last_byte;
	// Trace: design.sv:75861:3
	wire state_changing;
	// Trace: design.sv:75862:3
	wire byte_starting;
	wire byte_starting_cpha0;
	reg byte_starting_cpha0_q;
	wire byte_starting_cpha1;
	// Trace: design.sv:75863:3
	wire bit_shifting;
	wire bit_shifting_cpha0;
	reg bit_shifting_cpha0_q;
	wire bit_shifting_cpha1;
	// Trace: design.sv:75864:3
	wire byte_ending;
	wire byte_ending_cpha0;
	reg byte_ending_cpha0_q;
	wire byte_ending_cpha1;
	// Trace: design.sv:75866:3
	wire sample_en_d;
	reg sample_en_q;
	reg sample_en_q2;
	// Trace: design.sv:75868:3
	wire config_changed;
	// Trace: design.sv:75869:3
	wire fsm_en;
	// Trace: design.sv:75874:3
	wire new_command;
	reg new_command_cpha1;
	// Trace: design.sv:75876:3
	reg csb_single_d;
	// Trace: design.sv:75877:3
	reg [NumCS - 1:0] csb_q;
	// Trace: design.sv:75878:3
	wire sck_d;
	wire sck_q;
	// Trace: design.sv:75880:3
	wire wr_en_internal;
	wire rd_en_internal;
	wire sample_en_internal;
	wire shift_en_internal;
	// Trace: design.sv:75882:3
	wire stall;
	// Trace: design.sv:75884:3
	assign stall = rx_stall_o | tx_stall_o;
	// Trace: design.sv:75887:3
	assign wr_en_o = wr_en_internal & ~stall;
	// Trace: design.sv:75888:3
	assign rd_en_o = rd_en_internal & ~stall;
	// Trace: design.sv:75889:3
	assign sample_en_o = sample_en_internal & ~stall;
	// Trace: design.sv:75890:3
	assign shift_en_o = shift_en_internal & ~stall;
	// Trace: design.sv:75892:3
	// removed localparam type spi_host_st_e
	// Trace: design.sv:75903:3
	reg [2:0] state_q;
	reg [2:0] state_d;
	// Trace: design.sv:75905:3
	reg command_ready_int;
	// Trace: design.sv:75906:3
	assign command_ready_o = command_ready_int & ~stall;
	// Trace: design.sv:75909:3
	assign new_command = command_valid_i && command_ready_int;
	// Trace: design.sv:75910:3
	assign config_changed = ((((((command_i[0] != cpol_q) || (command_i[1] != cpha_q)) || (command_i[2] != full_cyc_q)) || (command_i[14-:4] != csnidle_q)) || (command_i[6-:4] != csntrail_q)) || (command_i[10-:4] != csnlead_q)) || (command_i[30-:16] != clkdiv_q);
	// Trace: design.sv:75918:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:75919:5
		csid = (new_command ? command_i[spi_host_cmd_pkg_CSW + 59-:((spi_host_cmd_pkg_CSW + 59) >= 60 ? spi_host_cmd_pkg_CSW + 0 : 61 - (spi_host_cmd_pkg_CSW + 59))] : csid_q);
		// Trace: design.sv:75920:5
		cpol = (new_command ? command_i[0] : cpol_q);
		// Trace: design.sv:75921:5
		cpha = (new_command ? command_i[1] : cpha_q);
		// Trace: design.sv:75922:5
		full_cyc = (new_command ? command_i[2] : full_cyc_q);
		// Trace: design.sv:75923:5
		csnidle = (new_command ? command_i[14-:4] : csnidle_q);
		// Trace: design.sv:75924:5
		csnlead = (new_command ? command_i[10-:4] : csnlead_q);
		// Trace: design.sv:75925:5
		csntrail = (new_command ? command_i[6-:4] : csntrail_q);
		// Trace: design.sv:75926:5
		clkdiv = (new_command ? command_i[30-:16] : clkdiv_q);
		// Trace: design.sv:75927:5
		csaat = (new_command ? command_i[31] : csaat_q);
		// Trace: design.sv:75928:5
		cmd_len_d = (new_command ? command_i[55-:24] : cmd_len_q);
		// Trace: design.sv:75929:5
		cmd_wr_en_d = (new_command ? command_i[57] : cmd_wr_en_q);
		// Trace: design.sv:75930:5
		cmd_rd_en_d = (new_command ? command_i[56] : cmd_rd_en_q);
		// Trace: design.sv:75931:5
		cmd_speed_d = (new_command ? command_i[59-:2] : cmd_speed_q);
	end
	// Trace: design.sv:75934:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:75935:5
		if (!rst_ni) begin
			// Trace: design.sv:75936:7
			csid_q <= {spi_host_cmd_pkg_CSW {1'b0}};
			// Trace: design.sv:75937:7
			cpol_q <= 1'b0;
			// Trace: design.sv:75938:7
			cpha_q <= 1'b0;
			// Trace: design.sv:75939:7
			full_cyc_q <= 1'b0;
			// Trace: design.sv:75940:7
			csnidle_q <= 4'h0;
			// Trace: design.sv:75941:7
			csnlead_q <= 4'h0;
			// Trace: design.sv:75942:7
			csntrail_q <= 4'h0;
			// Trace: design.sv:75943:7
			clkdiv_q <= 16'h0000;
			// Trace: design.sv:75944:7
			csaat_q <= 1'b0;
			// Trace: design.sv:75945:7
			cmd_rd_en_q <= 1'b0;
			// Trace: design.sv:75946:7
			cmd_wr_en_q <= 1'b0;
			// Trace: design.sv:75947:7
			cmd_speed_q <= 2'b00;
			// Trace: design.sv:75948:7
			cmd_len_q <= 24'h000000;
		end
		else begin
			// Trace: design.sv:75950:7
			csid_q <= (new_command && !stall ? csid : csid_q);
			// Trace: design.sv:75951:7
			cpol_q <= (new_command && !stall ? cpol : cpol_q);
			// Trace: design.sv:75952:7
			cpha_q <= (new_command && !stall ? cpha : cpha_q);
			// Trace: design.sv:75953:7
			full_cyc_q <= (new_command && !stall ? full_cyc : full_cyc_q);
			// Trace: design.sv:75954:7
			csnidle_q <= (new_command && !stall ? csnidle : csnidle_q);
			// Trace: design.sv:75955:7
			csnlead_q <= (new_command && !stall ? csnlead : csnlead_q);
			// Trace: design.sv:75956:7
			csntrail_q <= (new_command && !stall ? csntrail : csntrail_q);
			// Trace: design.sv:75957:7
			clkdiv_q <= (new_command && !stall ? clkdiv : clkdiv_q);
			// Trace: design.sv:75958:7
			csaat_q <= (new_command && !stall ? csaat : csaat_q);
			// Trace: design.sv:75959:7
			cmd_wr_en_q <= (new_command && !stall ? cmd_wr_en_d : cmd_wr_en_q);
			// Trace: design.sv:75960:7
			cmd_rd_en_q <= (new_command && !stall ? cmd_rd_en_d : cmd_rd_en_q);
			// Trace: design.sv:75961:7
			cmd_speed_q <= (new_command && !stall ? cmd_speed_d : cmd_speed_q);
			// Trace: design.sv:75962:7
			cmd_len_q <= (new_command && !stall ? cmd_len_d : cmd_len_q);
		end
	// Trace: design.sv:75966:3
	assign is_idle = (state_q == 3'd0) || (state_q == 3'd7);
	// Trace: design.sv:75968:3
	assign active_o = ~is_idle;
	// Trace: design.sv:75970:3
	assign clk_cntr_d = (sw_rst_i ? 16'h0000 : (!clk_cntr_en ? clk_cntr_q : (is_idle ? 16'h0000 : (new_command ? clkdiv : (clk_cntr_q == 16'h0000 ? clkdiv : clk_cntr_q - 1)))));
	// Trace: design.sv:75977:3
	assign tx_stall_o = wr_en_internal & ~sr_wr_ready_i;
	// Trace: design.sv:75978:3
	assign rx_stall_o = rd_en_internal & ~sr_rd_ready_i;
	// Trace: design.sv:75979:3
	assign clk_cntr_en = en_i;
	// Trace: design.sv:75980:3
	assign fsm_en = clk_cntr_en && (clk_cntr_q == 0);
	// Trace: design.sv:75982:3
	reg [2:0] next_state_after_idle;
	// Trace: design.sv:75983:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:75984:5
		if (command_valid_i) begin
			begin
				// Trace: design.sv:75985:7
				if (config_changed)
					// Trace: design.sv:75986:10
					next_state_after_idle = 3'd6;
				else
					// Trace: design.sv:75988:10
					next_state_after_idle = 3'd1;
			end
		end
		else
			// Trace: design.sv:75991:7
			next_state_after_idle = 3'd0;
	end
	// Trace: design.sv:75995:3
	reg [2:0] next_state_after_idle_csb_active;
	// Trace: design.sv:75996:3
	reg command_ready_idle_csb_active;
	// Trace: design.sv:75997:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:75998:5
		if (command_valid_i) begin
			begin
				// Trace: design.sv:75999:7
				if (command_i[spi_host_cmd_pkg_CSW + 59-:((spi_host_cmd_pkg_CSW + 59) >= 60 ? spi_host_cmd_pkg_CSW + 0 : 61 - (spi_host_cmd_pkg_CSW + 59))] != csid_q) begin
					// Trace: design.sv:76006:9
					next_state_after_idle_csb_active = 3'd4;
					// Trace: design.sv:76008:9
					command_ready_idle_csb_active = 1'b0;
				end
				else begin
					// Trace: design.sv:76010:9
					next_state_after_idle_csb_active = 3'd2;
					// Trace: design.sv:76011:9
					command_ready_idle_csb_active = 1'b1;
				end
			end
		end
		else begin
			// Trace: design.sv:76014:7
			next_state_after_idle_csb_active = 3'd7;
			// Trace: design.sv:76015:7
			command_ready_idle_csb_active = 1'b1;
		end
	end
	// Trace: design.sv:76022:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:76023:5
		state_d = state_q;
		// Trace: design.sv:76024:5
		command_ready_int = 1'b0;
		// Trace: design.sv:76025:5
		if (sw_rst_i)
			// Trace: design.sv:76026:7
			state_d = 3'd0;
		else if (fsm_en)
			// Trace: design.sv:76028:7
			(* full_case, parallel_case *)
			case (state_q)
				3'd0: begin
					// Trace: design.sv:76031:11
					command_ready_int = 1'b1;
					// Trace: design.sv:76032:11
					state_d = next_state_after_idle;
				end
				3'd1:
					// Trace: design.sv:76036:11
					if (wait_cntr_q == 4'h0)
						// Trace: design.sv:76037:13
						state_d = 3'd3;
				3'd2:
					// Trace: design.sv:76042:11
					state_d = 3'd3;
				3'd3:
					// Trace: design.sv:76048:11
					if (!last_bit || !last_byte)
						// Trace: design.sv:76049:13
						state_d = 3'd2;
					else if (!csaat_q)
						// Trace: design.sv:76052:13
						state_d = 3'd4;
					else begin
						// Trace: design.sv:76054:13
						state_d = next_state_after_idle_csb_active;
						// Trace: design.sv:76055:13
						command_ready_int = command_ready_idle_csb_active;
					end
				3'd4:
					// Trace: design.sv:76060:11
					if (wait_cntr_q == 4'h0)
						// Trace: design.sv:76061:13
						state_d = 3'd5;
				3'd5:
					// Trace: design.sv:76066:11
					if (wait_cntr_q == 4'h0) begin
						// Trace: design.sv:76068:13
						command_ready_int = 1'b1;
						// Trace: design.sv:76069:13
						state_d = next_state_after_idle;
					end
				3'd6:
					// Trace: design.sv:76076:11
					if (wait_cntr_q == 4'h0)
						// Trace: design.sv:76077:13
						state_d = 3'd1;
					else
						// Trace: design.sv:76079:13
						state_d = 3'd6;
				3'd7: begin
					// Trace: design.sv:76084:11
					state_d = next_state_after_idle_csb_active;
					// Trace: design.sv:76085:11
					command_ready_int = command_ready_idle_csb_active;
				end
				default: begin
					// Trace: design.sv:76088:11
					command_ready_int = 1'b0;
					// Trace: design.sv:76089:11
					state_d = 3'd0;
				end
			endcase
	end
	// Trace: design.sv:76100:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:76101:5
		if (!rst_ni) begin
			// Trace: design.sv:76102:7
			state_q <= 3'd0;
			// Trace: design.sv:76103:7
			clk_cntr_q <= 16'h0000;
		end
		else begin
			// Trace: design.sv:76105:7
			state_q <= (stall ? state_q : state_d);
			// Trace: design.sv:76106:7
			clk_cntr_q <= (stall ? clk_cntr_q : clk_cntr_d);
		end
	// Trace: design.sv:76110:3
	wire segment_rd_en;
	wire segment_rd_en_cpha0;
	reg segment_rd_en_cpha1;
	// Trace: design.sv:76112:3
	assign state_changing = state_q != state_d;
	// Trace: design.sv:76113:3
	assign byte_starting_cpha0 = (~sw_rst_i & state_changing) & ((state_d == 3'd1) | ((state_d == 3'd2) & (bit_cntr_q == 0)));
	// Trace: design.sv:76116:3
	assign bit_shifting_cpha0 = (~sw_rst_i & state_changing) & ((state_d == 3'd2) & (bit_cntr_q != 0));
	// Trace: design.sv:76118:3
	assign byte_ending_cpha0 = (~sw_rst_i & state_changing) & ((state_q == 3'd3) & (bit_cntr_q == 0));
	// Trace: design.sv:76121:3
	assign speed_cpha0 = cmd_speed_q;
	// Trace: design.sv:76122:3
	assign segment_rd_en_cpha0 = cmd_rd_en_q;
	// Trace: design.sv:76129:3
	// removed localparam type spi_host_cmd_pkg_speed_t
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:76130:5
		if (!rst_ni) begin
			// Trace: design.sv:76131:7
			byte_starting_cpha0_q <= 1'b0;
			// Trace: design.sv:76132:7
			byte_ending_cpha0_q <= 1'b0;
			// Trace: design.sv:76133:7
			bit_shifting_cpha0_q <= 1'b0;
			// Trace: design.sv:76134:7
			speed_cpha1 <= 2'b00;
			// Trace: design.sv:76135:7
			segment_rd_en_cpha1 <= 1'b0;
			// Trace: design.sv:76136:7
			new_command_cpha1 <= 1'b0;
		end
		else if (state_changing && !stall) begin
			// Trace: design.sv:76138:7
			byte_ending_cpha0_q <= byte_ending_cpha0;
			// Trace: design.sv:76139:7
			byte_starting_cpha0_q <= byte_starting_cpha0;
			// Trace: design.sv:76140:7
			bit_shifting_cpha0_q <= bit_shifting_cpha0;
			// Trace: design.sv:76141:7
			speed_cpha1 <= speed_cpha0;
			// Trace: design.sv:76142:7
			segment_rd_en_cpha1 <= segment_rd_en_cpha0;
			// Trace: design.sv:76143:7
			new_command_cpha1 <= new_command;
		end
	// Trace: design.sv:76150:3
	assign byte_starting_cpha1 = byte_starting_cpha0_q & state_changing;
	// Trace: design.sv:76151:3
	assign byte_ending_cpha1 = byte_ending_cpha0_q & state_changing;
	// Trace: design.sv:76152:3
	assign bit_shifting_cpha1 = bit_shifting_cpha0_q & state_changing;
	// Trace: design.sv:76154:3
	assign byte_starting = (cpha == 1'b0 ? byte_starting_cpha0 : byte_starting_cpha1);
	// Trace: design.sv:76157:3
	assign byte_ending = (cpha == 1'b0 ? byte_ending_cpha0 : byte_ending_cpha1);
	// Trace: design.sv:76160:3
	assign bit_shifting = (cpha == 1'b0 ? bit_shifting_cpha0 : bit_shifting_cpha1);
	// Trace: design.sv:76163:3
	assign speed_o = (cpha == 1'b0 ? speed_cpha0 : speed_cpha1);
	// Trace: design.sv:76166:3
	assign segment_rd_en = (cpha == 1'b0 ? segment_rd_en_cpha0 : segment_rd_en_cpha1);
	// Trace: design.sv:76169:3
	assign byte_cntr_early = (cpha == 1'b0 ? byte_cntr_cpha0_d : byte_cntr_cpha1_d);
	// Trace: design.sv:76171:3
	assign byte_cntr_late = (cpha == 1'b0 ? byte_cntr_cpha0_q : byte_cntr_cpha1_q);
	// Trace: design.sv:76174:3
	reg [2:0] shift_size;
	// Trace: design.sv:76175:3
	reg [2:0] start_bit;
	// Trace: design.sv:76177:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:76178:5
		if (!cmd_rd_en_d && !cmd_wr_en_d) begin
			// Trace: design.sv:76184:7
			shift_size = 0;
			// Trace: design.sv:76185:7
			start_bit = 3'h0;
		end
		else
			// Trace: design.sv:76187:7
			(* full_case, parallel_case *)
			case (cmd_speed_d)
				2'b00: begin
					// Trace: design.sv:76189:11
					shift_size = 3'h1;
					// Trace: design.sv:76190:11
					start_bit = 3'h7;
				end
				2'b01: begin
					// Trace: design.sv:76193:11
					shift_size = 3'h2;
					// Trace: design.sv:76194:11
					start_bit = 3'h6;
				end
				2'b10: begin
					// Trace: design.sv:76197:11
					shift_size = 3'h4;
					// Trace: design.sv:76198:11
					start_bit = 3'h4;
				end
				default: begin
					// Trace: design.sv:76202:11
					shift_size = 3'h1;
					// Trace: design.sv:76203:11
					start_bit = 3'h1;
				end
			endcase
	end
	// Trace: design.sv:76209:3
	assign bit_cntr_d = (sw_rst_i ? 3'h0 : (!fsm_en ? bit_cntr_q : (byte_starting ? start_bit : (bit_shifting ? bit_cntr_q - shift_size : bit_cntr_q))));
	// Trace: design.sv:76215:3
	assign last_bit = bit_cntr_q == 3'h0;
	// Trace: design.sv:76222:3
	assign last_byte = byte_cntr_cpha0_q == 24'h000000;
	// Trace: design.sv:76226:3
	assign byte_cntr_cpha0_d = (sw_rst_i ? 24'h000000 : (!fsm_en ? byte_cntr_cpha0_q : (new_command ? cmd_len_d : (byte_ending_cpha0 ? byte_cntr_cpha0_q - 1 : byte_cntr_cpha0_q))));
	// Trace: design.sv:76235:3
	assign byte_cntr_cpha1_d = (sw_rst_i ? 24'h000000 : (!fsm_en ? byte_cntr_cpha1_q : (new_command_cpha1 ? cmd_len_q : (byte_ending_cpha1 ? byte_cntr_cpha1_q - 1 : byte_cntr_cpha1_q))));
	// Trace: design.sv:76241:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:76242:5
		if (sw_rst_i)
			// Trace: design.sv:76243:7
			wait_cntr_d = 4'b0000;
		else if (!fsm_en)
			// Trace: design.sv:76245:7
			wait_cntr_d = wait_cntr_q;
		else if (state_changing)
			// Trace: design.sv:76247:7
			(* full_case, parallel_case *)
			case (state_d)
				3'd1:
					// Trace: design.sv:76249:12
					wait_cntr_d = csnlead;
				3'd4:
					// Trace: design.sv:76252:12
					wait_cntr_d = csntrail;
				3'd5:
					// Trace: design.sv:76255:12
					wait_cntr_d = csnidle;
				3'd6:
					// Trace: design.sv:76258:12
					wait_cntr_d = csnidle;
				default:
					// Trace: design.sv:76263:12
					wait_cntr_d = 4'b0000;
			endcase
		else if (wait_cntr_q == 0)
			// Trace: design.sv:76267:7
			wait_cntr_d = 4'h0;
		else
			// Trace: design.sv:76269:7
			wait_cntr_d = wait_cntr_q - 1;
	end
	// Trace: design.sv:76273:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:76274:5
		if (!rst_ni) begin
			// Trace: design.sv:76275:7
			bit_cntr_q <= 3'h0;
			// Trace: design.sv:76276:7
			byte_cntr_cpha0_q <= 24'h000000;
			// Trace: design.sv:76277:7
			byte_cntr_cpha1_q <= 24'h000000;
			// Trace: design.sv:76278:7
			wait_cntr_q <= 4'h0;
		end
		else begin
			// Trace: design.sv:76280:7
			bit_cntr_q <= (stall ? bit_cntr_q : bit_cntr_d);
			// Trace: design.sv:76281:7
			byte_cntr_cpha0_q <= (stall ? byte_cntr_cpha0_q : byte_cntr_cpha0_d);
			// Trace: design.sv:76282:7
			byte_cntr_cpha1_q <= (stall ? byte_cntr_cpha1_q : byte_cntr_cpha1_d);
			// Trace: design.sv:76283:7
			wait_cntr_q <= (stall ? wait_cntr_q : wait_cntr_d);
		end
	// Trace: design.sv:76287:3
	assign wr_en_internal = byte_starting & cmd_wr_en_d;
	// Trace: design.sv:76288:3
	assign shift_en_internal = bit_shifting;
	// Trace: design.sv:76290:3
	assign rd_en_internal = byte_ending & segment_rd_en;
	// Trace: design.sv:76291:3
	assign sample_en_d = byte_starting | shift_en_o;
	// Trace: design.sv:76292:3
	assign full_cyc_o = full_cyc;
	// Trace: design.sv:76293:3
	assign last_read_o = ((byte_cntr_late == 'h0) & rd_en_o) & sr_rd_ready_i;
	// Trace: design.sv:76295:3
	assign last_write_o = ((byte_cntr_early == 'h0) & wr_en_o) & sr_wr_ready_i;
	// Trace: design.sv:76297:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:76298:5
		if (!rst_ni) begin
			// Trace: design.sv:76299:7
			sample_en_q <= 1'b0;
			// Trace: design.sv:76300:7
			sample_en_q2 <= 1'b0;
		end
		else begin
			// Trace: design.sv:76302:7
			sample_en_q <= (fsm_en && !stall ? sample_en_d : sample_en_q);
			// Trace: design.sv:76303:7
			sample_en_q2 <= (fsm_en && !stall ? sample_en_q : sample_en_q2);
		end
	// Trace: design.sv:76307:3
	assign sample_en_internal = (full_cyc_o ? sample_en_q2 : sample_en_q);
	// Trace: design.sv:76309:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:76310:5
		(* full_case, parallel_case *)
		case (state_d)
			3'd1, 3'd2, 3'd3, 3'd7, 3'd4:
				// Trace: design.sv:76312:9
				csb_single_d = 1'b0;
			default:
				// Trace: design.sv:76314:9
				csb_single_d = 1'b1;
		endcase
	end
	// Trace: design.sv:76318:3
	assign sck_d = (cpol ? state_d != 3'd3 : state_d == 3'd3);
	// Trace: design.sv:76321:3
	assign sck_o = sck_q;
	// Trace: design.sv:76323:3
	prim_flop_en u_sck_flop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.en_i(~stall),
		.d_i(sck_d),
		.q_o(sck_q)
	);
	// Trace: design.sv:76331:3
	genvar _gv_ii_3;
	generate
		for (_gv_ii_3 = 0; _gv_ii_3 < NumCS; _gv_ii_3 = _gv_ii_3 + 1) begin : gen_csb_gen
			localparam ii = _gv_ii_3;
			// Trace: design.sv:76332:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: design.sv:76333:7
				if (!rst_ni)
					// Trace: design.sv:76334:9
					csb_q[ii] <= 1'b1;
				else
					// Trace: design.sv:76336:9
					csb_q[ii] <= (csid != ii ? 1'b1 : (!stall ? csb_single_d : csb_q[ii]));
		end
	endgenerate
	// Trace: design.sv:76343:3
	assign csb_o = csb_q;
	// Trace: design.sv:76345:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:76346:5
		if (&csb_o)
			// Trace: design.sv:76347:7
			sd_en_o[3:0] = 4'h0;
		else
			// Trace: design.sv:76349:7
			(* full_case, parallel_case *)
			case (speed_o)
				2'b00: begin
					// Trace: design.sv:76351:11
					sd_en_o[0] = 1'b1;
					// Trace: design.sv:76352:11
					sd_en_o[1] = 1'b0;
					// Trace: design.sv:76353:11
					sd_en_o[3:2] = 2'b00;
				end
				2'b01: begin
					// Trace: design.sv:76356:11
					sd_en_o[1:0] = {2 {cmd_wr_en_q}};
					// Trace: design.sv:76357:11
					sd_en_o[3:2] = 2'b00;
				end
				2'b10:
					// Trace: design.sv:76360:11
					sd_en_o[3:0] = {4 {cmd_wr_en_q}};
				default:
					// Trace: design.sv:76364:11
					sd_en_o[3:0] = 4'h0;
			endcase
	end
	initial _sv2v_0 = 0;
endmodule
module spi_host_core (
	clk_i,
	rst_ni,
	command_i,
	command_valid_i,
	command_ready_o,
	en_i,
	tx_data_i,
	tx_be_i,
	tx_valid_i,
	tx_ready_o,
	rx_data_o,
	rx_valid_o,
	rx_ready_i,
	sw_rst_i,
	sck_o,
	csb_o,
	sd_o,
	sd_en_o,
	sd_i,
	rx_stall_o,
	tx_stall_o,
	active_o
);
	// Trace: design.sv:76387:14
	parameter signed [31:0] NumCS = 1;
	// Trace: design.sv:76389:3
	input clk_i;
	// Trace: design.sv:76390:3
	input rst_ni;
	// Trace: design.sv:76392:3
	function automatic integer prim_util_pkg_vbits;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:74:36
		input integer value;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:85:5
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] spi_host_reg_pkg_NumCS = 2;
	localparam signed [31:0] spi_host_cmd_pkg_CSW = prim_util_pkg_vbits(spi_host_reg_pkg_NumCS);
	// removed localparam type spi_host_cmd_pkg_configopts_t
	// removed localparam type spi_host_cmd_pkg_segment_t
	// removed localparam type spi_host_cmd_pkg_command_t
	input wire [spi_host_cmd_pkg_CSW + 59:0] command_i;
	// Trace: design.sv:76393:3
	input command_valid_i;
	// Trace: design.sv:76394:3
	output wire command_ready_o;
	// Trace: design.sv:76395:3
	input en_i;
	// Trace: design.sv:76397:3
	input [31:0] tx_data_i;
	// Trace: design.sv:76398:3
	input [3:0] tx_be_i;
	// Trace: design.sv:76399:3
	input tx_valid_i;
	// Trace: design.sv:76400:3
	output wire tx_ready_o;
	// Trace: design.sv:76402:3
	output wire [31:0] rx_data_o;
	// Trace: design.sv:76403:3
	output wire rx_valid_o;
	// Trace: design.sv:76404:3
	input rx_ready_i;
	// Trace: design.sv:76406:3
	input sw_rst_i;
	// Trace: design.sv:76409:3
	output wire sck_o;
	// Trace: design.sv:76410:3
	output wire [NumCS - 1:0] csb_o;
	// Trace: design.sv:76411:3
	output wire [3:0] sd_o;
	// Trace: design.sv:76412:3
	output wire [3:0] sd_en_o;
	// Trace: design.sv:76413:3
	input [3:0] sd_i;
	// Trace: design.sv:76416:3
	output wire rx_stall_o;
	// Trace: design.sv:76417:3
	output wire tx_stall_o;
	// Trace: design.sv:76418:3
	output wire active_o;
	// Trace: design.sv:76421:3
	wire rx_valid_sr;
	// Trace: design.sv:76422:3
	wire rx_ready_sr;
	// Trace: design.sv:76423:3
	wire rx_last_sr;
	// Trace: design.sv:76424:3
	wire [7:0] rx_data_sr;
	// Trace: design.sv:76425:3
	wire tx_valid_sr;
	// Trace: design.sv:76426:3
	wire tx_ready_sr;
	// Trace: design.sv:76427:3
	wire tx_flush_sr;
	// Trace: design.sv:76428:3
	wire [7:0] tx_data_sr;
	// Trace: design.sv:76430:3
	wire wr_en;
	// Trace: design.sv:76431:3
	wire rd_en;
	// Trace: design.sv:76432:3
	wire wr_ready;
	// Trace: design.sv:76433:3
	wire rd_ready;
	// Trace: design.sv:76435:3
	wire sample_en;
	// Trace: design.sv:76436:3
	wire shift_en;
	// Trace: design.sv:76437:3
	wire [1:0] speed;
	// Trace: design.sv:76438:3
	wire full_cyc;
	// Trace: design.sv:76439:3
	wire last_read;
	// Trace: design.sv:76440:3
	wire last_write;
	// Trace: design.sv:76442:3
	spi_host_byte_merge u_merge(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.byte_i(rx_data_sr),
		.byte_last_i(rx_last_sr),
		.byte_valid_i(rx_valid_sr),
		.byte_ready_o(rx_ready_sr),
		.word_o(rx_data_o),
		.word_valid_o(rx_valid_o),
		.word_ready_i(rx_ready_i),
		.sw_rst_i(sw_rst_i)
	);
	// Trace: design.sv:76455:3
	spi_host_byte_select u_select(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.word_i(tx_data_i),
		.word_be_i(tx_be_i),
		.word_valid_i(tx_valid_i),
		.word_ready_o(tx_ready_o),
		.byte_o(tx_data_sr),
		.byte_valid_o(tx_valid_sr),
		.byte_ready_i(tx_ready_sr),
		.flush_i(tx_flush_sr),
		.sw_rst_i(sw_rst_i)
	);
	// Trace: design.sv:76469:3
	spi_host_shift_register u_shift_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_en_i(wr_en),
		.wr_ready_o(wr_ready),
		.rd_en_i(rd_en),
		.rd_ready_o(rd_ready),
		.speed_i(speed),
		.shift_en_i(shift_en),
		.sample_en_i(sample_en),
		.last_read_i(last_read),
		.last_write_i(last_write),
		.full_cyc_i(full_cyc),
		.tx_data_i(tx_data_sr),
		.tx_valid_i(tx_valid_sr),
		.tx_ready_o(tx_ready_sr),
		.tx_flush_o(tx_flush_sr),
		.rx_data_o(rx_data_sr),
		.rx_valid_o(rx_valid_sr),
		.rx_ready_i(rx_ready_sr),
		.rx_last_o(rx_last_sr),
		.sw_rst_i(sw_rst_i),
		.sd_o(sd_o),
		.sd_i(sd_i)
	);
	// Trace: design.sv:76495:3
	spi_host_fsm #(.NumCS(NumCS)) u_fsm(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.en_i(en_i),
		.command_i(command_i),
		.command_valid_i(command_valid_i),
		.command_ready_o(command_ready_o),
		.sck_o(sck_o),
		.csb_o(csb_o),
		.sd_en_o(sd_en_o),
		.last_read_o(last_read),
		.last_write_o(last_write),
		.wr_en_o(wr_en),
		.sr_wr_ready_i(wr_ready),
		.rd_en_o(rd_en),
		.sr_rd_ready_i(rd_ready),
		.sample_en_o(sample_en),
		.shift_en_o(shift_en),
		.speed_o(speed),
		.full_cyc_o(full_cyc),
		.sw_rst_i(sw_rst_i),
		.rx_stall_o(rx_stall_o),
		.tx_stall_o(tx_stall_o),
		.active_o(active_o)
	);
endmodule
module spi_host_command_queue (
	clk_i,
	rst_ni,
	command_i,
	command_valid_i,
	command_busy_o,
	core_command_o,
	core_command_valid_o,
	core_command_ready_i,
	qd_o,
	error_busy_o,
	sw_rst_i
);
	// Trace: design.sv:76532:13
	parameter signed [31:0] CmdDepth = 4;
	// Trace: design.sv:76534:3
	input clk_i;
	// Trace: design.sv:76535:3
	input rst_ni;
	// Trace: design.sv:76537:3
	function automatic integer prim_util_pkg_vbits;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:74:36
		input integer value;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:85:5
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] spi_host_reg_pkg_NumCS = 2;
	localparam signed [31:0] spi_host_cmd_pkg_CSW = prim_util_pkg_vbits(spi_host_reg_pkg_NumCS);
	// removed localparam type spi_host_cmd_pkg_configopts_t
	// removed localparam type spi_host_cmd_pkg_segment_t
	// removed localparam type spi_host_cmd_pkg_command_t
	input wire [spi_host_cmd_pkg_CSW + 59:0] command_i;
	// Trace: design.sv:76538:3
	input command_valid_i;
	// Trace: design.sv:76539:3
	output wire command_busy_o;
	// Trace: design.sv:76541:3
	output wire [spi_host_cmd_pkg_CSW + 59:0] core_command_o;
	// Trace: design.sv:76542:3
	output wire core_command_valid_o;
	// Trace: design.sv:76543:3
	input core_command_ready_i;
	// Trace: design.sv:76545:3
	output wire [3:0] qd_o;
	// Trace: design.sv:76547:3
	output wire error_busy_o;
	// Trace: design.sv:76549:3
	input sw_rst_i;
	// Trace: design.sv:76552:3
	localparam signed [31:0] CmdDepthW = prim_util_pkg_vbits(CmdDepth + 1);
	// Trace: design.sv:76554:3
	wire command_ready;
	// Trace: design.sv:76556:3
	assign command_busy_o = ~command_ready;
	// Trace: design.sv:76557:3
	assign error_busy_o = command_valid_i & command_busy_o;
	// Trace: design.sv:76559:3
	wire [CmdDepthW - 1:0] cmd_depth;
	// Trace: design.sv:76561:3
	localparam signed [31:0] spi_host_cmd_pkg_CmdSize = spi_host_cmd_pkg_CSW + 60;
	prim_fifo_sync #(
		.Width(spi_host_cmd_pkg_CmdSize),
		.Pass(1),
		.Depth(CmdDepth)
	) cmd_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(sw_rst_i),
		.wvalid_i(command_valid_i),
		.wready_o(command_ready),
		.wdata_i(command_i),
		.rvalid_o(core_command_valid_o),
		.rready_i(core_command_ready_i),
		.rdata_o(core_command_o),
		.full_o(),
		.depth_o(cmd_depth)
	);
	// Trace: design.sv:76579:3
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	assign qd_o = sv2v_cast_4(cmd_depth);
endmodule
module spi_host_data_fifos (
	clk_i,
	rst_ni,
	tx_data_i,
	tx_be_i,
	tx_valid_i,
	tx_ready_o,
	tx_watermark_i,
	core_tx_data_o,
	core_tx_be_o,
	core_tx_valid_o,
	core_tx_ready_i,
	core_rx_data_i,
	core_rx_valid_i,
	core_rx_ready_o,
	rx_data_o,
	rx_valid_o,
	rx_ready_i,
	rx_watermark_i,
	sw_rst_i,
	tx_empty_o,
	tx_full_o,
	tx_qd_o,
	tx_wm_o,
	rx_empty_o,
	rx_full_o,
	rx_qd_o,
	rx_wm_o
);
	// Trace: design.sv:76590:13
	parameter signed [31:0] TxDepth = 72;
	// Trace: design.sv:76591:13
	parameter signed [31:0] RxDepth = 64;
	// Trace: design.sv:76592:13
	parameter [0:0] SwapBytes = 0;
	// Trace: design.sv:76594:3
	input clk_i;
	// Trace: design.sv:76595:3
	input rst_ni;
	// Trace: design.sv:76597:3
	input [31:0] tx_data_i;
	// Trace: design.sv:76598:3
	input [3:0] tx_be_i;
	// Trace: design.sv:76599:3
	input tx_valid_i;
	// Trace: design.sv:76600:3
	output wire tx_ready_o;
	// Trace: design.sv:76601:3
	input [7:0] tx_watermark_i;
	// Trace: design.sv:76603:3
	output wire [31:0] core_tx_data_o;
	// Trace: design.sv:76604:3
	output wire [3:0] core_tx_be_o;
	// Trace: design.sv:76605:3
	output wire core_tx_valid_o;
	// Trace: design.sv:76606:3
	input core_tx_ready_i;
	// Trace: design.sv:76608:3
	input [31:0] core_rx_data_i;
	// Trace: design.sv:76609:3
	input core_rx_valid_i;
	// Trace: design.sv:76610:3
	output wire core_rx_ready_o;
	// Trace: design.sv:76612:3
	output wire [31:0] rx_data_o;
	// Trace: design.sv:76613:3
	output wire rx_valid_o;
	// Trace: design.sv:76614:3
	input rx_ready_i;
	// Trace: design.sv:76615:3
	input [7:0] rx_watermark_i;
	// Trace: design.sv:76617:3
	input sw_rst_i;
	// Trace: design.sv:76619:3
	output wire tx_empty_o;
	// Trace: design.sv:76620:3
	output wire tx_full_o;
	// Trace: design.sv:76621:3
	output wire [7:0] tx_qd_o;
	// Trace: design.sv:76622:3
	output wire tx_wm_o;
	// Trace: design.sv:76623:3
	output wire rx_empty_o;
	// Trace: design.sv:76624:3
	output wire rx_full_o;
	// Trace: design.sv:76625:3
	output wire [7:0] rx_qd_o;
	// Trace: design.sv:76626:3
	output wire rx_wm_o;
	// Trace: design.sv:76629:3
	function automatic integer prim_util_pkg_vbits;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:74:36
		input integer value;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:85:5
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] RxDepthW = prim_util_pkg_vbits(RxDepth + 1);
	// Trace: design.sv:76630:3
	localparam signed [31:0] TxDepthW = prim_util_pkg_vbits(TxDepth + 1);
	// Trace: design.sv:76632:3
	wire [31:0] tx_data_ordered;
	// Trace: design.sv:76633:3
	wire [3:0] tx_be_ordered;
	// Trace: design.sv:76634:3
	wire [31:0] rx_data_unordered;
	// Trace: design.sv:76636:3
	generate
		if (SwapBytes) begin : gen_swap
			// Trace: design.sv:76637:5
			function automatic [31:0] _sv2v_strm_AB923;
				input reg [31:0] inp;
				reg [31:0] _sv2v_strm_39B78_inp;
				reg [31:0] _sv2v_strm_39B78_out;
				integer _sv2v_strm_39B78_idx;
				begin
					_sv2v_strm_39B78_inp = {inp};
					for (_sv2v_strm_39B78_idx = 0; _sv2v_strm_39B78_idx <= 24; _sv2v_strm_39B78_idx = _sv2v_strm_39B78_idx + 8)
						_sv2v_strm_39B78_out[31 - _sv2v_strm_39B78_idx-:8] = _sv2v_strm_39B78_inp[_sv2v_strm_39B78_idx+:8];
					_sv2v_strm_AB923 = _sv2v_strm_39B78_out << 0;
				end
			endfunction
			assign tx_data_ordered = _sv2v_strm_AB923({tx_data_i});
			// Trace: design.sv:76638:5
			function automatic [3:0] _sv2v_strm_2D57E;
				input reg [3:0] inp;
				reg [3:0] _sv2v_strm_BEEC1_inp;
				reg [3:0] _sv2v_strm_BEEC1_out;
				integer _sv2v_strm_BEEC1_idx;
				begin
					_sv2v_strm_BEEC1_inp = {inp};
					for (_sv2v_strm_BEEC1_idx = 0; _sv2v_strm_BEEC1_idx <= 3; _sv2v_strm_BEEC1_idx = _sv2v_strm_BEEC1_idx + 1)
						_sv2v_strm_BEEC1_out[3 - _sv2v_strm_BEEC1_idx-:1] = _sv2v_strm_BEEC1_inp[_sv2v_strm_BEEC1_idx+:1];
					_sv2v_strm_2D57E = _sv2v_strm_BEEC1_out << 0;
				end
			endfunction
			assign tx_be_ordered = _sv2v_strm_2D57E({tx_be_i});
			// Trace: design.sv:76639:5
			function automatic [31:0] _sv2v_strm_695D0;
				input reg [31:0] inp;
				reg [31:0] _sv2v_strm_39B78_inp;
				reg [31:0] _sv2v_strm_39B78_out;
				integer _sv2v_strm_39B78_idx;
				begin
					_sv2v_strm_39B78_inp = {inp};
					for (_sv2v_strm_39B78_idx = 0; _sv2v_strm_39B78_idx <= 24; _sv2v_strm_39B78_idx = _sv2v_strm_39B78_idx + 8)
						_sv2v_strm_39B78_out[31 - _sv2v_strm_39B78_idx-:8] = _sv2v_strm_39B78_inp[_sv2v_strm_39B78_idx+:8];
					_sv2v_strm_695D0 = _sv2v_strm_39B78_out << 0;
				end
			endfunction
			assign rx_data_o = _sv2v_strm_695D0({rx_data_unordered});
		end
		else begin : gen_do_not_swap
			// Trace: design.sv:76641:5
			assign tx_data_ordered = tx_data_i;
			// Trace: design.sv:76642:5
			assign tx_be_ordered = tx_be_i;
			// Trace: design.sv:76643:5
			assign rx_data_o = rx_data_unordered;
		end
	endgenerate
	// Trace: design.sv:76646:3
	wire [35:0] tx_data_be;
	// Trace: design.sv:76647:3
	wire [35:0] core_tx_data_be;
	// Trace: design.sv:76649:3
	wire [TxDepthW - 1:0] tx_depth;
	// Trace: design.sv:76651:3
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	assign tx_qd_o = sv2v_cast_8(tx_depth);
	// Trace: design.sv:76653:3
	assign tx_data_be = {tx_data_ordered, tx_be_ordered};
	// Trace: design.sv:76654:3
	assign {core_tx_data_o, core_tx_be_o} = core_tx_data_be;
	// Trace: design.sv:76656:3
	prim_fifo_sync #(
		.Width(36),
		.Pass(1),
		.Depth(TxDepth)
	) u_tx_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(sw_rst_i),
		.wvalid_i(tx_valid_i),
		.wready_o(tx_ready_o),
		.wdata_i(tx_data_be),
		.rvalid_o(core_tx_valid_o),
		.rready_i(core_tx_ready_i),
		.rdata_o(core_tx_data_be),
		.full_o(),
		.depth_o(tx_depth)
	);
	// Trace: design.sv:76674:3
	wire [RxDepthW - 1:0] rx_depth;
	// Trace: design.sv:76676:3
	assign rx_qd_o = sv2v_cast_8(rx_depth);
	// Trace: design.sv:76678:3
	prim_fifo_sync #(
		.Width(32),
		.Pass(1),
		.Depth(RxDepth)
	) u_rx_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(sw_rst_i),
		.wvalid_i(core_rx_valid_i),
		.wready_o(core_rx_ready_o),
		.wdata_i(core_rx_data_i),
		.rvalid_o(rx_valid_o),
		.rready_i(rx_ready_i),
		.rdata_o(rx_data_unordered),
		.full_o(),
		.depth_o(rx_depth)
	);
	// Trace: design.sv:76696:3
	assign tx_empty_o = tx_qd_o == 0;
	// Trace: design.sv:76697:3
	assign rx_empty_o = rx_qd_o == 0;
	// Trace: design.sv:76698:3
	function automatic signed [7:0] sv2v_cast_8_signed;
		input reg signed [7:0] inp;
		sv2v_cast_8_signed = inp;
	endfunction
	assign tx_full_o = tx_qd_o >= sv2v_cast_8_signed(TxDepth);
	// Trace: design.sv:76699:3
	assign rx_full_o = rx_qd_o >= sv2v_cast_8_signed(RxDepth);
	// Trace: design.sv:76700:3
	assign tx_wm_o = tx_qd_o < tx_watermark_i;
	// Trace: design.sv:76701:3
	assign rx_wm_o = rx_qd_o >= rx_watermark_i;
endmodule
module spi_host_reg_top_3E795 (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	reg_req_win_o,
	reg_rsp_win_i,
	reg2hw,
	hw2reg,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:76714:20
	// removed localparam type reg_req_t
	// Trace: design.sv:76715:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:76716:15
	parameter signed [31:0] AW = 6;
	// Trace: design.sv:76718:3
	input clk_i;
	// Trace: design.sv:76719:3
	input rst_ni;
	// Trace: design.sv:76720:3
	input wire [69:0] reg_req_i;
	// Trace: design.sv:76721:3
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:76724:3
	output wire [139:0] reg_req_win_o;
	// Trace: design.sv:76725:3
	input wire [67:0] reg_rsp_win_i;
	// Trace: design.sv:76728:3
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_alert_test_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_command_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_configopts_mreg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_control_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_csid_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_error_enable_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_error_status_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_event_enable_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_intr_enable_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_intr_state_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_intr_test_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_t
	output wire [172:0] reg2hw;
	// Trace: design.sv:76729:3
	// removed localparam type spi_host_reg_pkg_spi_host_hw2reg_error_status_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_hw2reg_intr_state_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_hw2reg_status_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_hw2reg_t
	input wire [60:0] hw2reg;
	// Trace: design.sv:76733:3
	input devmode_i;
	// Trace: design.sv:76736:3
	// removed import spi_host_reg_pkg::*;
	// Trace: design.sv:76738:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:76739:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:76742:3
	wire reg_we;
	// Trace: design.sv:76743:3
	wire reg_re;
	// Trace: design.sv:76744:3
	wire [AW - 1:0] reg_addr;
	// Trace: design.sv:76745:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:76746:3
	wire [3:0] reg_be;
	// Trace: design.sv:76747:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:76748:3
	wire reg_error;
	// Trace: design.sv:76750:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:76752:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:76755:3
	wire [69:0] reg_intf_req;
	// Trace: design.sv:76756:3
	wire [33:0] reg_intf_rsp;
	// Trace: design.sv:76759:3
	reg [1:0] reg_steer;
	// Trace: design.sv:76761:3
	wire [209:0] reg_intf_demux_req;
	// Trace: design.sv:76762:3
	wire [101:0] reg_intf_demux_rsp;
	// Trace: design.sv:76765:3
	assign reg_intf_req = reg_intf_demux_req[140+:70];
	// Trace: design.sv:76766:3
	assign reg_intf_demux_rsp[68+:34] = reg_intf_rsp;
	// Trace: design.sv:76768:3
	assign reg_req_win_o[0+:70] = reg_intf_demux_req[0+:70];
	// Trace: design.sv:76769:3
	assign reg_intf_demux_rsp[0+:34] = reg_rsp_win_i[0+:34];
	// Trace: design.sv:76770:3
	assign reg_req_win_o[70+:70] = reg_intf_demux_req[70+:70];
	// Trace: design.sv:76771:3
	assign reg_intf_demux_rsp[34+:34] = reg_rsp_win_i[34+:34];
	// Trace: design.sv:76774:3
	reg_demux_64ED6 #(.NoPorts(3)) i_reg_demux(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.in_req_i(reg_req_i),
		.in_rsp_o(reg_rsp_o),
		.out_req_o(reg_intf_demux_req),
		.out_rsp_i(reg_intf_demux_rsp),
		.in_select_i(reg_steer)
	);
	// Trace: design.sv:76790:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:76791:5
		reg_steer = 2;
		// Trace: design.sv:76794:5
		if ((reg_req_i[31 + AW:32] >= 40) && (reg_req_i[31 + AW:32] < 44))
			// Trace: design.sv:76795:7
			reg_steer = 0;
		if ((reg_req_i[31 + AW:32] >= 44) && (reg_req_i[31 + AW:32] < 48))
			// Trace: design.sv:76798:7
			reg_steer = 1;
	end
	// Trace: design.sv:76803:3
	assign reg_we = reg_intf_req[69] & reg_intf_req[68];
	// Trace: design.sv:76804:3
	assign reg_re = reg_intf_req[69] & ~reg_intf_req[68];
	// Trace: design.sv:76805:3
	assign reg_addr = reg_intf_req[63-:32];
	// Trace: design.sv:76806:3
	assign reg_wdata = reg_intf_req[31-:32];
	// Trace: design.sv:76807:3
	assign reg_be = reg_intf_req[67-:4];
	// Trace: design.sv:76808:3
	assign reg_intf_rsp[31-:32] = reg_rdata;
	// Trace: design.sv:76809:3
	assign reg_intf_rsp[33] = reg_error;
	// Trace: design.sv:76810:3
	assign reg_intf_rsp[32] = 1'b1;
	// Trace: design.sv:76812:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:76813:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:76819:3
	wire intr_state_error_qs;
	// Trace: design.sv:76820:3
	wire intr_state_error_wd;
	// Trace: design.sv:76821:3
	wire intr_state_error_we;
	// Trace: design.sv:76822:3
	wire intr_state_spi_event_qs;
	// Trace: design.sv:76823:3
	wire intr_state_spi_event_wd;
	// Trace: design.sv:76824:3
	wire intr_state_spi_event_we;
	// Trace: design.sv:76825:3
	wire intr_enable_error_qs;
	// Trace: design.sv:76826:3
	wire intr_enable_error_wd;
	// Trace: design.sv:76827:3
	wire intr_enable_error_we;
	// Trace: design.sv:76828:3
	wire intr_enable_spi_event_qs;
	// Trace: design.sv:76829:3
	wire intr_enable_spi_event_wd;
	// Trace: design.sv:76830:3
	wire intr_enable_spi_event_we;
	// Trace: design.sv:76831:3
	wire intr_test_error_wd;
	// Trace: design.sv:76832:3
	wire intr_test_error_we;
	// Trace: design.sv:76833:3
	wire intr_test_spi_event_wd;
	// Trace: design.sv:76834:3
	wire intr_test_spi_event_we;
	// Trace: design.sv:76835:3
	wire alert_test_wd;
	// Trace: design.sv:76836:3
	wire alert_test_we;
	// Trace: design.sv:76837:3
	wire [7:0] control_rx_watermark_qs;
	// Trace: design.sv:76838:3
	wire [7:0] control_rx_watermark_wd;
	// Trace: design.sv:76839:3
	wire control_rx_watermark_we;
	// Trace: design.sv:76840:3
	wire [7:0] control_tx_watermark_qs;
	// Trace: design.sv:76841:3
	wire [7:0] control_tx_watermark_wd;
	// Trace: design.sv:76842:3
	wire control_tx_watermark_we;
	// Trace: design.sv:76843:3
	wire control_output_en_qs;
	// Trace: design.sv:76844:3
	wire control_output_en_wd;
	// Trace: design.sv:76845:3
	wire control_output_en_we;
	// Trace: design.sv:76846:3
	wire control_sw_rst_qs;
	// Trace: design.sv:76847:3
	wire control_sw_rst_wd;
	// Trace: design.sv:76848:3
	wire control_sw_rst_we;
	// Trace: design.sv:76849:3
	wire control_spien_qs;
	// Trace: design.sv:76850:3
	wire control_spien_wd;
	// Trace: design.sv:76851:3
	wire control_spien_we;
	// Trace: design.sv:76852:3
	wire [7:0] status_txqd_qs;
	// Trace: design.sv:76853:3
	wire [7:0] status_rxqd_qs;
	// Trace: design.sv:76854:3
	wire [3:0] status_cmdqd_qs;
	// Trace: design.sv:76855:3
	wire status_rxwm_qs;
	// Trace: design.sv:76856:3
	wire status_byteorder_qs;
	// Trace: design.sv:76857:3
	wire status_rxstall_qs;
	// Trace: design.sv:76858:3
	wire status_rxempty_qs;
	// Trace: design.sv:76859:3
	wire status_rxfull_qs;
	// Trace: design.sv:76860:3
	wire status_txwm_qs;
	// Trace: design.sv:76861:3
	wire status_txstall_qs;
	// Trace: design.sv:76862:3
	wire status_txempty_qs;
	// Trace: design.sv:76863:3
	wire status_txfull_qs;
	// Trace: design.sv:76864:3
	wire status_active_qs;
	// Trace: design.sv:76865:3
	wire status_ready_qs;
	// Trace: design.sv:76866:3
	wire [15:0] configopts_0_clkdiv_0_qs;
	// Trace: design.sv:76867:3
	wire [15:0] configopts_0_clkdiv_0_wd;
	// Trace: design.sv:76868:3
	wire configopts_0_clkdiv_0_we;
	// Trace: design.sv:76869:3
	wire [3:0] configopts_0_csnidle_0_qs;
	// Trace: design.sv:76870:3
	wire [3:0] configopts_0_csnidle_0_wd;
	// Trace: design.sv:76871:3
	wire configopts_0_csnidle_0_we;
	// Trace: design.sv:76872:3
	wire [3:0] configopts_0_csntrail_0_qs;
	// Trace: design.sv:76873:3
	wire [3:0] configopts_0_csntrail_0_wd;
	// Trace: design.sv:76874:3
	wire configopts_0_csntrail_0_we;
	// Trace: design.sv:76875:3
	wire [3:0] configopts_0_csnlead_0_qs;
	// Trace: design.sv:76876:3
	wire [3:0] configopts_0_csnlead_0_wd;
	// Trace: design.sv:76877:3
	wire configopts_0_csnlead_0_we;
	// Trace: design.sv:76878:3
	wire configopts_0_fullcyc_0_qs;
	// Trace: design.sv:76879:3
	wire configopts_0_fullcyc_0_wd;
	// Trace: design.sv:76880:3
	wire configopts_0_fullcyc_0_we;
	// Trace: design.sv:76881:3
	wire configopts_0_cpha_0_qs;
	// Trace: design.sv:76882:3
	wire configopts_0_cpha_0_wd;
	// Trace: design.sv:76883:3
	wire configopts_0_cpha_0_we;
	// Trace: design.sv:76884:3
	wire configopts_0_cpol_0_qs;
	// Trace: design.sv:76885:3
	wire configopts_0_cpol_0_wd;
	// Trace: design.sv:76886:3
	wire configopts_0_cpol_0_we;
	// Trace: design.sv:76887:3
	wire [15:0] configopts_1_clkdiv_1_qs;
	// Trace: design.sv:76888:3
	wire [15:0] configopts_1_clkdiv_1_wd;
	// Trace: design.sv:76889:3
	wire configopts_1_clkdiv_1_we;
	// Trace: design.sv:76890:3
	wire [3:0] configopts_1_csnidle_1_qs;
	// Trace: design.sv:76891:3
	wire [3:0] configopts_1_csnidle_1_wd;
	// Trace: design.sv:76892:3
	wire configopts_1_csnidle_1_we;
	// Trace: design.sv:76893:3
	wire [3:0] configopts_1_csntrail_1_qs;
	// Trace: design.sv:76894:3
	wire [3:0] configopts_1_csntrail_1_wd;
	// Trace: design.sv:76895:3
	wire configopts_1_csntrail_1_we;
	// Trace: design.sv:76896:3
	wire [3:0] configopts_1_csnlead_1_qs;
	// Trace: design.sv:76897:3
	wire [3:0] configopts_1_csnlead_1_wd;
	// Trace: design.sv:76898:3
	wire configopts_1_csnlead_1_we;
	// Trace: design.sv:76899:3
	wire configopts_1_fullcyc_1_qs;
	// Trace: design.sv:76900:3
	wire configopts_1_fullcyc_1_wd;
	// Trace: design.sv:76901:3
	wire configopts_1_fullcyc_1_we;
	// Trace: design.sv:76902:3
	wire configopts_1_cpha_1_qs;
	// Trace: design.sv:76903:3
	wire configopts_1_cpha_1_wd;
	// Trace: design.sv:76904:3
	wire configopts_1_cpha_1_we;
	// Trace: design.sv:76905:3
	wire configopts_1_cpol_1_qs;
	// Trace: design.sv:76906:3
	wire configopts_1_cpol_1_wd;
	// Trace: design.sv:76907:3
	wire configopts_1_cpol_1_we;
	// Trace: design.sv:76908:3
	wire [31:0] csid_qs;
	// Trace: design.sv:76909:3
	wire [31:0] csid_wd;
	// Trace: design.sv:76910:3
	wire csid_we;
	// Trace: design.sv:76911:3
	wire [23:0] command_len_wd;
	// Trace: design.sv:76912:3
	wire command_len_we;
	// Trace: design.sv:76913:3
	wire command_csaat_wd;
	// Trace: design.sv:76914:3
	wire command_csaat_we;
	// Trace: design.sv:76915:3
	wire [1:0] command_speed_wd;
	// Trace: design.sv:76916:3
	wire command_speed_we;
	// Trace: design.sv:76917:3
	wire [1:0] command_direction_wd;
	// Trace: design.sv:76918:3
	wire command_direction_we;
	// Trace: design.sv:76919:3
	wire error_enable_cmdbusy_qs;
	// Trace: design.sv:76920:3
	wire error_enable_cmdbusy_wd;
	// Trace: design.sv:76921:3
	wire error_enable_cmdbusy_we;
	// Trace: design.sv:76922:3
	wire error_enable_overflow_qs;
	// Trace: design.sv:76923:3
	wire error_enable_overflow_wd;
	// Trace: design.sv:76924:3
	wire error_enable_overflow_we;
	// Trace: design.sv:76925:3
	wire error_enable_underflow_qs;
	// Trace: design.sv:76926:3
	wire error_enable_underflow_wd;
	// Trace: design.sv:76927:3
	wire error_enable_underflow_we;
	// Trace: design.sv:76928:3
	wire error_enable_cmdinval_qs;
	// Trace: design.sv:76929:3
	wire error_enable_cmdinval_wd;
	// Trace: design.sv:76930:3
	wire error_enable_cmdinval_we;
	// Trace: design.sv:76931:3
	wire error_enable_csidinval_qs;
	// Trace: design.sv:76932:3
	wire error_enable_csidinval_wd;
	// Trace: design.sv:76933:3
	wire error_enable_csidinval_we;
	// Trace: design.sv:76934:3
	wire error_status_cmdbusy_qs;
	// Trace: design.sv:76935:3
	wire error_status_cmdbusy_wd;
	// Trace: design.sv:76936:3
	wire error_status_cmdbusy_we;
	// Trace: design.sv:76937:3
	wire error_status_overflow_qs;
	// Trace: design.sv:76938:3
	wire error_status_overflow_wd;
	// Trace: design.sv:76939:3
	wire error_status_overflow_we;
	// Trace: design.sv:76940:3
	wire error_status_underflow_qs;
	// Trace: design.sv:76941:3
	wire error_status_underflow_wd;
	// Trace: design.sv:76942:3
	wire error_status_underflow_we;
	// Trace: design.sv:76943:3
	wire error_status_cmdinval_qs;
	// Trace: design.sv:76944:3
	wire error_status_cmdinval_wd;
	// Trace: design.sv:76945:3
	wire error_status_cmdinval_we;
	// Trace: design.sv:76946:3
	wire error_status_csidinval_qs;
	// Trace: design.sv:76947:3
	wire error_status_csidinval_wd;
	// Trace: design.sv:76948:3
	wire error_status_csidinval_we;
	// Trace: design.sv:76949:3
	wire error_status_accessinval_qs;
	// Trace: design.sv:76950:3
	wire error_status_accessinval_wd;
	// Trace: design.sv:76951:3
	wire error_status_accessinval_we;
	// Trace: design.sv:76952:3
	wire event_enable_rxfull_qs;
	// Trace: design.sv:76953:3
	wire event_enable_rxfull_wd;
	// Trace: design.sv:76954:3
	wire event_enable_rxfull_we;
	// Trace: design.sv:76955:3
	wire event_enable_txempty_qs;
	// Trace: design.sv:76956:3
	wire event_enable_txempty_wd;
	// Trace: design.sv:76957:3
	wire event_enable_txempty_we;
	// Trace: design.sv:76958:3
	wire event_enable_rxwm_qs;
	// Trace: design.sv:76959:3
	wire event_enable_rxwm_wd;
	// Trace: design.sv:76960:3
	wire event_enable_rxwm_we;
	// Trace: design.sv:76961:3
	wire event_enable_txwm_qs;
	// Trace: design.sv:76962:3
	wire event_enable_txwm_wd;
	// Trace: design.sv:76963:3
	wire event_enable_txwm_we;
	// Trace: design.sv:76964:3
	wire event_enable_ready_qs;
	// Trace: design.sv:76965:3
	wire event_enable_ready_wd;
	// Trace: design.sv:76966:3
	wire event_enable_ready_we;
	// Trace: design.sv:76967:3
	wire event_enable_idle_qs;
	// Trace: design.sv:76968:3
	wire event_enable_idle_wd;
	// Trace: design.sv:76969:3
	wire event_enable_idle_we;
	// Trace: design.sv:76975:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_error(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_error_we),
		.wd(intr_state_error_wd),
		.de(hw2reg[59]),
		.d(hw2reg[60]),
		.qe(),
		.q(reg2hw[172]),
		.qs(intr_state_error_qs)
	);
	// Trace: design.sv:77001:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_spi_event(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_spi_event_we),
		.wd(intr_state_spi_event_wd),
		.de(hw2reg[57]),
		.d(hw2reg[58]),
		.qe(),
		.q(reg2hw[171]),
		.qs(intr_state_spi_event_qs)
	);
	// Trace: design.sv:77029:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_error_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_error_d
	localparam [0:0] sv2v_uu_u_intr_enable_error_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_error(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_error_we),
		.wd(intr_enable_error_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_error_ext_d_0),
		.qe(),
		.q(reg2hw[170]),
		.qs(intr_enable_error_qs)
	);
	// Trace: design.sv:77055:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_spi_event_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_spi_event_d
	localparam [0:0] sv2v_uu_u_intr_enable_spi_event_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_spi_event(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_spi_event_we),
		.wd(intr_enable_spi_event_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_spi_event_ext_d_0),
		.qe(),
		.q(reg2hw[169]),
		.qs(intr_enable_spi_event_qs)
	);
	// Trace: design.sv:77083:3
	localparam [31:0] sv2v_uu_u_intr_test_error_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_error_d
	localparam [0:0] sv2v_uu_u_intr_test_error_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_error(
		.re(1'b0),
		.we(intr_test_error_we),
		.wd(intr_test_error_wd),
		.d(sv2v_uu_u_intr_test_error_ext_d_0),
		.qre(),
		.qe(reg2hw[167]),
		.q(reg2hw[168]),
		.qs()
	);
	// Trace: design.sv:77098:3
	localparam [31:0] sv2v_uu_u_intr_test_spi_event_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_spi_event_d
	localparam [0:0] sv2v_uu_u_intr_test_spi_event_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_spi_event(
		.re(1'b0),
		.we(intr_test_spi_event_we),
		.wd(intr_test_spi_event_wd),
		.d(sv2v_uu_u_intr_test_spi_event_ext_d_0),
		.qre(),
		.qe(reg2hw[165]),
		.q(reg2hw[166]),
		.qs()
	);
	// Trace: design.sv:77114:3
	localparam [31:0] sv2v_uu_u_alert_test_DW = 1;
	// removed localparam type sv2v_uu_u_alert_test_d
	localparam [0:0] sv2v_uu_u_alert_test_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_alert_test(
		.re(1'b0),
		.we(alert_test_we),
		.wd(alert_test_wd),
		.d(sv2v_uu_u_alert_test_ext_d_0),
		.qre(),
		.qe(reg2hw[163]),
		.q(reg2hw[164]),
		.qs()
	);
	// Trace: design.sv:77131:3
	localparam signed [31:0] sv2v_uu_u_control_rx_watermark_DW = 8;
	// removed localparam type sv2v_uu_u_control_rx_watermark_d
	localparam [7:0] sv2v_uu_u_control_rx_watermark_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("RW"),
		.RESVAL(8'h7f)
	) u_control_rx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_rx_watermark_we),
		.wd(control_rx_watermark_wd),
		.de(1'b0),
		.d(sv2v_uu_u_control_rx_watermark_ext_d_0),
		.qe(),
		.q(reg2hw[162-:8]),
		.qs(control_rx_watermark_qs)
	);
	// Trace: design.sv:77157:3
	localparam signed [31:0] sv2v_uu_u_control_tx_watermark_DW = 8;
	// removed localparam type sv2v_uu_u_control_tx_watermark_d
	localparam [7:0] sv2v_uu_u_control_tx_watermark_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("RW"),
		.RESVAL(8'h00)
	) u_control_tx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_tx_watermark_we),
		.wd(control_tx_watermark_wd),
		.de(1'b0),
		.d(sv2v_uu_u_control_tx_watermark_ext_d_0),
		.qe(),
		.q(reg2hw[154-:8]),
		.qs(control_tx_watermark_qs)
	);
	// Trace: design.sv:77183:3
	localparam signed [31:0] sv2v_uu_u_control_output_en_DW = 1;
	// removed localparam type sv2v_uu_u_control_output_en_d
	localparam [0:0] sv2v_uu_u_control_output_en_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_control_output_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_output_en_we),
		.wd(control_output_en_wd),
		.de(1'b0),
		.d(sv2v_uu_u_control_output_en_ext_d_0),
		.qe(),
		.q(reg2hw[146]),
		.qs(control_output_en_qs)
	);
	// Trace: design.sv:77209:3
	localparam signed [31:0] sv2v_uu_u_control_sw_rst_DW = 1;
	// removed localparam type sv2v_uu_u_control_sw_rst_d
	localparam [0:0] sv2v_uu_u_control_sw_rst_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_control_sw_rst(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_sw_rst_we),
		.wd(control_sw_rst_wd),
		.de(1'b0),
		.d(sv2v_uu_u_control_sw_rst_ext_d_0),
		.qe(),
		.q(reg2hw[145]),
		.qs(control_sw_rst_qs)
	);
	// Trace: design.sv:77235:3
	localparam signed [31:0] sv2v_uu_u_control_spien_DW = 1;
	// removed localparam type sv2v_uu_u_control_spien_d
	localparam [0:0] sv2v_uu_u_control_spien_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_control_spien(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_spien_we),
		.wd(control_spien_wd),
		.de(1'b0),
		.d(sv2v_uu_u_control_spien_ext_d_0),
		.qe(),
		.q(reg2hw[144]),
		.qs(control_spien_qs)
	);
	// Trace: design.sv:77263:3
	localparam signed [31:0] sv2v_uu_u_status_txqd_DW = 8;
	// removed localparam type sv2v_uu_u_status_txqd_wd
	localparam [7:0] sv2v_uu_u_status_txqd_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("RO"),
		.RESVAL(8'h00)
	) u_status_txqd(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txqd_ext_wd_0),
		.de(hw2reg[48]),
		.d(hw2reg[56-:8]),
		.qe(),
		.q(),
		.qs(status_txqd_qs)
	);
	// Trace: design.sv:77288:3
	localparam signed [31:0] sv2v_uu_u_status_rxqd_DW = 8;
	// removed localparam type sv2v_uu_u_status_rxqd_wd
	localparam [7:0] sv2v_uu_u_status_rxqd_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("RO"),
		.RESVAL(8'h00)
	) u_status_rxqd(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxqd_ext_wd_0),
		.de(hw2reg[39]),
		.d(hw2reg[47-:8]),
		.qe(),
		.q(),
		.qs(status_rxqd_qs)
	);
	// Trace: design.sv:77313:3
	localparam signed [31:0] sv2v_uu_u_status_cmdqd_DW = 4;
	// removed localparam type sv2v_uu_u_status_cmdqd_wd
	localparam [3:0] sv2v_uu_u_status_cmdqd_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(4),
		.SWACCESS("RO"),
		.RESVAL(4'h0)
	) u_status_cmdqd(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_cmdqd_ext_wd_0),
		.de(hw2reg[34]),
		.d(hw2reg[38-:4]),
		.qe(),
		.q(),
		.qs(status_cmdqd_qs)
	);
	// Trace: design.sv:77338:3
	localparam signed [31:0] sv2v_uu_u_status_rxwm_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxwm_wd
	localparam [0:0] sv2v_uu_u_status_rxwm_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_rxwm(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxwm_ext_wd_0),
		.de(hw2reg[32]),
		.d(hw2reg[33]),
		.qe(),
		.q(),
		.qs(status_rxwm_qs)
	);
	// Trace: design.sv:77363:3
	localparam signed [31:0] sv2v_uu_u_status_byteorder_DW = 1;
	// removed localparam type sv2v_uu_u_status_byteorder_wd
	localparam [0:0] sv2v_uu_u_status_byteorder_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_byteorder(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_byteorder_ext_wd_0),
		.de(hw2reg[30]),
		.d(hw2reg[31]),
		.qe(),
		.q(),
		.qs(status_byteorder_qs)
	);
	// Trace: design.sv:77388:3
	localparam signed [31:0] sv2v_uu_u_status_rxstall_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxstall_wd
	localparam [0:0] sv2v_uu_u_status_rxstall_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_rxstall(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxstall_ext_wd_0),
		.de(hw2reg[28]),
		.d(hw2reg[29]),
		.qe(),
		.q(),
		.qs(status_rxstall_qs)
	);
	// Trace: design.sv:77413:3
	localparam signed [31:0] sv2v_uu_u_status_rxempty_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxempty_wd
	localparam [0:0] sv2v_uu_u_status_rxempty_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_rxempty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxempty_ext_wd_0),
		.de(hw2reg[26]),
		.d(hw2reg[27]),
		.qe(),
		.q(),
		.qs(status_rxempty_qs)
	);
	// Trace: design.sv:77438:3
	localparam signed [31:0] sv2v_uu_u_status_rxfull_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxfull_wd
	localparam [0:0] sv2v_uu_u_status_rxfull_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_rxfull(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxfull_ext_wd_0),
		.de(hw2reg[24]),
		.d(hw2reg[25]),
		.qe(),
		.q(),
		.qs(status_rxfull_qs)
	);
	// Trace: design.sv:77463:3
	localparam signed [31:0] sv2v_uu_u_status_txwm_DW = 1;
	// removed localparam type sv2v_uu_u_status_txwm_wd
	localparam [0:0] sv2v_uu_u_status_txwm_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_txwm(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txwm_ext_wd_0),
		.de(hw2reg[22]),
		.d(hw2reg[23]),
		.qe(),
		.q(),
		.qs(status_txwm_qs)
	);
	// Trace: design.sv:77488:3
	localparam signed [31:0] sv2v_uu_u_status_txstall_DW = 1;
	// removed localparam type sv2v_uu_u_status_txstall_wd
	localparam [0:0] sv2v_uu_u_status_txstall_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_txstall(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txstall_ext_wd_0),
		.de(hw2reg[20]),
		.d(hw2reg[21]),
		.qe(),
		.q(),
		.qs(status_txstall_qs)
	);
	// Trace: design.sv:77513:3
	localparam signed [31:0] sv2v_uu_u_status_txempty_DW = 1;
	// removed localparam type sv2v_uu_u_status_txempty_wd
	localparam [0:0] sv2v_uu_u_status_txempty_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_txempty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txempty_ext_wd_0),
		.de(hw2reg[18]),
		.d(hw2reg[19]),
		.qe(),
		.q(),
		.qs(status_txempty_qs)
	);
	// Trace: design.sv:77538:3
	localparam signed [31:0] sv2v_uu_u_status_txfull_DW = 1;
	// removed localparam type sv2v_uu_u_status_txfull_wd
	localparam [0:0] sv2v_uu_u_status_txfull_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_txfull(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txfull_ext_wd_0),
		.de(hw2reg[16]),
		.d(hw2reg[17]),
		.qe(),
		.q(),
		.qs(status_txfull_qs)
	);
	// Trace: design.sv:77563:3
	localparam signed [31:0] sv2v_uu_u_status_active_DW = 1;
	// removed localparam type sv2v_uu_u_status_active_wd
	localparam [0:0] sv2v_uu_u_status_active_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_active(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_active_ext_wd_0),
		.de(hw2reg[14]),
		.d(hw2reg[15]),
		.qe(),
		.q(),
		.qs(status_active_qs)
	);
	// Trace: design.sv:77588:3
	localparam signed [31:0] sv2v_uu_u_status_ready_DW = 1;
	// removed localparam type sv2v_uu_u_status_ready_wd
	localparam [0:0] sv2v_uu_u_status_ready_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_status_ready(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_status_ready_ext_wd_0),
		.de(hw2reg[12]),
		.d(hw2reg[13]),
		.qe(),
		.q(),
		.qs(status_ready_qs)
	);
	// Trace: design.sv:77617:3
	localparam signed [31:0] sv2v_uu_u_configopts_0_clkdiv_0_DW = 16;
	// removed localparam type sv2v_uu_u_configopts_0_clkdiv_0_d
	localparam [15:0] sv2v_uu_u_configopts_0_clkdiv_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_configopts_0_clkdiv_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_0_clkdiv_0_we),
		.wd(configopts_0_clkdiv_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_0_clkdiv_0_ext_d_0),
		.qe(),
		.q(reg2hw[112-:16]),
		.qs(configopts_0_clkdiv_0_qs)
	);
	// Trace: design.sv:77643:3
	localparam signed [31:0] sv2v_uu_u_configopts_0_csnidle_0_DW = 4;
	// removed localparam type sv2v_uu_u_configopts_0_csnidle_0_d
	localparam [3:0] sv2v_uu_u_configopts_0_csnidle_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(4),
		.SWACCESS("RW"),
		.RESVAL(4'h0)
	) u_configopts_0_csnidle_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_0_csnidle_0_we),
		.wd(configopts_0_csnidle_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_0_csnidle_0_ext_d_0),
		.qe(),
		.q(reg2hw[96-:4]),
		.qs(configopts_0_csnidle_0_qs)
	);
	// Trace: design.sv:77669:3
	localparam signed [31:0] sv2v_uu_u_configopts_0_csntrail_0_DW = 4;
	// removed localparam type sv2v_uu_u_configopts_0_csntrail_0_d
	localparam [3:0] sv2v_uu_u_configopts_0_csntrail_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(4),
		.SWACCESS("RW"),
		.RESVAL(4'h0)
	) u_configopts_0_csntrail_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_0_csntrail_0_we),
		.wd(configopts_0_csntrail_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_0_csntrail_0_ext_d_0),
		.qe(),
		.q(reg2hw[92-:4]),
		.qs(configopts_0_csntrail_0_qs)
	);
	// Trace: design.sv:77695:3
	localparam signed [31:0] sv2v_uu_u_configopts_0_csnlead_0_DW = 4;
	// removed localparam type sv2v_uu_u_configopts_0_csnlead_0_d
	localparam [3:0] sv2v_uu_u_configopts_0_csnlead_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(4),
		.SWACCESS("RW"),
		.RESVAL(4'h0)
	) u_configopts_0_csnlead_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_0_csnlead_0_we),
		.wd(configopts_0_csnlead_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_0_csnlead_0_ext_d_0),
		.qe(),
		.q(reg2hw[88-:4]),
		.qs(configopts_0_csnlead_0_qs)
	);
	// Trace: design.sv:77721:3
	localparam signed [31:0] sv2v_uu_u_configopts_0_fullcyc_0_DW = 1;
	// removed localparam type sv2v_uu_u_configopts_0_fullcyc_0_d
	localparam [0:0] sv2v_uu_u_configopts_0_fullcyc_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_configopts_0_fullcyc_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_0_fullcyc_0_we),
		.wd(configopts_0_fullcyc_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_0_fullcyc_0_ext_d_0),
		.qe(),
		.q(reg2hw[84]),
		.qs(configopts_0_fullcyc_0_qs)
	);
	// Trace: design.sv:77747:3
	localparam signed [31:0] sv2v_uu_u_configopts_0_cpha_0_DW = 1;
	// removed localparam type sv2v_uu_u_configopts_0_cpha_0_d
	localparam [0:0] sv2v_uu_u_configopts_0_cpha_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_configopts_0_cpha_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_0_cpha_0_we),
		.wd(configopts_0_cpha_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_0_cpha_0_ext_d_0),
		.qe(),
		.q(reg2hw[83]),
		.qs(configopts_0_cpha_0_qs)
	);
	// Trace: design.sv:77773:3
	localparam signed [31:0] sv2v_uu_u_configopts_0_cpol_0_DW = 1;
	// removed localparam type sv2v_uu_u_configopts_0_cpol_0_d
	localparam [0:0] sv2v_uu_u_configopts_0_cpol_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_configopts_0_cpol_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_0_cpol_0_we),
		.wd(configopts_0_cpol_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_0_cpol_0_ext_d_0),
		.qe(),
		.q(reg2hw[82]),
		.qs(configopts_0_cpol_0_qs)
	);
	// Trace: design.sv:77802:3
	localparam signed [31:0] sv2v_uu_u_configopts_1_clkdiv_1_DW = 16;
	// removed localparam type sv2v_uu_u_configopts_1_clkdiv_1_d
	localparam [15:0] sv2v_uu_u_configopts_1_clkdiv_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_configopts_1_clkdiv_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_1_clkdiv_1_we),
		.wd(configopts_1_clkdiv_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_1_clkdiv_1_ext_d_0),
		.qe(),
		.q(reg2hw[143-:16]),
		.qs(configopts_1_clkdiv_1_qs)
	);
	// Trace: design.sv:77828:3
	localparam signed [31:0] sv2v_uu_u_configopts_1_csnidle_1_DW = 4;
	// removed localparam type sv2v_uu_u_configopts_1_csnidle_1_d
	localparam [3:0] sv2v_uu_u_configopts_1_csnidle_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(4),
		.SWACCESS("RW"),
		.RESVAL(4'h0)
	) u_configopts_1_csnidle_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_1_csnidle_1_we),
		.wd(configopts_1_csnidle_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_1_csnidle_1_ext_d_0),
		.qe(),
		.q(reg2hw[127-:4]),
		.qs(configopts_1_csnidle_1_qs)
	);
	// Trace: design.sv:77854:3
	localparam signed [31:0] sv2v_uu_u_configopts_1_csntrail_1_DW = 4;
	// removed localparam type sv2v_uu_u_configopts_1_csntrail_1_d
	localparam [3:0] sv2v_uu_u_configopts_1_csntrail_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(4),
		.SWACCESS("RW"),
		.RESVAL(4'h0)
	) u_configopts_1_csntrail_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_1_csntrail_1_we),
		.wd(configopts_1_csntrail_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_1_csntrail_1_ext_d_0),
		.qe(),
		.q(reg2hw[123-:4]),
		.qs(configopts_1_csntrail_1_qs)
	);
	// Trace: design.sv:77880:3
	localparam signed [31:0] sv2v_uu_u_configopts_1_csnlead_1_DW = 4;
	// removed localparam type sv2v_uu_u_configopts_1_csnlead_1_d
	localparam [3:0] sv2v_uu_u_configopts_1_csnlead_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(4),
		.SWACCESS("RW"),
		.RESVAL(4'h0)
	) u_configopts_1_csnlead_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_1_csnlead_1_we),
		.wd(configopts_1_csnlead_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_1_csnlead_1_ext_d_0),
		.qe(),
		.q(reg2hw[119-:4]),
		.qs(configopts_1_csnlead_1_qs)
	);
	// Trace: design.sv:77906:3
	localparam signed [31:0] sv2v_uu_u_configopts_1_fullcyc_1_DW = 1;
	// removed localparam type sv2v_uu_u_configopts_1_fullcyc_1_d
	localparam [0:0] sv2v_uu_u_configopts_1_fullcyc_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_configopts_1_fullcyc_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_1_fullcyc_1_we),
		.wd(configopts_1_fullcyc_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_1_fullcyc_1_ext_d_0),
		.qe(),
		.q(reg2hw[115]),
		.qs(configopts_1_fullcyc_1_qs)
	);
	// Trace: design.sv:77932:3
	localparam signed [31:0] sv2v_uu_u_configopts_1_cpha_1_DW = 1;
	// removed localparam type sv2v_uu_u_configopts_1_cpha_1_d
	localparam [0:0] sv2v_uu_u_configopts_1_cpha_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_configopts_1_cpha_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_1_cpha_1_we),
		.wd(configopts_1_cpha_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_1_cpha_1_ext_d_0),
		.qe(),
		.q(reg2hw[114]),
		.qs(configopts_1_cpha_1_qs)
	);
	// Trace: design.sv:77958:3
	localparam signed [31:0] sv2v_uu_u_configopts_1_cpol_1_DW = 1;
	// removed localparam type sv2v_uu_u_configopts_1_cpol_1_d
	localparam [0:0] sv2v_uu_u_configopts_1_cpol_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_configopts_1_cpol_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(configopts_1_cpol_1_we),
		.wd(configopts_1_cpol_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_configopts_1_cpol_1_ext_d_0),
		.qe(),
		.q(reg2hw[113]),
		.qs(configopts_1_cpol_1_qs)
	);
	// Trace: design.sv:77986:3
	localparam signed [31:0] sv2v_uu_u_csid_DW = 32;
	// removed localparam type sv2v_uu_u_csid_d
	localparam [31:0] sv2v_uu_u_csid_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_csid(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(csid_we),
		.wd(csid_wd),
		.de(1'b0),
		.d(sv2v_uu_u_csid_ext_d_0),
		.qe(),
		.q(reg2hw[81-:32]),
		.qs(csid_qs)
	);
	// Trace: design.sv:78014:3
	localparam [31:0] sv2v_uu_u_command_len_DW = 24;
	// removed localparam type sv2v_uu_u_command_len_d
	localparam [23:0] sv2v_uu_u_command_len_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(24)) u_command_len(
		.re(1'b0),
		.we(command_len_we),
		.wd(command_len_wd),
		.d(sv2v_uu_u_command_len_ext_d_0),
		.qre(),
		.qe(reg2hw[25]),
		.q(reg2hw[49-:24]),
		.qs()
	);
	// Trace: design.sv:78029:3
	localparam [31:0] sv2v_uu_u_command_csaat_DW = 1;
	// removed localparam type sv2v_uu_u_command_csaat_d
	localparam [0:0] sv2v_uu_u_command_csaat_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_command_csaat(
		.re(1'b0),
		.we(command_csaat_we),
		.wd(command_csaat_wd),
		.d(sv2v_uu_u_command_csaat_ext_d_0),
		.qre(),
		.qe(reg2hw[23]),
		.q(reg2hw[24]),
		.qs()
	);
	// Trace: design.sv:78044:3
	localparam [31:0] sv2v_uu_u_command_speed_DW = 2;
	// removed localparam type sv2v_uu_u_command_speed_d
	localparam [1:0] sv2v_uu_u_command_speed_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(2)) u_command_speed(
		.re(1'b0),
		.we(command_speed_we),
		.wd(command_speed_wd),
		.d(sv2v_uu_u_command_speed_ext_d_0),
		.qre(),
		.qe(reg2hw[20]),
		.q(reg2hw[22-:2]),
		.qs()
	);
	// Trace: design.sv:78059:3
	localparam [31:0] sv2v_uu_u_command_direction_DW = 2;
	// removed localparam type sv2v_uu_u_command_direction_d
	localparam [1:0] sv2v_uu_u_command_direction_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(2)) u_command_direction(
		.re(1'b0),
		.we(command_direction_we),
		.wd(command_direction_wd),
		.d(sv2v_uu_u_command_direction_ext_d_0),
		.qre(),
		.qe(reg2hw[17]),
		.q(reg2hw[19-:2]),
		.qs()
	);
	// Trace: design.sv:78076:3
	localparam signed [31:0] sv2v_uu_u_error_enable_cmdbusy_DW = 1;
	// removed localparam type sv2v_uu_u_error_enable_cmdbusy_d
	localparam [0:0] sv2v_uu_u_error_enable_cmdbusy_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h1)
	) u_error_enable_cmdbusy(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_enable_cmdbusy_we),
		.wd(error_enable_cmdbusy_wd),
		.de(1'b0),
		.d(sv2v_uu_u_error_enable_cmdbusy_ext_d_0),
		.qe(),
		.q(reg2hw[16]),
		.qs(error_enable_cmdbusy_qs)
	);
	// Trace: design.sv:78102:3
	localparam signed [31:0] sv2v_uu_u_error_enable_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_error_enable_overflow_d
	localparam [0:0] sv2v_uu_u_error_enable_overflow_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h1)
	) u_error_enable_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_enable_overflow_we),
		.wd(error_enable_overflow_wd),
		.de(1'b0),
		.d(sv2v_uu_u_error_enable_overflow_ext_d_0),
		.qe(),
		.q(reg2hw[15]),
		.qs(error_enable_overflow_qs)
	);
	// Trace: design.sv:78128:3
	localparam signed [31:0] sv2v_uu_u_error_enable_underflow_DW = 1;
	// removed localparam type sv2v_uu_u_error_enable_underflow_d
	localparam [0:0] sv2v_uu_u_error_enable_underflow_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h1)
	) u_error_enable_underflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_enable_underflow_we),
		.wd(error_enable_underflow_wd),
		.de(1'b0),
		.d(sv2v_uu_u_error_enable_underflow_ext_d_0),
		.qe(),
		.q(reg2hw[14]),
		.qs(error_enable_underflow_qs)
	);
	// Trace: design.sv:78154:3
	localparam signed [31:0] sv2v_uu_u_error_enable_cmdinval_DW = 1;
	// removed localparam type sv2v_uu_u_error_enable_cmdinval_d
	localparam [0:0] sv2v_uu_u_error_enable_cmdinval_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h1)
	) u_error_enable_cmdinval(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_enable_cmdinval_we),
		.wd(error_enable_cmdinval_wd),
		.de(1'b0),
		.d(sv2v_uu_u_error_enable_cmdinval_ext_d_0),
		.qe(),
		.q(reg2hw[13]),
		.qs(error_enable_cmdinval_qs)
	);
	// Trace: design.sv:78180:3
	localparam signed [31:0] sv2v_uu_u_error_enable_csidinval_DW = 1;
	// removed localparam type sv2v_uu_u_error_enable_csidinval_d
	localparam [0:0] sv2v_uu_u_error_enable_csidinval_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h1)
	) u_error_enable_csidinval(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_enable_csidinval_we),
		.wd(error_enable_csidinval_wd),
		.de(1'b0),
		.d(sv2v_uu_u_error_enable_csidinval_ext_d_0),
		.qe(),
		.q(reg2hw[12]),
		.qs(error_enable_csidinval_qs)
	);
	// Trace: design.sv:78208:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_error_status_cmdbusy(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_status_cmdbusy_we),
		.wd(error_status_cmdbusy_wd),
		.de(hw2reg[10]),
		.d(hw2reg[11]),
		.qe(),
		.q(reg2hw[11]),
		.qs(error_status_cmdbusy_qs)
	);
	// Trace: design.sv:78234:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_error_status_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_status_overflow_we),
		.wd(error_status_overflow_wd),
		.de(hw2reg[8]),
		.d(hw2reg[9]),
		.qe(),
		.q(reg2hw[10]),
		.qs(error_status_overflow_qs)
	);
	// Trace: design.sv:78260:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_error_status_underflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_status_underflow_we),
		.wd(error_status_underflow_wd),
		.de(hw2reg[6]),
		.d(hw2reg[7]),
		.qe(),
		.q(reg2hw[9]),
		.qs(error_status_underflow_qs)
	);
	// Trace: design.sv:78286:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_error_status_cmdinval(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_status_cmdinval_we),
		.wd(error_status_cmdinval_wd),
		.de(hw2reg[4]),
		.d(hw2reg[5]),
		.qe(),
		.q(reg2hw[8]),
		.qs(error_status_cmdinval_qs)
	);
	// Trace: design.sv:78312:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_error_status_csidinval(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_status_csidinval_we),
		.wd(error_status_csidinval_wd),
		.de(hw2reg[2]),
		.d(hw2reg[3]),
		.qe(),
		.q(reg2hw[7]),
		.qs(error_status_csidinval_qs)
	);
	// Trace: design.sv:78338:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_error_status_accessinval(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(error_status_accessinval_we),
		.wd(error_status_accessinval_wd),
		.de(hw2reg[0]),
		.d(hw2reg[1]),
		.qe(),
		.q(reg2hw[6]),
		.qs(error_status_accessinval_qs)
	);
	// Trace: design.sv:78366:3
	localparam signed [31:0] sv2v_uu_u_event_enable_rxfull_DW = 1;
	// removed localparam type sv2v_uu_u_event_enable_rxfull_d
	localparam [0:0] sv2v_uu_u_event_enable_rxfull_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_event_enable_rxfull(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(event_enable_rxfull_we),
		.wd(event_enable_rxfull_wd),
		.de(1'b0),
		.d(sv2v_uu_u_event_enable_rxfull_ext_d_0),
		.qe(),
		.q(reg2hw[5]),
		.qs(event_enable_rxfull_qs)
	);
	// Trace: design.sv:78392:3
	localparam signed [31:0] sv2v_uu_u_event_enable_txempty_DW = 1;
	// removed localparam type sv2v_uu_u_event_enable_txempty_d
	localparam [0:0] sv2v_uu_u_event_enable_txempty_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_event_enable_txempty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(event_enable_txempty_we),
		.wd(event_enable_txempty_wd),
		.de(1'b0),
		.d(sv2v_uu_u_event_enable_txempty_ext_d_0),
		.qe(),
		.q(reg2hw[4]),
		.qs(event_enable_txempty_qs)
	);
	// Trace: design.sv:78418:3
	localparam signed [31:0] sv2v_uu_u_event_enable_rxwm_DW = 1;
	// removed localparam type sv2v_uu_u_event_enable_rxwm_d
	localparam [0:0] sv2v_uu_u_event_enable_rxwm_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_event_enable_rxwm(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(event_enable_rxwm_we),
		.wd(event_enable_rxwm_wd),
		.de(1'b0),
		.d(sv2v_uu_u_event_enable_rxwm_ext_d_0),
		.qe(),
		.q(reg2hw[3]),
		.qs(event_enable_rxwm_qs)
	);
	// Trace: design.sv:78444:3
	localparam signed [31:0] sv2v_uu_u_event_enable_txwm_DW = 1;
	// removed localparam type sv2v_uu_u_event_enable_txwm_d
	localparam [0:0] sv2v_uu_u_event_enable_txwm_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_event_enable_txwm(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(event_enable_txwm_we),
		.wd(event_enable_txwm_wd),
		.de(1'b0),
		.d(sv2v_uu_u_event_enable_txwm_ext_d_0),
		.qe(),
		.q(reg2hw[2]),
		.qs(event_enable_txwm_qs)
	);
	// Trace: design.sv:78470:3
	localparam signed [31:0] sv2v_uu_u_event_enable_ready_DW = 1;
	// removed localparam type sv2v_uu_u_event_enable_ready_d
	localparam [0:0] sv2v_uu_u_event_enable_ready_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_event_enable_ready(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(event_enable_ready_we),
		.wd(event_enable_ready_wd),
		.de(1'b0),
		.d(sv2v_uu_u_event_enable_ready_ext_d_0),
		.qe(),
		.q(reg2hw[1]),
		.qs(event_enable_ready_qs)
	);
	// Trace: design.sv:78496:3
	localparam signed [31:0] sv2v_uu_u_event_enable_idle_DW = 1;
	// removed localparam type sv2v_uu_u_event_enable_idle_d
	localparam [0:0] sv2v_uu_u_event_enable_idle_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_event_enable_idle(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(event_enable_idle_we),
		.wd(event_enable_idle_wd),
		.de(1'b0),
		.d(sv2v_uu_u_event_enable_idle_ext_d_0),
		.qe(),
		.q(reg2hw[0]),
		.qs(event_enable_idle_qs)
	);
	// Trace: design.sv:78523:3
	reg [12:0] addr_hit;
	// Trace: design.sv:78524:3
	localparam signed [31:0] spi_host_reg_pkg_BlockAw = 6;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_ALERT_TEST_OFFSET = 6'h0c;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_COMMAND_OFFSET = 6'h24;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_CONFIGOPTS_0_OFFSET = 6'h18;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_CONFIGOPTS_1_OFFSET = 6'h1c;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_CONTROL_OFFSET = 6'h10;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_CSID_OFFSET = 6'h20;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_ERROR_ENABLE_OFFSET = 6'h30;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_ERROR_STATUS_OFFSET = 6'h34;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_EVENT_ENABLE_OFFSET = 6'h38;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_INTR_ENABLE_OFFSET = 6'h04;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_INTR_STATE_OFFSET = 6'h00;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_INTR_TEST_OFFSET = 6'h08;
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_STATUS_OFFSET = 6'h14;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:78525:5
		addr_hit = 1'sb0;
		// Trace: design.sv:78526:5
		addr_hit[0] = reg_addr == spi_host_reg_pkg_SPI_HOST_INTR_STATE_OFFSET;
		// Trace: design.sv:78527:5
		addr_hit[1] = reg_addr == spi_host_reg_pkg_SPI_HOST_INTR_ENABLE_OFFSET;
		// Trace: design.sv:78528:5
		addr_hit[2] = reg_addr == spi_host_reg_pkg_SPI_HOST_INTR_TEST_OFFSET;
		// Trace: design.sv:78529:5
		addr_hit[3] = reg_addr == spi_host_reg_pkg_SPI_HOST_ALERT_TEST_OFFSET;
		// Trace: design.sv:78530:5
		addr_hit[4] = reg_addr == spi_host_reg_pkg_SPI_HOST_CONTROL_OFFSET;
		// Trace: design.sv:78531:5
		addr_hit[5] = reg_addr == spi_host_reg_pkg_SPI_HOST_STATUS_OFFSET;
		// Trace: design.sv:78532:5
		addr_hit[6] = reg_addr == spi_host_reg_pkg_SPI_HOST_CONFIGOPTS_0_OFFSET;
		// Trace: design.sv:78533:5
		addr_hit[7] = reg_addr == spi_host_reg_pkg_SPI_HOST_CONFIGOPTS_1_OFFSET;
		// Trace: design.sv:78534:5
		addr_hit[8] = reg_addr == spi_host_reg_pkg_SPI_HOST_CSID_OFFSET;
		// Trace: design.sv:78535:5
		addr_hit[9] = reg_addr == spi_host_reg_pkg_SPI_HOST_COMMAND_OFFSET;
		// Trace: design.sv:78536:5
		addr_hit[10] = reg_addr == spi_host_reg_pkg_SPI_HOST_ERROR_ENABLE_OFFSET;
		// Trace: design.sv:78537:5
		addr_hit[11] = reg_addr == spi_host_reg_pkg_SPI_HOST_ERROR_STATUS_OFFSET;
		// Trace: design.sv:78538:5
		addr_hit[12] = reg_addr == spi_host_reg_pkg_SPI_HOST_EVENT_ENABLE_OFFSET;
	end
	// Trace: design.sv:78541:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:78544:3
	localparam [51:0] spi_host_reg_pkg_SPI_HOST_PERMIT = 52'b0001000100010001111111111111111111111111000100010001;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:78545:5
		wr_err = reg_we & (((((((((((((addr_hit[0] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[48+:4] & ~reg_be)) | (addr_hit[1] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[44+:4] & ~reg_be))) | (addr_hit[2] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[40+:4] & ~reg_be))) | (addr_hit[3] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[36+:4] & ~reg_be))) | (addr_hit[4] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[32+:4] & ~reg_be))) | (addr_hit[5] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[28+:4] & ~reg_be))) | (addr_hit[6] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[24+:4] & ~reg_be))) | (addr_hit[7] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[20+:4] & ~reg_be))) | (addr_hit[8] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[16+:4] & ~reg_be))) | (addr_hit[9] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[12+:4] & ~reg_be))) | (addr_hit[10] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[8+:4] & ~reg_be))) | (addr_hit[11] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[4+:4] & ~reg_be))) | (addr_hit[12] & |(spi_host_reg_pkg_SPI_HOST_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:78561:3
	assign intr_state_error_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:78562:3
	assign intr_state_error_wd = reg_wdata[0];
	// Trace: design.sv:78564:3
	assign intr_state_spi_event_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:78565:3
	assign intr_state_spi_event_wd = reg_wdata[1];
	// Trace: design.sv:78567:3
	assign intr_enable_error_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:78568:3
	assign intr_enable_error_wd = reg_wdata[0];
	// Trace: design.sv:78570:3
	assign intr_enable_spi_event_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:78571:3
	assign intr_enable_spi_event_wd = reg_wdata[1];
	// Trace: design.sv:78573:3
	assign intr_test_error_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:78574:3
	assign intr_test_error_wd = reg_wdata[0];
	// Trace: design.sv:78576:3
	assign intr_test_spi_event_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:78577:3
	assign intr_test_spi_event_wd = reg_wdata[1];
	// Trace: design.sv:78579:3
	assign alert_test_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:78580:3
	assign alert_test_wd = reg_wdata[0];
	// Trace: design.sv:78582:3
	assign control_rx_watermark_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:78583:3
	assign control_rx_watermark_wd = reg_wdata[7:0];
	// Trace: design.sv:78585:3
	assign control_tx_watermark_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:78586:3
	assign control_tx_watermark_wd = reg_wdata[15:8];
	// Trace: design.sv:78588:3
	assign control_output_en_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:78589:3
	assign control_output_en_wd = reg_wdata[29];
	// Trace: design.sv:78591:3
	assign control_sw_rst_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:78592:3
	assign control_sw_rst_wd = reg_wdata[30];
	// Trace: design.sv:78594:3
	assign control_spien_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:78595:3
	assign control_spien_wd = reg_wdata[31];
	// Trace: design.sv:78597:3
	assign configopts_0_clkdiv_0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:78598:3
	assign configopts_0_clkdiv_0_wd = reg_wdata[15:0];
	// Trace: design.sv:78600:3
	assign configopts_0_csnidle_0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:78601:3
	assign configopts_0_csnidle_0_wd = reg_wdata[19:16];
	// Trace: design.sv:78603:3
	assign configopts_0_csntrail_0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:78604:3
	assign configopts_0_csntrail_0_wd = reg_wdata[23:20];
	// Trace: design.sv:78606:3
	assign configopts_0_csnlead_0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:78607:3
	assign configopts_0_csnlead_0_wd = reg_wdata[27:24];
	// Trace: design.sv:78609:3
	assign configopts_0_fullcyc_0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:78610:3
	assign configopts_0_fullcyc_0_wd = reg_wdata[29];
	// Trace: design.sv:78612:3
	assign configopts_0_cpha_0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:78613:3
	assign configopts_0_cpha_0_wd = reg_wdata[30];
	// Trace: design.sv:78615:3
	assign configopts_0_cpol_0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:78616:3
	assign configopts_0_cpol_0_wd = reg_wdata[31];
	// Trace: design.sv:78618:3
	assign configopts_1_clkdiv_1_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:78619:3
	assign configopts_1_clkdiv_1_wd = reg_wdata[15:0];
	// Trace: design.sv:78621:3
	assign configopts_1_csnidle_1_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:78622:3
	assign configopts_1_csnidle_1_wd = reg_wdata[19:16];
	// Trace: design.sv:78624:3
	assign configopts_1_csntrail_1_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:78625:3
	assign configopts_1_csntrail_1_wd = reg_wdata[23:20];
	// Trace: design.sv:78627:3
	assign configopts_1_csnlead_1_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:78628:3
	assign configopts_1_csnlead_1_wd = reg_wdata[27:24];
	// Trace: design.sv:78630:3
	assign configopts_1_fullcyc_1_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:78631:3
	assign configopts_1_fullcyc_1_wd = reg_wdata[29];
	// Trace: design.sv:78633:3
	assign configopts_1_cpha_1_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:78634:3
	assign configopts_1_cpha_1_wd = reg_wdata[30];
	// Trace: design.sv:78636:3
	assign configopts_1_cpol_1_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:78637:3
	assign configopts_1_cpol_1_wd = reg_wdata[31];
	// Trace: design.sv:78639:3
	assign csid_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:78640:3
	assign csid_wd = reg_wdata[31:0];
	// Trace: design.sv:78642:3
	assign command_len_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:78643:3
	assign command_len_wd = reg_wdata[23:0];
	// Trace: design.sv:78645:3
	assign command_csaat_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:78646:3
	assign command_csaat_wd = reg_wdata[24];
	// Trace: design.sv:78648:3
	assign command_speed_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:78649:3
	assign command_speed_wd = reg_wdata[26:25];
	// Trace: design.sv:78651:3
	assign command_direction_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:78652:3
	assign command_direction_wd = reg_wdata[28:27];
	// Trace: design.sv:78654:3
	assign error_enable_cmdbusy_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:78655:3
	assign error_enable_cmdbusy_wd = reg_wdata[0];
	// Trace: design.sv:78657:3
	assign error_enable_overflow_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:78658:3
	assign error_enable_overflow_wd = reg_wdata[1];
	// Trace: design.sv:78660:3
	assign error_enable_underflow_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:78661:3
	assign error_enable_underflow_wd = reg_wdata[2];
	// Trace: design.sv:78663:3
	assign error_enable_cmdinval_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:78664:3
	assign error_enable_cmdinval_wd = reg_wdata[3];
	// Trace: design.sv:78666:3
	assign error_enable_csidinval_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:78667:3
	assign error_enable_csidinval_wd = reg_wdata[4];
	// Trace: design.sv:78669:3
	assign error_status_cmdbusy_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:78670:3
	assign error_status_cmdbusy_wd = reg_wdata[0];
	// Trace: design.sv:78672:3
	assign error_status_overflow_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:78673:3
	assign error_status_overflow_wd = reg_wdata[1];
	// Trace: design.sv:78675:3
	assign error_status_underflow_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:78676:3
	assign error_status_underflow_wd = reg_wdata[2];
	// Trace: design.sv:78678:3
	assign error_status_cmdinval_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:78679:3
	assign error_status_cmdinval_wd = reg_wdata[3];
	// Trace: design.sv:78681:3
	assign error_status_csidinval_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:78682:3
	assign error_status_csidinval_wd = reg_wdata[4];
	// Trace: design.sv:78684:3
	assign error_status_accessinval_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:78685:3
	assign error_status_accessinval_wd = reg_wdata[5];
	// Trace: design.sv:78687:3
	assign event_enable_rxfull_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:78688:3
	assign event_enable_rxfull_wd = reg_wdata[0];
	// Trace: design.sv:78690:3
	assign event_enable_txempty_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:78691:3
	assign event_enable_txempty_wd = reg_wdata[1];
	// Trace: design.sv:78693:3
	assign event_enable_rxwm_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:78694:3
	assign event_enable_rxwm_wd = reg_wdata[2];
	// Trace: design.sv:78696:3
	assign event_enable_txwm_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:78697:3
	assign event_enable_txwm_wd = reg_wdata[3];
	// Trace: design.sv:78699:3
	assign event_enable_ready_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:78700:3
	assign event_enable_ready_wd = reg_wdata[4];
	// Trace: design.sv:78702:3
	assign event_enable_idle_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:78703:3
	assign event_enable_idle_wd = reg_wdata[5];
	// Trace: design.sv:78706:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:78707:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:78708:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]: begin
				// Trace: design.sv:78710:9
				reg_rdata_next[0] = intr_state_error_qs;
				// Trace: design.sv:78711:9
				reg_rdata_next[1] = intr_state_spi_event_qs;
			end
			addr_hit[1]: begin
				// Trace: design.sv:78715:9
				reg_rdata_next[0] = intr_enable_error_qs;
				// Trace: design.sv:78716:9
				reg_rdata_next[1] = intr_enable_spi_event_qs;
			end
			addr_hit[2]: begin
				// Trace: design.sv:78720:9
				reg_rdata_next[0] = 1'sb0;
				// Trace: design.sv:78721:9
				reg_rdata_next[1] = 1'sb0;
			end
			addr_hit[3]:
				// Trace: design.sv:78725:9
				reg_rdata_next[0] = 1'sb0;
			addr_hit[4]: begin
				// Trace: design.sv:78729:9
				reg_rdata_next[7:0] = control_rx_watermark_qs;
				// Trace: design.sv:78730:9
				reg_rdata_next[15:8] = control_tx_watermark_qs;
				// Trace: design.sv:78731:9
				reg_rdata_next[29] = control_output_en_qs;
				// Trace: design.sv:78732:9
				reg_rdata_next[30] = control_sw_rst_qs;
				// Trace: design.sv:78733:9
				reg_rdata_next[31] = control_spien_qs;
			end
			addr_hit[5]: begin
				// Trace: design.sv:78737:9
				reg_rdata_next[7:0] = status_txqd_qs;
				// Trace: design.sv:78738:9
				reg_rdata_next[15:8] = status_rxqd_qs;
				// Trace: design.sv:78739:9
				reg_rdata_next[19:16] = status_cmdqd_qs;
				// Trace: design.sv:78740:9
				reg_rdata_next[20] = status_rxwm_qs;
				// Trace: design.sv:78741:9
				reg_rdata_next[22] = status_byteorder_qs;
				// Trace: design.sv:78742:9
				reg_rdata_next[23] = status_rxstall_qs;
				// Trace: design.sv:78743:9
				reg_rdata_next[24] = status_rxempty_qs;
				// Trace: design.sv:78744:9
				reg_rdata_next[25] = status_rxfull_qs;
				// Trace: design.sv:78745:9
				reg_rdata_next[26] = status_txwm_qs;
				// Trace: design.sv:78746:9
				reg_rdata_next[27] = status_txstall_qs;
				// Trace: design.sv:78747:9
				reg_rdata_next[28] = status_txempty_qs;
				// Trace: design.sv:78748:9
				reg_rdata_next[29] = status_txfull_qs;
				// Trace: design.sv:78749:9
				reg_rdata_next[30] = status_active_qs;
				// Trace: design.sv:78750:9
				reg_rdata_next[31] = status_ready_qs;
			end
			addr_hit[6]: begin
				// Trace: design.sv:78754:9
				reg_rdata_next[15:0] = configopts_0_clkdiv_0_qs;
				// Trace: design.sv:78755:9
				reg_rdata_next[19:16] = configopts_0_csnidle_0_qs;
				// Trace: design.sv:78756:9
				reg_rdata_next[23:20] = configopts_0_csntrail_0_qs;
				// Trace: design.sv:78757:9
				reg_rdata_next[27:24] = configopts_0_csnlead_0_qs;
				// Trace: design.sv:78758:9
				reg_rdata_next[29] = configopts_0_fullcyc_0_qs;
				// Trace: design.sv:78759:9
				reg_rdata_next[30] = configopts_0_cpha_0_qs;
				// Trace: design.sv:78760:9
				reg_rdata_next[31] = configopts_0_cpol_0_qs;
			end
			addr_hit[7]: begin
				// Trace: design.sv:78764:9
				reg_rdata_next[15:0] = configopts_1_clkdiv_1_qs;
				// Trace: design.sv:78765:9
				reg_rdata_next[19:16] = configopts_1_csnidle_1_qs;
				// Trace: design.sv:78766:9
				reg_rdata_next[23:20] = configopts_1_csntrail_1_qs;
				// Trace: design.sv:78767:9
				reg_rdata_next[27:24] = configopts_1_csnlead_1_qs;
				// Trace: design.sv:78768:9
				reg_rdata_next[29] = configopts_1_fullcyc_1_qs;
				// Trace: design.sv:78769:9
				reg_rdata_next[30] = configopts_1_cpha_1_qs;
				// Trace: design.sv:78770:9
				reg_rdata_next[31] = configopts_1_cpol_1_qs;
			end
			addr_hit[8]:
				// Trace: design.sv:78774:9
				reg_rdata_next[31:0] = csid_qs;
			addr_hit[9]: begin
				// Trace: design.sv:78778:9
				reg_rdata_next[23:0] = 1'sb0;
				// Trace: design.sv:78779:9
				reg_rdata_next[24] = 1'sb0;
				// Trace: design.sv:78780:9
				reg_rdata_next[26:25] = 1'sb0;
				// Trace: design.sv:78781:9
				reg_rdata_next[28:27] = 1'sb0;
			end
			addr_hit[10]: begin
				// Trace: design.sv:78785:9
				reg_rdata_next[0] = error_enable_cmdbusy_qs;
				// Trace: design.sv:78786:9
				reg_rdata_next[1] = error_enable_overflow_qs;
				// Trace: design.sv:78787:9
				reg_rdata_next[2] = error_enable_underflow_qs;
				// Trace: design.sv:78788:9
				reg_rdata_next[3] = error_enable_cmdinval_qs;
				// Trace: design.sv:78789:9
				reg_rdata_next[4] = error_enable_csidinval_qs;
			end
			addr_hit[11]: begin
				// Trace: design.sv:78793:9
				reg_rdata_next[0] = error_status_cmdbusy_qs;
				// Trace: design.sv:78794:9
				reg_rdata_next[1] = error_status_overflow_qs;
				// Trace: design.sv:78795:9
				reg_rdata_next[2] = error_status_underflow_qs;
				// Trace: design.sv:78796:9
				reg_rdata_next[3] = error_status_cmdinval_qs;
				// Trace: design.sv:78797:9
				reg_rdata_next[4] = error_status_csidinval_qs;
				// Trace: design.sv:78798:9
				reg_rdata_next[5] = error_status_accessinval_qs;
			end
			addr_hit[12]: begin
				// Trace: design.sv:78802:9
				reg_rdata_next[0] = event_enable_rxfull_qs;
				// Trace: design.sv:78803:9
				reg_rdata_next[1] = event_enable_txempty_qs;
				// Trace: design.sv:78804:9
				reg_rdata_next[2] = event_enable_rxwm_qs;
				// Trace: design.sv:78805:9
				reg_rdata_next[3] = event_enable_txwm_qs;
				// Trace: design.sv:78806:9
				reg_rdata_next[4] = event_enable_ready_qs;
				// Trace: design.sv:78807:9
				reg_rdata_next[5] = event_enable_idle_qs;
			end
			default:
				// Trace: design.sv:78811:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:78820:3
	wire unused_wdata;
	// Trace: design.sv:78821:3
	wire unused_be;
	// Trace: design.sv:78822:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:78823:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module spi_host_window_9C1FC (
	clk_i,
	rst_ni,
	rx_win_i,
	rx_win_o,
	tx_win_i,
	tx_win_o,
	tx_data_o,
	tx_be_o,
	tx_valid_o,
	rx_data_i,
	rx_ready_o
);
	// Trace: design.sv:78840:18
	// removed localparam type reg_req_t
	// Trace: design.sv:78841:18
	// removed localparam type reg_rsp_t
	// Trace: design.sv:78843:3
	input clk_i;
	// Trace: design.sv:78844:3
	input rst_ni;
	// Trace: design.sv:78845:3
	input wire [69:0] rx_win_i;
	// Trace: design.sv:78846:3
	output wire [33:0] rx_win_o;
	// Trace: design.sv:78847:3
	input wire [69:0] tx_win_i;
	// Trace: design.sv:78848:3
	output wire [33:0] tx_win_o;
	// Trace: design.sv:78849:3
	output wire [31:0] tx_data_o;
	// Trace: design.sv:78850:3
	output wire [3:0] tx_be_o;
	// Trace: design.sv:78851:3
	output wire tx_valid_o;
	// Trace: design.sv:78852:3
	input [31:0] rx_data_i;
	// Trace: design.sv:78853:3
	output wire rx_ready_o;
	// Trace: design.sv:78856:3
	localparam signed [31:0] spi_host_reg_pkg_BlockAw = 6;
	localparam signed [31:0] AW = spi_host_reg_pkg_BlockAw;
	// Trace: design.sv:78858:3
	wire [5:0] tx_addr;
	// Trace: design.sv:78860:3
	wire tx_win_error;
	// Trace: design.sv:78861:3
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_TXDATA_OFFSET = 6'h2c;
	assign tx_win_error = (tx_win_i[68] == 1'b0) && (tx_addr != spi_host_reg_pkg_SPI_HOST_TXDATA_OFFSET);
	// Trace: design.sv:78864:3
	wire [5:0] rx_addr;
	// Trace: design.sv:78866:3
	wire rx_win_error;
	// Trace: design.sv:78867:3
	localparam [5:0] spi_host_reg_pkg_SPI_HOST_RXDATA_OFFSET = 6'h28;
	assign rx_win_error = (rx_win_i[68] == 1'b1) && (rx_addr != spi_host_reg_pkg_SPI_HOST_RXDATA_OFFSET);
	// Trace: design.sv:78877:5
	assign rx_ready_o = rx_win_i[69] & ~rx_win_i[68];
	// Trace: design.sv:78878:5
	assign rx_win_o[31-:32] = rx_data_i;
	// Trace: design.sv:78880:5
	assign rx_win_o[33] = rx_win_error;
	// Trace: design.sv:78881:5
	assign rx_win_o[32] = 1'b1;
	// Trace: design.sv:78882:5
	assign rx_addr = rx_win_i[63-:32];
	// Trace: design.sv:78884:5
	assign tx_valid_o = tx_win_i[69] & tx_win_i[68];
	// Trace: design.sv:78885:5
	assign tx_data_o = tx_win_i[31-:32];
	// Trace: design.sv:78886:5
	assign tx_be_o = tx_win_i[67-:4];
	// Trace: design.sv:78888:5
	assign tx_win_o[33] = tx_win_error;
	// Trace: design.sv:78889:5
	assign tx_win_o[31-:32] = 32'h00000000;
	// Trace: design.sv:78890:5
	assign tx_win_o[32] = 1'b1;
	// Trace: design.sv:78891:5
	assign tx_addr = tx_win_i[63-:32];
endmodule
module spi_host_CA356 (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	alert_rx_i,
	alert_tx_o,
	cio_sck_o,
	cio_sck_en_o,
	cio_csb_o,
	cio_csb_en_o,
	cio_sd_o,
	cio_sd_en_o,
	cio_sd_i,
	passthrough_i,
	passthrough_o,
	rx_valid_o,
	tx_ready_o,
	intr_error_o,
	intr_spi_event_o
);
	reg _sv2v_0;
	// removed import spi_host_reg_pkg::*;
	// Trace: design.sv:78907:13
	localparam signed [31:0] spi_host_reg_pkg_NumAlerts = 1;
	parameter [0:0] AlertAsyncOn = {spi_host_reg_pkg_NumAlerts {1'b1}};
	// Trace: design.sv:78908:18
	// removed localparam type reg_req_t
	// Trace: design.sv:78909:18
	// removed localparam type reg_rsp_t
	// Trace: design.sv:78911:3
	input clk_i;
	// Trace: design.sv:78912:3
	input rst_ni;
	// Trace: design.sv:78915:3
	input wire [69:0] reg_req_i;
	// Trace: design.sv:78916:3
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:78919:3
	// removed localparam type prim_alert_pkg_alert_rx_t
	input wire [3:0] alert_rx_i;
	// Trace: design.sv:78920:3
	// removed localparam type prim_alert_pkg_alert_tx_t
	output wire [1:0] alert_tx_o;
	// Trace: design.sv:78923:3
	output wire cio_sck_o;
	// Trace: design.sv:78924:3
	output wire cio_sck_en_o;
	// Trace: design.sv:78925:3
	localparam signed [31:0] spi_host_reg_pkg_NumCS = 2;
	output wire [1:0] cio_csb_o;
	// Trace: design.sv:78926:3
	output wire [1:0] cio_csb_en_o;
	// Trace: design.sv:78927:3
	output wire [3:0] cio_sd_o;
	// Trace: design.sv:78928:3
	output wire [3:0] cio_sd_en_o;
	// Trace: design.sv:78929:3
	input [3:0] cio_sd_i;
	// Trace: design.sv:78932:3
	// removed localparam type spi_device_pkg_passthrough_req_t
	input wire [13:0] passthrough_i;
	// Trace: design.sv:78933:3
	// removed localparam type spi_device_pkg_passthrough_rsp_t
	output wire [3:0] passthrough_o;
	// Trace: design.sv:78936:3
	output wire rx_valid_o;
	// Trace: design.sv:78937:3
	output wire tx_ready_o;
	// Trace: design.sv:78939:3
	output wire intr_error_o;
	// Trace: design.sv:78940:3
	output wire intr_spi_event_o;
	// Trace: design.sv:78943:3
	// removed import spi_host_cmd_pkg::*;
	// Trace: design.sv:78945:3
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_alert_test_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_command_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_configopts_mreg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_control_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_csid_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_error_enable_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_error_status_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_event_enable_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_intr_enable_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_intr_state_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_intr_test_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_reg2hw_t
	wire [172:0] reg2hw;
	// Trace: design.sv:78946:3
	// removed localparam type spi_host_reg_pkg_spi_host_hw2reg_error_status_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_hw2reg_intr_state_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_hw2reg_status_reg_t
	// removed localparam type spi_host_reg_pkg_spi_host_hw2reg_t
	wire [60:0] hw2reg;
	// Trace: design.sv:78948:3
	wire [139:0] fifo_win_h2d;
	// Trace: design.sv:78949:3
	wire [67:0] fifo_win_d2h;
	// Trace: design.sv:78952:3
	wire [0:0] alert_test;
	wire [0:0] alerts;
	// Trace: design.sv:78953:3
	spi_host_reg_top_3E795 u_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(reg_req_i),
		.reg_rsp_o(reg_rsp_o),
		.reg_req_win_o(fifo_win_h2d),
		.reg_rsp_win_i(fifo_win_d2h),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:78970:3
	assign alerts[0] = 1'b0;
	// Trace: design.sv:78971:3
	assign alert_test = {reg2hw[164] & reg2hw[163]};
	// Trace: design.sv:78976:3
	genvar _gv_i_87;
	generate
		for (_gv_i_87 = 0; _gv_i_87 < spi_host_reg_pkg_NumAlerts; _gv_i_87 = _gv_i_87 + 1) begin : gen_alert_tx
			localparam i = _gv_i_87;
			// Trace: design.sv:78977:5
			prim_alert_sender #(
				.AsyncOn(AlertAsyncOn[i]),
				.IsFatal(1'b1)
			) u_prim_alert_sender(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.alert_test_i(alert_test[i]),
				.alert_req_i(alerts[0]),
				.alert_ack_o(),
				.alert_state_o(),
				.alert_rx_i(alert_rx_i[i * 4+:4]),
				.alert_tx_o(alert_tx_o[i * 2+:2])
			);
		end
	endgenerate
	// Trace: design.sv:78992:3
	wire sck;
	// Trace: design.sv:78993:3
	wire [1:0] csb;
	// Trace: design.sv:78994:3
	wire [3:0] sd_out;
	// Trace: design.sv:78995:3
	wire [3:0] sd_en;
	wire [3:0] sd_en_core;
	// Trace: design.sv:78996:3
	wire [3:0] sd_i;
	// Trace: design.sv:78997:3
	wire output_en;
	// Trace: design.sv:78999:3
	assign output_en = reg2hw[146];
	// Trace: design.sv:79001:3
	assign sd_en = (output_en ? sd_en_core : 4'h0);
	// Trace: design.sv:79003:3
	generate
		if (1) begin : gen_passthrough_ignore
			// Trace: design.sv:79033:5
			assign cio_sck_o = sck;
			// Trace: design.sv:79034:5
			assign cio_sck_en_o = output_en;
			// Trace: design.sv:79035:5
			assign cio_csb_o = csb;
			// Trace: design.sv:79036:5
			assign cio_csb_en_o = {spi_host_reg_pkg_NumCS {output_en}};
			// Trace: design.sv:79037:5
			assign cio_sd_o = sd_out;
			// Trace: design.sv:79038:5
			assign cio_sd_en_o = sd_en;
			// Trace: design.sv:79040:5
			wire unused_pt_en;
			// Trace: design.sv:79041:5
			wire unused_pt_sck;
			// Trace: design.sv:79042:5
			wire unused_pt_sck_en;
			// Trace: design.sv:79043:5
			wire unused_pt_csb;
			// Trace: design.sv:79044:5
			wire unused_pt_csb_en;
			// Trace: design.sv:79045:5
			wire [3:0] unused_pt_sd_out;
			// Trace: design.sv:79046:5
			wire [3:0] unused_pt_sd_en;
			// Trace: design.sv:79048:5
			assign unused_pt_en = passthrough_i[13];
			// Trace: design.sv:79049:5
			assign unused_pt_sck = passthrough_i[12];
			// Trace: design.sv:79050:5
			assign unused_pt_sck_en = passthrough_i[10];
			// Trace: design.sv:79051:5
			assign unused_pt_csb = passthrough_i[9];
			// Trace: design.sv:79052:5
			assign unused_pt_csb_en = passthrough_i[8];
			// Trace: design.sv:79053:5
			assign unused_pt_sd_out = passthrough_i[7-:4];
			// Trace: design.sv:79054:5
			assign unused_pt_sd_en = passthrough_i[3-:4];
		end
	endgenerate
	// Trace: design.sv:79058:3
	assign passthrough_o[3-:4] = cio_sd_i;
	// Trace: design.sv:79059:3
	assign sd_i = cio_sd_i;
	// Trace: design.sv:79061:3
	localparam [0:0] spi_host_reg_pkg_ByteOrder = 1;
	assign hw2reg[31] = spi_host_reg_pkg_ByteOrder;
	// Trace: design.sv:79062:3
	assign hw2reg[30] = 1'b1;
	// Trace: design.sv:79064:3
	wire command_valid;
	// Trace: design.sv:79065:3
	wire core_command_valid;
	// Trace: design.sv:79066:3
	wire command_busy;
	// Trace: design.sv:79067:3
	wire core_command_ready;
	// Trace: design.sv:79069:3
	function automatic integer prim_util_pkg_vbits;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:74:36
		input integer value;
		// Trace: ../src/lowrisc_prim_util_0.1/rtl/prim_util_pkg.sv:85:5
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] spi_host_cmd_pkg_CSW = prim_util_pkg_vbits(spi_host_reg_pkg_NumCS);
	// removed localparam type spi_host_cmd_pkg_configopts_t
	// removed localparam type spi_host_cmd_pkg_segment_t
	// removed localparam type spi_host_cmd_pkg_command_t
	wire [spi_host_cmd_pkg_CSW + 59:0] core_command;
	reg [spi_host_cmd_pkg_CSW + 59:0] command;
	// Trace: design.sv:79070:3
	wire error_csid_inval;
	// Trace: design.sv:79071:3
	wire error_cmd_inval;
	// Trace: design.sv:79072:3
	wire error_busy;
	// Trace: design.sv:79073:3
	wire test_csid_inval;
	// Trace: design.sv:79074:3
	reg test_dir_inval;
	// Trace: design.sv:79075:3
	reg test_speed_inval;
	// Trace: design.sv:79077:3
	assign test_csid_inval = reg2hw[81-:32] >= spi_host_reg_pkg_NumCS;
	// Trace: design.sv:79079:3
	// removed localparam type spi_host_cmd_pkg_reg_direction_t
	// removed localparam type spi_host_cmd_pkg_speed_t
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:79080:5
		test_speed_inval = 1'b1;
		// Trace: design.sv:79081:5
		test_dir_inval = 1'b1;
		// Trace: design.sv:79082:5
		(* full_case, parallel_case *)
		case (reg2hw[22-:2])
			2'b00: begin
				// Trace: design.sv:79084:9
				test_dir_inval = 1'b0;
				// Trace: design.sv:79085:9
				test_speed_inval = 1'b0;
			end
			2'b01, 2'b10: begin
				// Trace: design.sv:79088:9
				test_dir_inval = reg2hw[19-:2] == 2'b11;
				// Trace: design.sv:79089:9
				test_speed_inval = 1'b0;
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:79096:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:79097:5
		command[56] = 1'b0;
		// Trace: design.sv:79098:5
		command[57] = 1'b0;
		// Trace: design.sv:79099:5
		(* full_case, parallel_case *)
		case (reg2hw[19-:2])
			2'b01:
				// Trace: design.sv:79101:9
				command[56] = 1'b1;
			2'b10:
				// Trace: design.sv:79104:9
				command[57] = 1'b1;
			2'b11: begin
				// Trace: design.sv:79107:9
				command[56] = 1'b1;
				// Trace: design.sv:79108:9
				command[57] = 1'b1;
			end
			default:
				;
		endcase
	end
	// Trace: design.sv:79115:3
	assign error_csid_inval = (command_valid & ~command_busy) & test_csid_inval;
	// Trace: design.sv:79117:3
	assign error_cmd_inval = (command_valid & ~command_busy) & (test_speed_inval | test_dir_inval);
	// Trace: design.sv:79120:3
	wire [30:0] configopts;
	// Trace: design.sv:79122:3
	generate
		if (1) begin : gen_multiple_devices
			// Trace: design.sv:79126:5
			wire [spi_host_cmd_pkg_CSW - 1:0] csid;
			// Trace: design.sv:79127:5
			assign csid = (test_csid_inval ? {spi_host_cmd_pkg_CSW {1'sb0}} : reg2hw[spi_host_cmd_pkg_CSW + 49:50]);
			// Trace: design.sv:79128:5
			assign configopts = reg2hw[82 + (csid * 31)+:31];
			// Trace: design.sv:79129:5
			wire [((spi_host_cmd_pkg_CSW + 59) >= 60 ? spi_host_cmd_pkg_CSW + 0 : 61 - (spi_host_cmd_pkg_CSW + 59)) * 1:1] sv2v_tmp_D6B78;
			assign sv2v_tmp_D6B78 = csid;
			always @(*) command[spi_host_cmd_pkg_CSW + 59-:((spi_host_cmd_pkg_CSW + 59) >= 60 ? spi_host_cmd_pkg_CSW + 0 : 61 - (spi_host_cmd_pkg_CSW + 59))] = sv2v_tmp_D6B78;
		end
	endgenerate
	// Trace: design.sv:79132:3
	wire [16:1] sv2v_tmp_8C1C9;
	assign sv2v_tmp_8C1C9 = configopts[30-:16];
	always @(*) command[30-:16] = sv2v_tmp_8C1C9;
	// Trace: design.sv:79133:3
	wire [4:1] sv2v_tmp_3279F;
	assign sv2v_tmp_3279F = configopts[14-:4];
	always @(*) command[14-:4] = sv2v_tmp_3279F;
	// Trace: design.sv:79134:3
	wire [4:1] sv2v_tmp_4844B;
	assign sv2v_tmp_4844B = configopts[6-:4];
	always @(*) command[10-:4] = sv2v_tmp_4844B;
	// Trace: design.sv:79135:3
	wire [4:1] sv2v_tmp_BC40B;
	assign sv2v_tmp_BC40B = configopts[10-:4];
	always @(*) command[6-:4] = sv2v_tmp_BC40B;
	// Trace: design.sv:79136:3
	wire [1:1] sv2v_tmp_4FA47;
	assign sv2v_tmp_4FA47 = configopts[2];
	always @(*) command[2] = sv2v_tmp_4FA47;
	// Trace: design.sv:79137:3
	wire [1:1] sv2v_tmp_1B667;
	assign sv2v_tmp_1B667 = configopts[1];
	always @(*) command[1] = sv2v_tmp_1B667;
	// Trace: design.sv:79138:3
	wire [1:1] sv2v_tmp_45EDB;
	assign sv2v_tmp_45EDB = configopts[-0];
	always @(*) command[0] = sv2v_tmp_45EDB;
	// Trace: design.sv:79140:3
	wire [24:1] sv2v_tmp_49692;
	assign sv2v_tmp_49692 = reg2hw[49-:24];
	always @(*) command[55-:24] = sv2v_tmp_49692;
	// Trace: design.sv:79141:3
	wire [1:1] sv2v_tmp_55901;
	assign sv2v_tmp_55901 = reg2hw[24];
	always @(*) command[31] = sv2v_tmp_55901;
	// Trace: design.sv:79142:3
	wire [2:1] sv2v_tmp_C9B77;
	assign sv2v_tmp_C9B77 = reg2hw[22-:2];
	always @(*) command[59-:2] = sv2v_tmp_C9B77;
	// Trace: design.sv:79145:3
	wire [3:0] cmd_qes;
	// Trace: design.sv:79147:3
	assign cmd_qes = {reg2hw[25], reg2hw[20], reg2hw[17], reg2hw[23]};
	// Trace: design.sv:79155:3
	assign command_valid = |cmd_qes;
	// Trace: design.sv:79157:3
	wire active;
	// Trace: design.sv:79158:3
	wire rx_stall;
	// Trace: design.sv:79159:3
	wire tx_stall;
	// Trace: design.sv:79161:3
	assign hw2reg[13] = ~command_busy;
	// Trace: design.sv:79162:3
	assign hw2reg[15] = active;
	// Trace: design.sv:79163:3
	assign hw2reg[29] = rx_stall;
	// Trace: design.sv:79164:3
	assign hw2reg[21] = tx_stall;
	// Trace: design.sv:79166:3
	assign hw2reg[12] = 1'b1;
	// Trace: design.sv:79167:3
	assign hw2reg[14] = 1'b1;
	// Trace: design.sv:79168:3
	assign hw2reg[28] = 1'b1;
	// Trace: design.sv:79169:3
	assign hw2reg[20] = 1'b1;
	// Trace: design.sv:79171:3
	wire sw_rst;
	// Trace: design.sv:79173:3
	wire [3:0] cmd_qd;
	// Trace: design.sv:79175:3
	localparam signed [31:0] spi_host_reg_pkg_CmdDepth = 4;
	spi_host_command_queue #(.CmdDepth(spi_host_reg_pkg_CmdDepth)) u_cmd_queue(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.command_i(command),
		.command_valid_i(command_valid),
		.command_busy_o(command_busy),
		.core_command_o(core_command),
		.core_command_valid_o(core_command_valid),
		.core_command_ready_i(core_command_ready),
		.error_busy_o(error_busy),
		.qd_o(cmd_qd),
		.sw_rst_i(sw_rst)
	);
	// Trace: design.sv:79191:3
	wire [31:0] tx_data;
	// Trace: design.sv:79192:3
	wire [3:0] tx_be;
	// Trace: design.sv:79193:3
	wire tx_valid;
	// Trace: design.sv:79194:3
	wire tx_ready;
	// Trace: design.sv:79196:3
	wire [31:0] rx_data;
	// Trace: design.sv:79197:3
	wire rx_valid;
	// Trace: design.sv:79198:3
	wire rx_ready;
	// Trace: design.sv:79200:3
	spi_host_window_9C1FC u_window(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rx_win_i(fifo_win_h2d[0+:70]),
		.rx_win_o(fifo_win_d2h[0+:34]),
		.tx_win_i(fifo_win_h2d[70+:70]),
		.tx_win_o(fifo_win_d2h[34+:34]),
		.tx_data_o(tx_data),
		.tx_be_o(tx_be),
		.tx_valid_o(tx_valid),
		.rx_data_i(rx_data),
		.rx_ready_o(rx_ready)
	);
	// Trace: design.sv:79217:3
	wire [31:0] core_tx_data;
	// Trace: design.sv:79218:3
	wire [3:0] core_tx_be;
	// Trace: design.sv:79219:3
	wire core_tx_valid;
	// Trace: design.sv:79220:3
	wire core_tx_ready;
	// Trace: design.sv:79222:3
	wire [31:0] core_rx_data;
	// Trace: design.sv:79223:3
	wire core_rx_valid;
	// Trace: design.sv:79224:3
	wire core_rx_ready;
	// Trace: design.sv:79226:3
	wire [7:0] rx_watermark;
	// Trace: design.sv:79227:3
	wire [7:0] tx_watermark;
	// Trace: design.sv:79228:3
	wire [7:0] rx_qd;
	// Trace: design.sv:79229:3
	wire [7:0] tx_qd;
	// Trace: design.sv:79231:3
	wire tx_empty;
	wire tx_full;
	wire tx_wm;
	// Trace: design.sv:79232:3
	wire rx_empty;
	wire rx_full;
	wire rx_wm;
	// Trace: design.sv:79234:3
	assign rx_valid_o = rx_valid;
	// Trace: design.sv:79235:3
	assign tx_ready_o = tx_ready;
	// Trace: design.sv:79237:3
	assign rx_watermark = reg2hw[162-:8];
	// Trace: design.sv:79238:3
	assign tx_watermark = reg2hw[154-:8];
	// Trace: design.sv:79240:3
	assign hw2reg[56-:8] = tx_qd;
	// Trace: design.sv:79241:3
	assign hw2reg[47-:8] = rx_qd;
	// Trace: design.sv:79242:3
	assign hw2reg[38-:4] = cmd_qd;
	// Trace: design.sv:79243:3
	assign hw2reg[23] = tx_wm;
	// Trace: design.sv:79244:3
	assign hw2reg[33] = rx_wm;
	// Trace: design.sv:79245:3
	assign hw2reg[27] = rx_empty;
	// Trace: design.sv:79246:3
	assign hw2reg[19] = tx_empty;
	// Trace: design.sv:79247:3
	assign hw2reg[25] = rx_full;
	// Trace: design.sv:79248:3
	assign hw2reg[17] = tx_full;
	// Trace: design.sv:79250:3
	assign hw2reg[48] = 1'b1;
	// Trace: design.sv:79251:3
	assign hw2reg[39] = 1'b1;
	// Trace: design.sv:79252:3
	assign hw2reg[34] = 1'b1;
	// Trace: design.sv:79253:3
	assign hw2reg[22] = 1'b1;
	// Trace: design.sv:79254:3
	assign hw2reg[32] = 1'b1;
	// Trace: design.sv:79255:3
	assign hw2reg[26] = 1'b1;
	// Trace: design.sv:79256:3
	assign hw2reg[18] = 1'b1;
	// Trace: design.sv:79257:3
	assign hw2reg[24] = 1'b1;
	// Trace: design.sv:79258:3
	assign hw2reg[16] = 1'b1;
	// Trace: design.sv:79260:3
	wire error_overflow;
	wire error_underflow;
	// Trace: design.sv:79261:3
	wire error_access_inval;
	// Trace: design.sv:79265:3
	assign error_overflow = tx_valid & ~tx_ready;
	// Trace: design.sv:79266:3
	assign error_underflow = rx_ready & ~rx_valid;
	// Trace: design.sv:79267:3
	reg access_valid;
	// Trace: design.sv:79268:3
	assign error_access_inval = tx_valid & ~access_valid;
	// Trace: design.sv:79270:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:79271:5
		(* full_case, parallel_case *)
		case (tx_be)
			4'b1000, 4'b0100, 4'b0010, 4'b0001, 4'b1100, 4'b0110, 4'b0011, 4'b1111:
				// Trace: design.sv:79280:9
				access_valid = 1'b1;
			default:
				// Trace: design.sv:79283:9
				access_valid = 1'b0;
		endcase
	end
	// Trace: design.sv:79288:3
	wire tx_valid_checked;
	// Trace: design.sv:79289:3
	assign tx_valid_checked = (tx_valid & ~error_overflow) & ~error_access_inval;
	// Trace: design.sv:79295:3
	localparam signed [31:0] spi_host_reg_pkg_RxDepth = 64;
	localparam signed [31:0] spi_host_reg_pkg_TxDepth = 72;
	spi_host_data_fifos #(
		.TxDepth(spi_host_reg_pkg_TxDepth),
		.RxDepth(spi_host_reg_pkg_RxDepth),
		.SwapBytes(~spi_host_reg_pkg_ByteOrder)
	) u_data_fifos(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tx_data_i(tx_data),
		.tx_be_i(tx_be),
		.tx_valid_i(tx_valid_checked),
		.tx_ready_o(tx_ready),
		.tx_watermark_i(tx_watermark),
		.core_tx_data_o(core_tx_data),
		.core_tx_be_o(core_tx_be),
		.core_tx_valid_o(core_tx_valid),
		.core_tx_ready_i(core_tx_ready),
		.core_rx_data_i(core_rx_data),
		.core_rx_valid_i(core_rx_valid),
		.core_rx_ready_o(core_rx_ready),
		.rx_data_o(rx_data),
		.rx_valid_o(rx_valid),
		.rx_ready_i(rx_ready),
		.rx_watermark_i(rx_watermark),
		.tx_empty_o(tx_empty),
		.tx_full_o(tx_full),
		.tx_qd_o(tx_qd),
		.tx_wm_o(tx_wm),
		.rx_empty_o(rx_empty),
		.rx_full_o(rx_full),
		.rx_qd_o(rx_qd),
		.rx_wm_o(rx_wm),
		.sw_rst_i(sw_rst)
	);
	// Trace: design.sv:79335:3
	wire en_sw;
	// Trace: design.sv:79336:3
	wire enb_error;
	// Trace: design.sv:79337:3
	wire en;
	// Trace: design.sv:79339:3
	assign en = en_sw & ~enb_error;
	// Trace: design.sv:79340:3
	assign sw_rst = reg2hw[145];
	// Trace: design.sv:79341:3
	assign en_sw = reg2hw[144];
	// Trace: design.sv:79343:3
	spi_host_core #(.NumCS(spi_host_reg_pkg_NumCS)) u_spi_core(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.command_i(core_command),
		.command_valid_i(core_command_valid),
		.command_ready_o(core_command_ready),
		.en_i(en),
		.tx_data_i(core_tx_data),
		.tx_be_i(core_tx_be),
		.tx_valid_i(core_tx_valid),
		.tx_ready_o(core_tx_ready),
		.rx_data_o(core_rx_data),
		.rx_valid_o(core_rx_valid),
		.rx_ready_i(core_rx_ready),
		.sck_o(sck),
		.csb_o(csb),
		.sd_o(sd_out),
		.sd_en_o(sd_en_core),
		.sd_i(sd_i),
		.rx_stall_o(rx_stall),
		.tx_stall_o(tx_stall),
		.sw_rst_i(sw_rst),
		.active_o(active)
	);
	// Trace: design.sv:79371:3
	wire event_error;
	// Trace: design.sv:79373:3
	wire [5:0] error_vec;
	// Trace: design.sv:79374:3
	wire [5:0] error_mask;
	// Trace: design.sv:79375:3
	wire [5:0] sw_error_status;
	// Trace: design.sv:79377:3
	assign error_vec = {error_access_inval, error_csid_inval, error_cmd_inval, error_underflow, error_overflow, error_busy};
	// Trace: design.sv:79391:3
	assign error_mask = {1'b1, reg2hw[12], reg2hw[13], reg2hw[14], reg2hw[15], reg2hw[16]};
	// Trace: design.sv:79400:3
	assign hw2reg[1] = error_access_inval;
	// Trace: design.sv:79401:3
	assign hw2reg[3] = error_csid_inval;
	// Trace: design.sv:79402:3
	assign hw2reg[5] = error_cmd_inval;
	// Trace: design.sv:79403:3
	assign hw2reg[7] = error_underflow;
	// Trace: design.sv:79404:3
	assign hw2reg[9] = error_overflow;
	// Trace: design.sv:79405:3
	assign hw2reg[11] = error_busy;
	// Trace: design.sv:79409:3
	assign hw2reg[0] = error_access_inval;
	// Trace: design.sv:79410:3
	assign hw2reg[2] = error_csid_inval;
	// Trace: design.sv:79411:3
	assign hw2reg[4] = error_cmd_inval;
	// Trace: design.sv:79412:3
	assign hw2reg[6] = error_underflow;
	// Trace: design.sv:79413:3
	assign hw2reg[8] = error_overflow;
	// Trace: design.sv:79414:3
	assign hw2reg[10] = error_busy;
	// Trace: design.sv:79416:3
	assign sw_error_status[5] = reg2hw[6];
	// Trace: design.sv:79417:3
	assign sw_error_status[4] = reg2hw[7];
	// Trace: design.sv:79418:3
	assign sw_error_status[3] = reg2hw[8];
	// Trace: design.sv:79419:3
	assign sw_error_status[2] = reg2hw[9];
	// Trace: design.sv:79420:3
	assign sw_error_status[1] = reg2hw[10];
	// Trace: design.sv:79421:3
	assign sw_error_status[0] = reg2hw[11];
	// Trace: design.sv:79423:3
	assign event_error = |(error_vec & error_mask);
	// Trace: design.sv:79424:3
	assign enb_error = |sw_error_status;
	// Trace: design.sv:79426:3
	prim_intr_hw #(.Width(1)) intr_hw_error(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_error),
		.reg2hw_intr_enable_q_i(reg2hw[170]),
		.reg2hw_intr_test_q_i(reg2hw[168]),
		.reg2hw_intr_test_qe_i(reg2hw[167]),
		.reg2hw_intr_state_q_i(reg2hw[172]),
		.hw2reg_intr_state_de_o(hw2reg[59]),
		.hw2reg_intr_state_d_o(hw2reg[60]),
		.intr_o(intr_error_o)
	);
	// Trace: design.sv:79439:3
	wire event_spi_event;
	// Trace: design.sv:79440:3
	wire event_idle;
	wire event_ready;
	wire event_tx_wm;
	wire event_rx_wm;
	wire event_tx_empty;
	wire event_rx_full;
	// Trace: design.sv:79441:3
	wire [5:0] event_vector;
	// Trace: design.sv:79442:3
	wire [5:0] event_mask;
	// Trace: design.sv:79444:3
	assign event_vector = {event_idle, event_ready, event_tx_wm, event_rx_wm, event_tx_empty, event_rx_full};
	// Trace: design.sv:79449:3
	assign event_mask = {reg2hw[0], reg2hw[1], reg2hw[2], reg2hw[3], reg2hw[4], reg2hw[5]};
	// Trace: design.sv:79458:3
	assign event_spi_event = |(event_vector & event_mask);
	// Trace: design.sv:79460:3
	wire idle_d;
	reg idle_q;
	// Trace: design.sv:79461:3
	wire ready_d;
	reg ready_q;
	// Trace: design.sv:79462:3
	wire tx_wm_d;
	reg tx_wm_q;
	// Trace: design.sv:79463:3
	wire rx_wm_d;
	reg rx_wm_q;
	// Trace: design.sv:79464:3
	wire tx_empty_d;
	reg tx_empty_q;
	// Trace: design.sv:79465:3
	wire rx_full_d;
	reg rx_full_q;
	// Trace: design.sv:79467:3
	assign event_idle = idle_d & ~idle_q;
	// Trace: design.sv:79468:3
	assign idle_d = ~active;
	// Trace: design.sv:79469:3
	assign event_ready = ready_d & ~ready_q;
	// Trace: design.sv:79470:3
	assign ready_d = ~command_busy;
	// Trace: design.sv:79471:3
	assign event_tx_wm = tx_wm_d & ~tx_wm_q;
	// Trace: design.sv:79472:3
	assign tx_wm_d = tx_wm;
	// Trace: design.sv:79473:3
	assign event_rx_wm = rx_wm_d & ~rx_wm_q;
	// Trace: design.sv:79474:3
	assign rx_wm_d = rx_wm;
	// Trace: design.sv:79475:3
	assign event_tx_empty = tx_empty_d & ~tx_empty_q;
	// Trace: design.sv:79476:3
	assign tx_empty_d = tx_empty;
	// Trace: design.sv:79477:3
	assign event_rx_full = rx_full_d & ~rx_full_q;
	// Trace: design.sv:79478:3
	assign rx_full_d = rx_full;
	// Trace: design.sv:79480:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:79481:5
		if (!rst_ni) begin
			// Trace: design.sv:79482:7
			idle_q <= 1'b0;
			// Trace: design.sv:79483:7
			ready_q <= 1'b0;
			// Trace: design.sv:79484:7
			tx_wm_q <= 1'b0;
			// Trace: design.sv:79485:7
			rx_wm_q <= 1'b0;
			// Trace: design.sv:79486:7
			tx_empty_q <= 1'b0;
			// Trace: design.sv:79487:7
			rx_full_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:79489:7
			idle_q <= idle_d;
			// Trace: design.sv:79490:7
			ready_q <= ready_d;
			// Trace: design.sv:79491:7
			tx_wm_q <= tx_wm_d;
			// Trace: design.sv:79492:7
			rx_wm_q <= rx_wm_d;
			// Trace: design.sv:79493:7
			tx_empty_q <= tx_empty_d;
			// Trace: design.sv:79494:7
			rx_full_q <= rx_full_d;
		end
	// Trace: design.sv:79498:3
	prim_intr_hw #(.Width(1)) intr_hw_spi_event(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_spi_event),
		.reg2hw_intr_enable_q_i(reg2hw[169]),
		.reg2hw_intr_test_q_i(reg2hw[166]),
		.reg2hw_intr_test_qe_i(reg2hw[165]),
		.reg2hw_intr_state_q_i(reg2hw[171]),
		.hw2reg_intr_state_de_o(hw2reg[57]),
		.hw2reg_intr_state_d_o(hw2reg[58]),
		.intr_o(intr_spi_event_o)
	);
	initial _sv2v_0 = 0;
endmodule
module tlul_err_resp (
	clk_i,
	rst_ni,
	tl_h_i,
	tl_h_o
);
	// Trace: design.sv:79536:3
	input clk_i;
	// Trace: design.sv:79537:3
	input rst_ni;
	// Trace: design.sv:79538:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_h_i;
	// Trace: design.sv:79539:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o;
	// Trace: design.sv:79541:3
	// removed import tlul_pkg::*;
	// Trace: design.sv:79543:3
	reg [2:0] err_opcode;
	// Trace: design.sv:79544:3
	reg [7:0] err_source;
	// Trace: design.sv:79545:3
	reg [top_pkg_TL_SZW - 1:0] err_size;
	// Trace: design.sv:79546:3
	reg err_req_pending;
	reg err_rsp_pending;
	// Trace: design.sv:79548:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:79549:5
		if (!rst_ni) begin
			// Trace: design.sv:79550:7
			err_req_pending <= 1'b0;
			// Trace: design.sv:79551:7
			err_source <= {top_pkg_TL_AIW {1'b0}};
			// Trace: design.sv:79552:7
			err_opcode <= 3'h4;
			// Trace: design.sv:79553:7
			err_size <= 1'sb0;
		end
		else if (tl_h_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] && tl_h_o[0]) begin
			// Trace: design.sv:79555:7
			err_req_pending <= 1'b1;
			// Trace: design.sv:79556:7
			err_source <= tl_h_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)];
			// Trace: design.sv:79557:7
			err_opcode <= tl_h_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)];
			// Trace: design.sv:79558:7
			err_size <= tl_h_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)];
		end
		else if (!err_rsp_pending)
			// Trace: design.sv:79560:7
			err_req_pending <= 1'b0;
	// Trace: design.sv:79564:3
	assign tl_h_o[0] = ~err_rsp_pending & ~(err_req_pending & ~tl_h_i[0]);
	// Trace: design.sv:79565:3
	assign tl_h_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] = err_req_pending | err_rsp_pending;
	// Trace: design.sv:79566:3
	assign tl_h_o[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)] = 1'sb1;
	// Trace: design.sv:79567:3
	assign tl_h_o[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)] = err_source;
	// Trace: design.sv:79568:3
	assign tl_h_o[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)] = 1'sb0;
	// Trace: design.sv:79569:3
	assign tl_h_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = 1'sb0;
	// Trace: design.sv:79570:3
	assign tl_h_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)] = err_size;
	// Trace: design.sv:79571:3
	assign tl_h_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = (err_opcode == 3'h4 ? 3'h1 : 3'h0);
	// Trace: design.sv:79572:3
	assign tl_h_o[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))] = 1'sb0;
	// Trace: design.sv:79573:3
	assign tl_h_o[1] = 1'b1;
	// Trace: design.sv:79575:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:79576:5
		if (!rst_ni)
			// Trace: design.sv:79577:7
			err_rsp_pending <= 1'b0;
		else if ((err_req_pending || err_rsp_pending) && !tl_h_i[0])
			// Trace: design.sv:79579:7
			err_rsp_pending <= 1'b1;
		else
			// Trace: design.sv:79581:7
			err_rsp_pending <= 1'b0;
	// Trace: design.sv:79586:3
	wire unused_tl_h;
	// Trace: design.sv:79587:3
	assign unused_tl_h = &{1'b0, tl_h_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)], tl_h_i[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)], tl_h_i[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))], tl_h_i[53-:32], tl_h_i[21-:21], tl_h_i[0]};
endmodule
module tlul_socket_1n (
	clk_i,
	rst_ni,
	tl_h_i,
	tl_h_o,
	tl_d_o,
	tl_d_i,
	dev_select_i
);
	reg _sv2v_0;
	// Trace: design.sv:79631:13
	parameter [31:0] N = 4;
	// Trace: design.sv:79632:13
	parameter [0:0] HReqPass = 1'b1;
	// Trace: design.sv:79633:13
	parameter [0:0] HRspPass = 1'b1;
	// Trace: design.sv:79634:13
	parameter [N - 1:0] DReqPass = {N {1'b1}};
	// Trace: design.sv:79635:13
	parameter [N - 1:0] DRspPass = {N {1'b1}};
	// Trace: design.sv:79636:13
	parameter [3:0] HReqDepth = 4'h2;
	// Trace: design.sv:79637:13
	parameter [3:0] HRspDepth = 4'h2;
	// Trace: design.sv:79638:13
	parameter [(N * 4) - 1:0] DReqDepth = {N {4'h2}};
	// Trace: design.sv:79639:13
	parameter [(N * 4) - 1:0] DRspDepth = {N {4'h2}};
	// Trace: design.sv:79640:14
	localparam [31:0] NWD = $clog2(N + 1);
	// Trace: design.sv:79642:3
	input clk_i;
	// Trace: design.sv:79643:3
	input rst_ni;
	// Trace: design.sv:79644:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_h_i;
	// Trace: design.sv:79645:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o;
	// Trace: design.sv:79646:3
	output wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? (N * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)) - 1 : (N * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 20)):(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21)] tl_d_o;
	// Trace: design.sv:79647:3
	input wire [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (N * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 1 : (N * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 0)):((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)] tl_d_i;
	// Trace: design.sv:79648:3
	input [NWD - 1:0] dev_select_i;
	// Trace: design.sv:79659:3
	wire [NWD - 1:0] dev_select_t;
	// Trace: design.sv:79661:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_t_o;
	// Trace: design.sv:79662:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_t_i;
	// Trace: design.sv:79664:3
	tlul_fifo_sync #(
		.ReqPass(HReqPass),
		.RspPass(HRspPass),
		.ReqDepth(HReqDepth),
		.RspDepth(HRspDepth),
		.SpareReqW(NWD)
	) fifo_h(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(tl_h_i),
		.tl_h_o(tl_h_o),
		.tl_d_o(tl_t_o),
		.tl_d_i(tl_t_i),
		.spare_req_i(dev_select_i),
		.spare_req_o(dev_select_t),
		.spare_rsp_i(1'b0),
		.spare_rsp_o()
	);
	// Trace: design.sv:79686:3
	localparam signed [31:0] MaxOutstanding = 256;
	// Trace: design.sv:79687:3
	localparam signed [31:0] OutstandingW = 9;
	// Trace: design.sv:79688:3
	reg [8:0] num_req_outstanding;
	// Trace: design.sv:79689:3
	reg [NWD - 1:0] dev_select_outstanding;
	// Trace: design.sv:79690:3
	wire hold_all_requests;
	// Trace: design.sv:79691:3
	wire accept_t_req;
	wire accept_t_rsp;
	// Trace: design.sv:79693:3
	assign accept_t_req = tl_t_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] & tl_t_i[0];
	// Trace: design.sv:79694:3
	assign accept_t_rsp = tl_t_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & tl_t_o[0];
	// Trace: design.sv:79696:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:79697:5
		if (!rst_ni) begin
			// Trace: design.sv:79698:7
			num_req_outstanding <= 1'sb0;
			// Trace: design.sv:79699:7
			dev_select_outstanding <= 1'sb0;
		end
		else if (accept_t_req) begin
			// Trace: design.sv:79701:7
			if (!accept_t_rsp)
				// Trace: design.sv:79703:9
				num_req_outstanding <= num_req_outstanding + 1'b1;
			// Trace: design.sv:79705:7
			dev_select_outstanding <= dev_select_t;
		end
		else if (accept_t_rsp)
			// Trace: design.sv:79707:7
			num_req_outstanding <= num_req_outstanding - 1'b1;
	// Trace: design.sv:79711:3
	assign hold_all_requests = (num_req_outstanding != {9 {1'sb0}}) & (dev_select_t != dev_select_outstanding);
	// Trace: design.sv:79718:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_u_o [0:N + 0];
	// Trace: design.sv:79719:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_u_i [0:N + 0];
	// Trace: design.sv:79721:3
	genvar _gv_i_88;
	function automatic signed [NWD - 1:0] sv2v_cast_1D9BB_signed;
		input reg signed [NWD - 1:0] inp;
		sv2v_cast_1D9BB_signed = inp;
	endfunction
	generate
		for (_gv_i_88 = 0; _gv_i_88 < N; _gv_i_88 = _gv_i_88 + 1) begin : gen_u_o
			localparam i = _gv_i_88;
			// Trace: design.sv:79722:5
			assign tl_u_o[i][7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] = (tl_t_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] & (dev_select_t == sv2v_cast_1D9BB_signed(i))) & ~hold_all_requests;
			// Trace: design.sv:79725:5
			assign tl_u_o[i][6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] = tl_t_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)];
			// Trace: design.sv:79726:5
			assign tl_u_o[i][3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] = tl_t_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)];
			// Trace: design.sv:79727:5
			assign tl_u_o[i][top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)] = tl_t_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)];
			// Trace: design.sv:79728:5
			assign tl_u_o[i][top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)] = tl_t_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)];
			// Trace: design.sv:79729:5
			assign tl_u_o[i][top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)] = tl_t_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)];
			// Trace: design.sv:79730:5
			assign tl_u_o[i][top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))] = tl_t_o[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))];
			// Trace: design.sv:79731:5
			assign tl_u_o[i][53-:32] = tl_t_o[53-:32];
			// Trace: design.sv:79732:5
			assign tl_u_o[i][21-:21] = tl_t_o[21-:21];
		end
	endgenerate
	// Trace: design.sv:79735:3
	reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_t_p;
	// Trace: design.sv:79738:3
	reg hfifo_reqready;
	// Trace: design.sv:79739:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:79740:5
		hfifo_reqready = tl_u_i[N][0];
		// Trace: design.sv:79741:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:79741:10
			reg signed [31:0] idx;
			// Trace: design.sv:79741:10
			for (idx = 0; idx < N; idx = idx + 1)
				begin
					// Trace: design.sv:79743:7
					if (dev_select_t == sv2v_cast_1D9BB_signed(idx))
						// Trace: design.sv:79743:38
						hfifo_reqready = tl_u_i[idx][0];
				end
		end
		if (hold_all_requests)
			// Trace: design.sv:79745:28
			hfifo_reqready = 1'b0;
	end
	// Trace: design.sv:79749:3
	assign tl_t_i[0] = tl_t_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] & hfifo_reqready;
	// Trace: design.sv:79751:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:79752:5
		tl_t_p = tl_u_i[N];
		// Trace: design.sv:79753:5
		begin : sv2v_autoblock_2
			// Trace: design.sv:79753:10
			reg signed [31:0] idx;
			// Trace: design.sv:79753:10
			for (idx = 0; idx < N; idx = idx + 1)
				begin
					// Trace: design.sv:79754:7
					if (dev_select_outstanding == sv2v_cast_1D9BB_signed(idx))
						// Trace: design.sv:79754:48
						tl_t_p = tl_u_i[idx];
				end
		end
	end
	// Trace: design.sv:79757:3
	assign tl_t_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] = tl_t_p[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))];
	// Trace: design.sv:79758:3
	assign tl_t_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = tl_t_p[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)];
	// Trace: design.sv:79759:3
	assign tl_t_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = tl_t_p[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)];
	// Trace: design.sv:79760:3
	assign tl_t_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)] = tl_t_p[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)];
	// Trace: design.sv:79761:3
	assign tl_t_i[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)] = tl_t_p[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)];
	// Trace: design.sv:79762:3
	assign tl_t_i[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)] = tl_t_p[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)];
	// Trace: design.sv:79763:3
	assign tl_t_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)] = tl_t_p[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)];
	// Trace: design.sv:79764:3
	assign tl_t_i[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))] = tl_t_p[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))];
	// Trace: design.sv:79765:3
	assign tl_t_i[1] = tl_t_p[1];
	// Trace: design.sv:79769:3
	genvar _gv_i_89;
	generate
		for (_gv_i_89 = 0; _gv_i_89 < (N + 1); _gv_i_89 = _gv_i_89 + 1) begin : gen_u_o_d_ready
			localparam i = _gv_i_89;
			// Trace: design.sv:79770:5
			assign tl_u_o[i][0] = tl_t_o[0];
		end
	endgenerate
	// Trace: design.sv:79774:3
	genvar _gv_i_90;
	generate
		for (_gv_i_90 = 0; _gv_i_90 < N; _gv_i_90 = _gv_i_90 + 1) begin : gen_dfifo
			localparam i = _gv_i_90;
			// Trace: design.sv:79775:5
			tlul_fifo_sync #(
				.ReqPass(DReqPass[i]),
				.RspPass(DRspPass[i]),
				.ReqDepth(DReqDepth[i * 4+:4]),
				.RspDepth(DRspDepth[i * 4+:4])
			) fifo_d(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.tl_h_i(tl_u_o[i]),
				.tl_h_o(tl_u_i[i]),
				.tl_d_o(tl_d_o[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21) + (((N - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21)))+:(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 53) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21))]),
				.tl_d_i(tl_d_i[((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1) + (((N - 1) - i) * ((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)))+:((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))]),
				.spare_req_i(1'b0),
				.spare_req_o(),
				.spare_rsp_i(1'b0),
				.spare_rsp_o()
			);
		end
	endgenerate
	// Trace: design.sv:79793:3
	function automatic [NWD - 1:0] sv2v_cast_1D9BB;
		input reg [NWD - 1:0] inp;
		sv2v_cast_1D9BB = inp;
	endfunction
	assign tl_u_o[N][7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] = (tl_t_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] & (dev_select_t == sv2v_cast_1D9BB(N))) & ~hold_all_requests;
	// Trace: design.sv:79796:3
	assign tl_u_o[N][6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] = tl_t_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)];
	// Trace: design.sv:79797:3
	assign tl_u_o[N][3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] = tl_t_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)];
	// Trace: design.sv:79798:3
	assign tl_u_o[N][top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)] = tl_t_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)];
	// Trace: design.sv:79799:3
	assign tl_u_o[N][top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)] = tl_t_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)];
	// Trace: design.sv:79800:3
	assign tl_u_o[N][top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)] = tl_t_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)];
	// Trace: design.sv:79801:3
	assign tl_u_o[N][top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))] = tl_t_o[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))];
	// Trace: design.sv:79802:3
	assign tl_u_o[N][53-:32] = tl_t_o[53-:32];
	// Trace: design.sv:79803:3
	assign tl_u_o[N][21-:21] = tl_t_o[21-:21];
	// Trace: design.sv:79804:3
	tlul_err_resp err_resp(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(tl_u_o[N]),
		.tl_h_o(tl_u_i[N])
	);
	initial _sv2v_0 = 0;
endmodule
module tlul_cmd_intg_gen (
	tl_i,
	tl_o
);
	reg _sv2v_0;
	// removed import tlul_pkg::*;
	// Trace: design.sv:79823:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:79824:3
	output reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_o;
	// Trace: design.sv:79827:3
	// removed localparam type tlul_pkg_tl_h2d_cmd_intg_t
	wire [(37 + top_pkg_TL_DBW) - 1:0] cmd;
	// Trace: design.sv:79828:3
	function automatic [(37 + top_pkg_TL_DBW) - 1:0] tlul_pkg_extract_h2d_cmd_intg;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:145:61
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:146:5
		reg [(37 + top_pkg_TL_DBW) - 1:0] payload;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:147:5
		reg unused_tlul;
		begin
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:148:5
			unused_tlul = ^tl;
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:149:5
			payload[top_pkg_TL_AW + (top_pkg_TL_DBW + 2)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) >= (3 + (top_pkg_TL_DBW + 0)) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) - (3 + (top_pkg_TL_DBW + 0))) + 1 : ((3 + (top_pkg_TL_DBW + 0)) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) + 1)] = tl[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:150:5
			payload[top_pkg_TL_DBW + 2-:((top_pkg_TL_DBW + 2) >= (top_pkg_TL_DBW + 0) ? ((top_pkg_TL_DBW + 2) - (top_pkg_TL_DBW + 0)) + 1 : ((top_pkg_TL_DBW + 0) - (top_pkg_TL_DBW + 2)) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:151:5
			payload[top_pkg_TL_DBW - 1-:top_pkg_TL_DBW] = tl[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:152:5
			payload[2 + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))-:((34 + (top_pkg_TL_DBW + 2)) >= (35 + (top_pkg_TL_DBW + 0)) ? ((2 + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) - (top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0)))) + 1 : ((top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0))) - (2 + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2)))) + 1)] = tl[16-:2];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:153:5
			tlul_pkg_extract_h2d_cmd_intg = payload;
		end
	endfunction
	assign cmd = tlul_pkg_extract_h2d_cmd_intg(tl_i);
	// Trace: design.sv:79829:3
	localparam signed [31:0] tlul_pkg_H2DCmdMaxWidth = 57;
	wire [56:0] unused_cmd_payload;
	// Trace: design.sv:79831:3
	wire [6:0] cmd_intg;
	// Trace: design.sv:79832:3
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	prim_secded_64_57_enc u_cmd_gen(
		.in(sv2v_cast_57(cmd)),
		.out({cmd_intg, unused_cmd_payload})
	);
	// Trace: design.sv:79837:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:79838:5
		tl_o = tl_i;
		// Trace: design.sv:79839:5
		tl_o[14-:7] = cmd_intg;
	end
	// Trace: design.sv:79842:3
	wire unused_tl;
	// Trace: design.sv:79843:3
	assign unused_tl = ^tl_i;
	initial _sv2v_0 = 0;
endmodule
module tlul_cmd_intg_chk (
	tl_i,
	err_o
);
	// removed import tlul_pkg::*;
	// Trace: design.sv:79860:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:79863:3
	output wire err_o;
	// Trace: design.sv:79866:3
	wire [1:0] err;
	// Trace: design.sv:79867:3
	// removed localparam type tlul_pkg_tl_h2d_cmd_intg_t
	wire [(37 + top_pkg_TL_DBW) - 1:0] cmd;
	// Trace: design.sv:79868:3
	function automatic [(37 + top_pkg_TL_DBW) - 1:0] tlul_pkg_extract_h2d_cmd_intg;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:145:61
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:146:5
		reg [(37 + top_pkg_TL_DBW) - 1:0] payload;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:147:5
		reg unused_tlul;
		begin
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:148:5
			unused_tlul = ^tl;
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:149:5
			payload[top_pkg_TL_AW + (top_pkg_TL_DBW + 2)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) >= (3 + (top_pkg_TL_DBW + 0)) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) - (3 + (top_pkg_TL_DBW + 0))) + 1 : ((3 + (top_pkg_TL_DBW + 0)) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) + 1)] = tl[top_pkg_TL_AW + (top_pkg_TL_DBW + 53)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) >= (top_pkg_TL_DBW + 54) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (top_pkg_TL_DBW + 54)) + 1 : ((top_pkg_TL_DBW + 54) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) + 1)];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:150:5
			payload[top_pkg_TL_DBW + 2-:((top_pkg_TL_DBW + 2) >= (top_pkg_TL_DBW + 0) ? ((top_pkg_TL_DBW + 2) - (top_pkg_TL_DBW + 0)) + 1 : ((top_pkg_TL_DBW + 0) - (top_pkg_TL_DBW + 2)) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:151:5
			payload[top_pkg_TL_DBW - 1-:top_pkg_TL_DBW] = tl[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:152:5
			payload[2 + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))-:((34 + (top_pkg_TL_DBW + 2)) >= (35 + (top_pkg_TL_DBW + 0)) ? ((2 + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) - (top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0)))) + 1 : ((top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0))) - (2 + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2)))) + 1)] = tl[16-:2];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:153:5
			tlul_pkg_extract_h2d_cmd_intg = payload;
		end
	endfunction
	assign cmd = tlul_pkg_extract_h2d_cmd_intg(tl_i);
	// Trace: design.sv:79870:3
	localparam signed [31:0] tlul_pkg_H2DCmdMaxWidth = 57;
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	prim_secded_64_57_dec u_chk(
		.in({tl_i[14-:7], sv2v_cast_57(cmd)}),
		.d_o(),
		.syndrome_o(),
		.err_o(err)
	);
	// Trace: design.sv:79879:3
	assign err_o = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] & |err;
	// Trace: design.sv:79881:3
	wire unused_tl;
	// Trace: design.sv:79882:3
	assign unused_tl = |tl_i;
endmodule
module tlul_rsp_intg_gen (
	tl_i,
	tl_o
);
	reg _sv2v_0;
	// removed import tlul_pkg::*;
	// Trace: design.sv:79898:13
	parameter [0:0] EnableRspIntgGen = 1'b1;
	// Trace: design.sv:79899:13
	parameter [0:0] EnableDataIntgGen = 1'b1;
	// Trace: design.sv:79902:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_d2h_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_i;
	// Trace: design.sv:79903:3
	output reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:79906:3
	wire [6:0] rsp_intg;
	// Trace: design.sv:79907:3
	localparam signed [31:0] tlul_pkg_D2HRspMaxWidth = 57;
	// removed localparam type tlul_pkg_tl_d2h_rsp_intg_t
	function automatic [(3 + top_pkg_TL_SZW) + 0:0] tlul_pkg_extract_d2h_rsp_intg;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:157:61
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:158:5
		reg [(3 + top_pkg_TL_SZW) + 0:0] payload;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:159:5
		reg unused_tlul;
		begin
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:160:5
			unused_tlul = ^tl;
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:161:5
			payload[3 + (top_pkg_TL_SZW + 0)-:((3 + (top_pkg_TL_SZW + 0)) >= (top_pkg_TL_SZW + 1) ? ((3 + (top_pkg_TL_SZW + 0)) - (top_pkg_TL_SZW + 1)) + 1 : ((top_pkg_TL_SZW + 1) - (3 + (top_pkg_TL_SZW + 0))) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:162:5
			payload[top_pkg_TL_SZW + 0-:((top_pkg_TL_SZW + 0) >= 1 ? top_pkg_TL_SZW + 0 : 2 - (top_pkg_TL_SZW + 0))] = tl[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:164:5
			payload[0] = tl[1];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:165:5
			tlul_pkg_extract_d2h_rsp_intg = payload;
		end
	endfunction
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	generate
		if (EnableRspIntgGen) begin : gen_rsp_intg
			// Trace: design.sv:79908:5
			wire [(3 + top_pkg_TL_SZW) + 0:0] rsp;
			// Trace: design.sv:79909:5
			wire [56:0] unused_payload;
			// Trace: design.sv:79911:5
			assign rsp = tlul_pkg_extract_d2h_rsp_intg(tl_i);
			// Trace: design.sv:79913:5
			prim_secded_64_57_enc u_rsp_gen(
				.in(sv2v_cast_57(rsp)),
				.out({rsp_intg, unused_payload})
			);
		end
		else begin : gen_passthrough_rsp_intg
			// Trace: design.sv:79918:5
			assign rsp_intg = tl_i[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 14)-:7];
		end
	endgenerate
	// Trace: design.sv:79921:3
	wire [6:0] data_intg;
	// Trace: design.sv:79922:3
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 57;
	generate
		if (EnableDataIntgGen) begin : gen_data_intg
			// Trace: design.sv:79923:5
			wire [56:0] unused_data;
			// Trace: design.sv:79925:5
			prim_secded_64_57_enc u_data_gen(
				.in(sv2v_cast_57(tl_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)])),
				.out({data_intg, unused_data})
			);
		end
		else begin : gen_passthrough_data_intg
			// Trace: design.sv:79930:5
			assign data_intg = tl_i[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 7)-:tlul_pkg_DataIntgWidth];
		end
	endgenerate
	// Trace: design.sv:79933:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:79934:5
		tl_o = tl_i;
		// Trace: design.sv:79935:5
		tl_o[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 14)-:7] = rsp_intg;
		// Trace: design.sv:79936:5
		tl_o[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 7)-:tlul_pkg_DataIntgWidth] = data_intg;
	end
	// Trace: design.sv:79939:3
	wire unused_tl;
	// Trace: design.sv:79940:3
	assign unused_tl = ^tl_i;
	initial _sv2v_0 = 0;
endmodule
module tlul_rsp_intg_chk (
	tl_i,
	err_o
);
	// removed import tlul_pkg::*;
	// Trace: design.sv:79959:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_d2h_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_i;
	// Trace: design.sv:79962:3
	output wire err_o;
	// Trace: design.sv:79965:3
	wire [1:0] err;
	// Trace: design.sv:79966:3
	// removed localparam type tlul_pkg_tl_d2h_rsp_intg_t
	wire [(3 + top_pkg_TL_SZW) + 0:0] rsp;
	// Trace: design.sv:79967:3
	function automatic [(3 + top_pkg_TL_SZW) + 0:0] tlul_pkg_extract_d2h_rsp_intg;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:157:61
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:158:5
		reg [(3 + top_pkg_TL_SZW) + 0:0] payload;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:159:5
		reg unused_tlul;
		begin
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:160:5
			unused_tlul = ^tl;
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:161:5
			payload[3 + (top_pkg_TL_SZW + 0)-:((3 + (top_pkg_TL_SZW + 0)) >= (top_pkg_TL_SZW + 1) ? ((3 + (top_pkg_TL_SZW + 0)) - (top_pkg_TL_SZW + 1)) + 1 : ((top_pkg_TL_SZW + 1) - (3 + (top_pkg_TL_SZW + 0))) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:162:5
			payload[top_pkg_TL_SZW + 0-:((top_pkg_TL_SZW + 0) >= 1 ? top_pkg_TL_SZW + 0 : 2 - (top_pkg_TL_SZW + 0))] = tl[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:164:5
			payload[0] = tl[1];
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:165:5
			tlul_pkg_extract_d2h_rsp_intg = payload;
		end
	endfunction
	assign rsp = tlul_pkg_extract_d2h_rsp_intg(tl_i);
	// Trace: design.sv:79969:3
	localparam signed [31:0] tlul_pkg_D2HRspMaxWidth = 57;
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	prim_secded_64_57_dec u_chk(
		.in({tl_i[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 14)-:7], sv2v_cast_57(rsp)}),
		.d_o(),
		.syndrome_o(),
		.err_o(err)
	);
	// Trace: design.sv:79981:3
	assign err_o = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & |err;
	// Trace: design.sv:79983:3
	wire unused_tl;
	// Trace: design.sv:79984:3
	assign unused_tl = |tl_i;
endmodule
// removed package "soc_ctrl_reg_pkg"
module soc_ctrl_reg_top_28969 (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	reg2hw,
	hw2reg,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:80097:20
	// removed localparam type reg_req_t
	// Trace: design.sv:80098:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:80099:15
	parameter signed [31:0] AW = 5;
	// Trace: design.sv:80101:5
	input clk_i;
	// Trace: design.sv:80102:5
	input rst_ni;
	// Trace: design.sv:80103:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:80104:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:80106:5
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_boot_address_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_boot_exit_loop_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_boot_select_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_enable_spi_sel_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_exit_valid_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_exit_value_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_use_spimemio_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_t
	output wire [68:0] reg2hw;
	// Trace: design.sv:80107:5
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_hw2reg_boot_exit_loop_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_hw2reg_boot_select_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_hw2reg_use_spimemio_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_hw2reg_t
	input wire [5:0] hw2reg;
	// Trace: design.sv:80111:5
	input devmode_i;
	// Trace: design.sv:80114:3
	// removed import soc_ctrl_reg_pkg::*;
	// Trace: design.sv:80116:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:80117:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:80120:3
	wire reg_we;
	// Trace: design.sv:80121:3
	wire reg_re;
	// Trace: design.sv:80122:3
	wire [AW - 1:0] reg_addr;
	// Trace: design.sv:80123:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:80124:3
	wire [3:0] reg_be;
	// Trace: design.sv:80125:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:80126:3
	wire reg_error;
	// Trace: design.sv:80128:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:80130:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:80133:3
	wire [69:0] reg_intf_req;
	// Trace: design.sv:80134:3
	wire [33:0] reg_intf_rsp;
	// Trace: design.sv:80137:3
	assign reg_intf_req = reg_req_i;
	// Trace: design.sv:80138:3
	assign reg_rsp_o = reg_intf_rsp;
	// Trace: design.sv:80141:3
	assign reg_we = reg_intf_req[69] & reg_intf_req[68];
	// Trace: design.sv:80142:3
	assign reg_re = reg_intf_req[69] & ~reg_intf_req[68];
	// Trace: design.sv:80143:3
	assign reg_addr = reg_intf_req[63-:32];
	// Trace: design.sv:80144:3
	assign reg_wdata = reg_intf_req[31-:32];
	// Trace: design.sv:80145:3
	assign reg_be = reg_intf_req[67-:4];
	// Trace: design.sv:80146:3
	assign reg_intf_rsp[31-:32] = reg_rdata;
	// Trace: design.sv:80147:3
	assign reg_intf_rsp[33] = reg_error;
	// Trace: design.sv:80148:3
	assign reg_intf_rsp[32] = 1'b1;
	// Trace: design.sv:80150:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:80151:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:80157:3
	wire exit_valid_qs;
	// Trace: design.sv:80158:3
	wire exit_valid_wd;
	// Trace: design.sv:80159:3
	wire exit_valid_we;
	// Trace: design.sv:80160:3
	wire [31:0] exit_value_qs;
	// Trace: design.sv:80161:3
	wire [31:0] exit_value_wd;
	// Trace: design.sv:80162:3
	wire exit_value_we;
	// Trace: design.sv:80163:3
	wire boot_select_qs;
	// Trace: design.sv:80164:3
	wire boot_exit_loop_qs;
	// Trace: design.sv:80165:3
	wire boot_exit_loop_wd;
	// Trace: design.sv:80166:3
	wire boot_exit_loop_we;
	// Trace: design.sv:80167:3
	wire [31:0] boot_address_qs;
	// Trace: design.sv:80168:3
	wire [31:0] boot_address_wd;
	// Trace: design.sv:80169:3
	wire boot_address_we;
	// Trace: design.sv:80170:3
	wire use_spimemio_qs;
	// Trace: design.sv:80171:3
	wire use_spimemio_wd;
	// Trace: design.sv:80172:3
	wire use_spimemio_we;
	// Trace: design.sv:80173:3
	wire enable_spi_sel_qs;
	// Trace: design.sv:80174:3
	wire enable_spi_sel_wd;
	// Trace: design.sv:80175:3
	wire enable_spi_sel_we;
	// Trace: design.sv:80176:3
	wire [31:0] system_frequency_hz_qs;
	// Trace: design.sv:80177:3
	wire [31:0] system_frequency_hz_wd;
	// Trace: design.sv:80178:3
	wire system_frequency_hz_we;
	// Trace: design.sv:80183:3
	localparam signed [31:0] sv2v_uu_u_exit_valid_DW = 1;
	// removed localparam type sv2v_uu_u_exit_valid_d
	localparam [0:0] sv2v_uu_u_exit_valid_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_exit_valid(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(exit_valid_we),
		.wd(exit_valid_wd),
		.de(1'b0),
		.d(sv2v_uu_u_exit_valid_ext_d_0),
		.qe(),
		.q(reg2hw[68]),
		.qs(exit_valid_qs)
	);
	// Trace: design.sv:80210:3
	localparam signed [31:0] sv2v_uu_u_exit_value_DW = 32;
	// removed localparam type sv2v_uu_u_exit_value_d
	localparam [31:0] sv2v_uu_u_exit_value_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_exit_value(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(exit_value_we),
		.wd(exit_value_wd),
		.de(1'b0),
		.d(sv2v_uu_u_exit_value_ext_d_0),
		.qe(),
		.q(reg2hw[67-:32]),
		.qs(exit_value_qs)
	);
	// Trace: design.sv:80237:3
	localparam signed [31:0] sv2v_uu_u_boot_select_DW = 1;
	// removed localparam type sv2v_uu_u_boot_select_wd
	localparam [0:0] sv2v_uu_u_boot_select_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_boot_select(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_boot_select_ext_wd_0),
		.de(hw2reg[4]),
		.d(hw2reg[5]),
		.qe(),
		.q(reg2hw[35]),
		.qs(boot_select_qs)
	);
	// Trace: design.sv:80263:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_boot_exit_loop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(boot_exit_loop_we),
		.wd(boot_exit_loop_wd),
		.de(hw2reg[2]),
		.d(hw2reg[3]),
		.qe(),
		.q(reg2hw[34]),
		.qs(boot_exit_loop_qs)
	);
	// Trace: design.sv:80290:3
	localparam signed [31:0] sv2v_uu_u_boot_address_DW = 32;
	// removed localparam type sv2v_uu_u_boot_address_d
	localparam [31:0] sv2v_uu_u_boot_address_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000180)
	) u_boot_address(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(boot_address_we),
		.wd(boot_address_wd),
		.de(1'b0),
		.d(sv2v_uu_u_boot_address_ext_d_0),
		.qe(),
		.q(reg2hw[33-:32]),
		.qs(boot_address_qs)
	);
	// Trace: design.sv:80317:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h1)
	) u_use_spimemio(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(use_spimemio_we),
		.wd(use_spimemio_wd),
		.de(hw2reg[0]),
		.d(hw2reg[1]),
		.qe(),
		.q(reg2hw[1]),
		.qs(use_spimemio_qs)
	);
	// Trace: design.sv:80344:3
	localparam signed [31:0] sv2v_uu_u_enable_spi_sel_DW = 1;
	// removed localparam type sv2v_uu_u_enable_spi_sel_d
	localparam [0:0] sv2v_uu_u_enable_spi_sel_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_enable_spi_sel(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(enable_spi_sel_we),
		.wd(enable_spi_sel_wd),
		.de(1'b0),
		.d(sv2v_uu_u_enable_spi_sel_ext_d_0),
		.qe(),
		.q(reg2hw[-0]),
		.qs(enable_spi_sel_qs)
	);
	// Trace: design.sv:80371:3
	localparam signed [31:0] sv2v_uu_u_system_frequency_hz_DW = 32;
	// removed localparam type sv2v_uu_u_system_frequency_hz_d
	localparam [31:0] sv2v_uu_u_system_frequency_hz_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000001)
	) u_system_frequency_hz(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(system_frequency_hz_we),
		.wd(system_frequency_hz_wd),
		.de(1'b0),
		.d(sv2v_uu_u_system_frequency_hz_ext_d_0),
		.qe(),
		.q(),
		.qs(system_frequency_hz_qs)
	);
	// Trace: design.sv:80398:3
	reg [7:0] addr_hit;
	// Trace: design.sv:80399:3
	localparam signed [31:0] soc_ctrl_reg_pkg_BlockAw = 5;
	localparam [4:0] soc_ctrl_reg_pkg_SOC_CTRL_BOOT_ADDRESS_OFFSET = 5'h10;
	localparam [4:0] soc_ctrl_reg_pkg_SOC_CTRL_BOOT_EXIT_LOOP_OFFSET = 5'h0c;
	localparam [4:0] soc_ctrl_reg_pkg_SOC_CTRL_BOOT_SELECT_OFFSET = 5'h08;
	localparam [4:0] soc_ctrl_reg_pkg_SOC_CTRL_ENABLE_SPI_SEL_OFFSET = 5'h18;
	localparam [4:0] soc_ctrl_reg_pkg_SOC_CTRL_EXIT_VALID_OFFSET = 5'h00;
	localparam [4:0] soc_ctrl_reg_pkg_SOC_CTRL_EXIT_VALUE_OFFSET = 5'h04;
	localparam [4:0] soc_ctrl_reg_pkg_SOC_CTRL_SYSTEM_FREQUENCY_HZ_OFFSET = 5'h1c;
	localparam [4:0] soc_ctrl_reg_pkg_SOC_CTRL_USE_SPIMEMIO_OFFSET = 5'h14;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:80400:5
		addr_hit = 1'sb0;
		// Trace: design.sv:80401:5
		addr_hit[0] = reg_addr == soc_ctrl_reg_pkg_SOC_CTRL_EXIT_VALID_OFFSET;
		// Trace: design.sv:80402:5
		addr_hit[1] = reg_addr == soc_ctrl_reg_pkg_SOC_CTRL_EXIT_VALUE_OFFSET;
		// Trace: design.sv:80403:5
		addr_hit[2] = reg_addr == soc_ctrl_reg_pkg_SOC_CTRL_BOOT_SELECT_OFFSET;
		// Trace: design.sv:80404:5
		addr_hit[3] = reg_addr == soc_ctrl_reg_pkg_SOC_CTRL_BOOT_EXIT_LOOP_OFFSET;
		// Trace: design.sv:80405:5
		addr_hit[4] = reg_addr == soc_ctrl_reg_pkg_SOC_CTRL_BOOT_ADDRESS_OFFSET;
		// Trace: design.sv:80406:5
		addr_hit[5] = reg_addr == soc_ctrl_reg_pkg_SOC_CTRL_USE_SPIMEMIO_OFFSET;
		// Trace: design.sv:80407:5
		addr_hit[6] = reg_addr == soc_ctrl_reg_pkg_SOC_CTRL_ENABLE_SPI_SEL_OFFSET;
		// Trace: design.sv:80408:5
		addr_hit[7] = reg_addr == soc_ctrl_reg_pkg_SOC_CTRL_SYSTEM_FREQUENCY_HZ_OFFSET;
	end
	// Trace: design.sv:80411:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:80414:3
	localparam [31:0] soc_ctrl_reg_pkg_SOC_CTRL_PERMIT = 32'b00011111000100011111000100011111;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:80415:5
		wr_err = reg_we & ((((((((addr_hit[0] & |(soc_ctrl_reg_pkg_SOC_CTRL_PERMIT[28+:4] & ~reg_be)) | (addr_hit[1] & |(soc_ctrl_reg_pkg_SOC_CTRL_PERMIT[24+:4] & ~reg_be))) | (addr_hit[2] & |(soc_ctrl_reg_pkg_SOC_CTRL_PERMIT[20+:4] & ~reg_be))) | (addr_hit[3] & |(soc_ctrl_reg_pkg_SOC_CTRL_PERMIT[16+:4] & ~reg_be))) | (addr_hit[4] & |(soc_ctrl_reg_pkg_SOC_CTRL_PERMIT[12+:4] & ~reg_be))) | (addr_hit[5] & |(soc_ctrl_reg_pkg_SOC_CTRL_PERMIT[8+:4] & ~reg_be))) | (addr_hit[6] & |(soc_ctrl_reg_pkg_SOC_CTRL_PERMIT[4+:4] & ~reg_be))) | (addr_hit[7] & |(soc_ctrl_reg_pkg_SOC_CTRL_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:80426:3
	assign exit_valid_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:80427:3
	assign exit_valid_wd = reg_wdata[0];
	// Trace: design.sv:80429:3
	assign exit_value_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:80430:3
	assign exit_value_wd = reg_wdata[31:0];
	// Trace: design.sv:80432:3
	assign boot_exit_loop_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:80433:3
	assign boot_exit_loop_wd = reg_wdata[0];
	// Trace: design.sv:80435:3
	assign boot_address_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:80436:3
	assign boot_address_wd = reg_wdata[31:0];
	// Trace: design.sv:80438:3
	assign use_spimemio_we = (addr_hit[5] & reg_we) & !reg_error;
	// Trace: design.sv:80439:3
	assign use_spimemio_wd = reg_wdata[0];
	// Trace: design.sv:80441:3
	assign enable_spi_sel_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:80442:3
	assign enable_spi_sel_wd = reg_wdata[0];
	// Trace: design.sv:80444:3
	assign system_frequency_hz_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:80445:3
	assign system_frequency_hz_wd = reg_wdata[31:0];
	// Trace: design.sv:80448:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:80449:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:80450:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]:
				// Trace: design.sv:80452:9
				reg_rdata_next[0] = exit_valid_qs;
			addr_hit[1]:
				// Trace: design.sv:80456:9
				reg_rdata_next[31:0] = exit_value_qs;
			addr_hit[2]:
				// Trace: design.sv:80460:9
				reg_rdata_next[0] = boot_select_qs;
			addr_hit[3]:
				// Trace: design.sv:80464:9
				reg_rdata_next[0] = boot_exit_loop_qs;
			addr_hit[4]:
				// Trace: design.sv:80468:9
				reg_rdata_next[31:0] = boot_address_qs;
			addr_hit[5]:
				// Trace: design.sv:80472:9
				reg_rdata_next[0] = use_spimemio_qs;
			addr_hit[6]:
				// Trace: design.sv:80476:9
				reg_rdata_next[0] = enable_spi_sel_qs;
			addr_hit[7]:
				// Trace: design.sv:80480:9
				reg_rdata_next[31:0] = system_frequency_hz_qs;
			default:
				// Trace: design.sv:80484:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:80493:3
	wire unused_wdata;
	// Trace: design.sv:80494:3
	wire unused_be;
	// Trace: design.sv:80495:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:80496:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module soc_ctrl_E136A (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	boot_select_i,
	execute_from_flash_i,
	use_spimemio_o,
	exit_valid_o,
	exit_value_o
);
	// Trace: design.sv:80509:20
	// removed localparam type reg_req_t
	// Trace: design.sv:80510:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:80512:5
	input wire clk_i;
	// Trace: design.sv:80513:5
	input wire rst_ni;
	// Trace: design.sv:80516:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:80517:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:80519:5
	input wire boot_select_i;
	// Trace: design.sv:80520:5
	input wire execute_from_flash_i;
	// Trace: design.sv:80521:5
	output wire use_spimemio_o;
	// Trace: design.sv:80523:5
	output wire exit_valid_o;
	// Trace: design.sv:80524:5
	output wire [31:0] exit_value_o;
	// Trace: design.sv:80527:3
	// removed import soc_ctrl_reg_pkg::*;
	// Trace: design.sv:80529:3
	wire enable_spi_sel;
	// Trace: design.sv:80531:3
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_boot_address_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_boot_exit_loop_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_boot_select_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_enable_spi_sel_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_exit_valid_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_exit_value_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_use_spimemio_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_reg2hw_t
	wire [68:0] reg2hw;
	// Trace: design.sv:80532:3
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_hw2reg_boot_exit_loop_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_hw2reg_boot_select_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_hw2reg_use_spimemio_reg_t
	// removed localparam type soc_ctrl_reg_pkg_soc_ctrl_hw2reg_t
	wire [5:0] hw2reg;
	// Trace: design.sv:80547:3
	assign hw2reg[3] = 1'b0;
	// Trace: design.sv:80548:3
	assign hw2reg[2] = 1'b0;
	// Trace: design.sv:80551:3
	assign hw2reg[4] = 1'b1;
	// Trace: design.sv:80552:3
	assign hw2reg[5] = boot_select_i;
	// Trace: design.sv:80554:3
	assign hw2reg[0] = ~enable_spi_sel;
	// Trace: design.sv:80555:3
	assign hw2reg[1] = execute_from_flash_i;
	// Trace: design.sv:80557:3
	soc_ctrl_reg_top_28969 soc_ctrl_reg_top_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(reg_req_i),
		.reg_rsp_o(reg_rsp_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:80570:3
	assign exit_valid_o = reg2hw[68];
	// Trace: design.sv:80571:3
	assign exit_value_o = reg2hw[67-:32];
	// Trace: design.sv:80572:3
	assign use_spimemio_o = reg2hw[1];
	// Trace: design.sv:80573:3
	assign enable_spi_sel = reg2hw[-0];
endmodule
// removed package "fast_intr_ctrl_reg_pkg"
module fast_intr_ctrl_reg_top_F39E6 (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	reg2hw,
	hw2reg,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:80645:20
	// removed localparam type reg_req_t
	// Trace: design.sv:80646:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:80647:15
	parameter signed [31:0] AW = 3;
	// Trace: design.sv:80649:5
	input clk_i;
	// Trace: design.sv:80650:5
	input rst_ni;
	// Trace: design.sv:80651:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:80652:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:80654:5
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_reg2hw_fast_intr_clear_reg_t
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_reg2hw_fast_intr_pending_reg_t
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_reg2hw_t
	output wire [31:0] reg2hw;
	// Trace: design.sv:80655:5
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_hw2reg_fast_intr_clear_reg_t
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_hw2reg_fast_intr_pending_reg_t
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_hw2reg_t
	input wire [33:0] hw2reg;
	// Trace: design.sv:80659:5
	input devmode_i;
	// Trace: design.sv:80662:3
	// removed import fast_intr_ctrl_reg_pkg::*;
	// Trace: design.sv:80664:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:80665:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:80668:3
	wire reg_we;
	// Trace: design.sv:80669:3
	wire reg_re;
	// Trace: design.sv:80670:3
	wire [AW - 1:0] reg_addr;
	// Trace: design.sv:80671:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:80672:3
	wire [3:0] reg_be;
	// Trace: design.sv:80673:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:80674:3
	wire reg_error;
	// Trace: design.sv:80676:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:80678:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:80681:3
	wire [69:0] reg_intf_req;
	// Trace: design.sv:80682:3
	wire [33:0] reg_intf_rsp;
	// Trace: design.sv:80685:3
	assign reg_intf_req = reg_req_i;
	// Trace: design.sv:80686:3
	assign reg_rsp_o = reg_intf_rsp;
	// Trace: design.sv:80689:3
	assign reg_we = reg_intf_req[69] & reg_intf_req[68];
	// Trace: design.sv:80690:3
	assign reg_re = reg_intf_req[69] & ~reg_intf_req[68];
	// Trace: design.sv:80691:3
	assign reg_addr = reg_intf_req[63-:32];
	// Trace: design.sv:80692:3
	assign reg_wdata = reg_intf_req[31-:32];
	// Trace: design.sv:80693:3
	assign reg_be = reg_intf_req[67-:4];
	// Trace: design.sv:80694:3
	assign reg_intf_rsp[31-:32] = reg_rdata;
	// Trace: design.sv:80695:3
	assign reg_intf_rsp[33] = reg_error;
	// Trace: design.sv:80696:3
	assign reg_intf_rsp[32] = 1'b1;
	// Trace: design.sv:80698:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:80699:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:80705:3
	wire [15:0] fast_intr_pending_qs;
	// Trace: design.sv:80706:3
	wire [15:0] fast_intr_clear_qs;
	// Trace: design.sv:80707:3
	wire [15:0] fast_intr_clear_wd;
	// Trace: design.sv:80708:3
	wire fast_intr_clear_we;
	// Trace: design.sv:80713:3
	localparam signed [31:0] sv2v_uu_u_fast_intr_pending_DW = 16;
	// removed localparam type sv2v_uu_u_fast_intr_pending_wd
	localparam [15:0] sv2v_uu_u_fast_intr_pending_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RO"),
		.RESVAL(16'h0000)
	) u_fast_intr_pending(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_fast_intr_pending_ext_wd_0),
		.de(hw2reg[17]),
		.d(hw2reg[33-:16]),
		.qe(),
		.q(reg2hw[31-:16]),
		.qs(fast_intr_pending_qs)
	);
	// Trace: design.sv:80739:3
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_fast_intr_clear(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fast_intr_clear_we),
		.wd(fast_intr_clear_wd),
		.de(hw2reg[0]),
		.d(hw2reg[16-:16]),
		.qe(),
		.q(reg2hw[15-:16]),
		.qs(fast_intr_clear_qs)
	);
	// Trace: design.sv:80766:3
	reg [1:0] addr_hit;
	// Trace: design.sv:80767:3
	localparam signed [31:0] fast_intr_ctrl_reg_pkg_BlockAw = 3;
	localparam [2:0] fast_intr_ctrl_reg_pkg_FAST_INTR_CTRL_FAST_INTR_CLEAR_OFFSET = 3'h4;
	localparam [2:0] fast_intr_ctrl_reg_pkg_FAST_INTR_CTRL_FAST_INTR_PENDING_OFFSET = 3'h0;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:80768:5
		addr_hit = 1'sb0;
		// Trace: design.sv:80769:5
		addr_hit[0] = reg_addr == fast_intr_ctrl_reg_pkg_FAST_INTR_CTRL_FAST_INTR_PENDING_OFFSET;
		// Trace: design.sv:80770:5
		addr_hit[1] = reg_addr == fast_intr_ctrl_reg_pkg_FAST_INTR_CTRL_FAST_INTR_CLEAR_OFFSET;
	end
	// Trace: design.sv:80773:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:80776:3
	localparam [7:0] fast_intr_ctrl_reg_pkg_FAST_INTR_CTRL_PERMIT = 8'b00110011;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:80777:5
		wr_err = reg_we & ((addr_hit[0] & |(fast_intr_ctrl_reg_pkg_FAST_INTR_CTRL_PERMIT[4+:4] & ~reg_be)) | (addr_hit[1] & |(fast_intr_ctrl_reg_pkg_FAST_INTR_CTRL_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:80782:3
	assign fast_intr_clear_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:80783:3
	assign fast_intr_clear_wd = reg_wdata[15:0];
	// Trace: design.sv:80786:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:80787:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:80788:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]:
				// Trace: design.sv:80790:9
				reg_rdata_next[15:0] = fast_intr_pending_qs;
			addr_hit[1]:
				// Trace: design.sv:80794:9
				reg_rdata_next[15:0] = fast_intr_clear_qs;
			default:
				// Trace: design.sv:80798:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:80807:3
	wire unused_wdata;
	// Trace: design.sv:80808:3
	wire unused_be;
	// Trace: design.sv:80809:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:80810:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module fast_intr_ctrl_65415 (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	fast_intr_i,
	fast_intr_o
);
	reg _sv2v_0;
	// Trace: design.sv:80823:20
	// removed localparam type reg_req_t
	// Trace: design.sv:80824:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:80826:5
	input wire clk_i;
	// Trace: design.sv:80827:5
	input wire rst_ni;
	// Trace: design.sv:80830:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:80831:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:80833:5
	input wire [14:0] fast_intr_i;
	// Trace: design.sv:80834:5
	output wire [14:0] fast_intr_o;
	// Trace: design.sv:80837:3
	// removed import fast_intr_ctrl_reg_pkg::*;
	// Trace: design.sv:80839:3
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_reg2hw_fast_intr_clear_reg_t
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_reg2hw_fast_intr_pending_reg_t
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_reg2hw_t
	wire [31:0] reg2hw;
	// Trace: design.sv:80840:3
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_hw2reg_fast_intr_clear_reg_t
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_hw2reg_fast_intr_pending_reg_t
	// removed localparam type fast_intr_ctrl_reg_pkg_fast_intr_ctrl_hw2reg_t
	reg [33:0] hw2reg;
	// Trace: design.sv:80842:3
	reg [14:0] fast_intr_pending_de;
	// Trace: design.sv:80843:3
	reg [14:0] fast_intr_clear_de;
	// Trace: design.sv:80845:3
	fast_intr_ctrl_reg_top_F39E6 fast_intr_ctrl_reg_top_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(reg_req_i),
		.reg_rsp_o(reg_rsp_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:80858:3
	genvar _gv_i_91;
	generate
		for (_gv_i_91 = 0; _gv_i_91 < 15; _gv_i_91 = _gv_i_91 + 1) begin : gen_fast_interrupt
			localparam i = _gv_i_91;
			// Trace: design.sv:80860:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: design.sv:80861:7
				if (reg2hw[0 + i]) begin
					// Trace: design.sv:80862:9
					fast_intr_pending_de[i] = 1'b1;
					// Trace: design.sv:80863:9
					hw2reg[18 + i] = 1'b0;
					// Trace: design.sv:80864:9
					fast_intr_clear_de[i] = 1'b1;
					// Trace: design.sv:80865:9
					hw2reg[1 + i] = 1'b0;
				end
				else
					// Trace: design.sv:80867:9
					if (fast_intr_i[i]) begin
						// Trace: design.sv:80868:11
						fast_intr_pending_de[i] = 1'b1;
						// Trace: design.sv:80869:11
						hw2reg[18 + i] = 1'b1;
						// Trace: design.sv:80870:11
						fast_intr_clear_de[i] = 1'b0;
						// Trace: design.sv:80871:11
						hw2reg[1 + i] = 1'b0;
					end
					else begin
						// Trace: design.sv:80873:11
						fast_intr_pending_de[i] = 1'b0;
						// Trace: design.sv:80874:11
						hw2reg[18 + i] = 1'b0;
						// Trace: design.sv:80875:11
						fast_intr_clear_de[i] = 1'b0;
						// Trace: design.sv:80876:11
						hw2reg[1 + i] = 1'b0;
					end
			end
		end
	endgenerate
	// Trace: design.sv:80883:3
	wire [1:1] sv2v_tmp_99126;
	assign sv2v_tmp_99126 = 1'b0;
	always @(*) hw2reg[33] = sv2v_tmp_99126;
	// Trace: design.sv:80884:3
	wire [1:1] sv2v_tmp_005A1;
	assign sv2v_tmp_005A1 = 1'b0;
	always @(*) hw2reg[16] = sv2v_tmp_005A1;
	// Trace: design.sv:80885:3
	assign fast_intr_o = reg2hw[30:16];
	// Trace: design.sv:80886:3
	wire [1:1] sv2v_tmp_940FB;
	assign sv2v_tmp_940FB = |fast_intr_pending_de;
	always @(*) hw2reg[17] = sv2v_tmp_940FB;
	// Trace: design.sv:80887:3
	wire [1:1] sv2v_tmp_8ABF6;
	assign sv2v_tmp_8ABF6 = |fast_intr_clear_de;
	always @(*) hw2reg[0] = sv2v_tmp_8ABF6;
	initial _sv2v_0 = 0;
endmodule
module power_manager_reg_top_E039C (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	reg2hw,
	hw2reg,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:80900:18
	// removed localparam type reg_req_t
	// Trace: design.sv:80901:18
	// removed localparam type reg_rsp_t
	// Trace: design.sv:80902:13
	parameter signed [31:0] AW = 8;
	// Trace: design.sv:80904:3
	input wire clk_i;
	// Trace: design.sv:80905:3
	input wire rst_ni;
	// Trace: design.sv:80906:3
	input wire [69:0] reg_req_i;
	// Trace: design.sv:80907:3
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:80909:3
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_counters_stop_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_iso_off_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_iso_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_reset_assert_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_reset_deassert_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_switch_off_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_switch_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_wait_ack_switch_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_en_wait_for_intr_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_intr_state_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_iso_off_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_iso_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_reset_assert_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_reset_deassert_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_switch_off_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_switch_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_clk_gate_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_iso_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_reset_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_switch_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_wait_ack_switch_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_core_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_core_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_periph_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_ram_block_0_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_ram_block_1_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_clk_gate_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_iso_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_retentive_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_switch_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_wait_ack_switch_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_clk_gate_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_iso_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_retentive_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_switch_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_wait_ack_switch_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_restore_address_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_wakeup_state_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_t
	output wire [321:0] reg2hw;
	// Trace: design.sv:80910:3
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_iso_off_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_iso_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_reset_assert_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_reset_deassert_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_switch_off_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_switch_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_intr_state_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_monitor_power_gate_core_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_monitor_power_gate_periph_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_monitor_power_gate_ram_block_0_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_monitor_power_gate_ram_block_1_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_power_gate_core_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_power_gate_periph_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_power_gate_ram_block_0_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_power_gate_ram_block_1_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_t
	input wire [252:0] hw2reg;
	// Trace: design.sv:80914:3
	input devmode_i;
	// Trace: design.sv:80917:3
	// removed import power_manager_reg_pkg::*;
	// Trace: design.sv:80919:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:80920:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:80923:3
	wire reg_we;
	// Trace: design.sv:80924:3
	wire reg_re;
	// Trace: design.sv:80925:3
	wire [AW - 1:0] reg_addr;
	// Trace: design.sv:80926:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:80927:3
	wire [3:0] reg_be;
	// Trace: design.sv:80928:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:80929:3
	wire reg_error;
	// Trace: design.sv:80931:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:80933:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:80936:3
	wire [69:0] reg_intf_req;
	// Trace: design.sv:80937:3
	wire [33:0] reg_intf_rsp;
	// Trace: design.sv:80940:3
	assign reg_intf_req = reg_req_i;
	// Trace: design.sv:80941:3
	assign reg_rsp_o = reg_intf_rsp;
	// Trace: design.sv:80944:3
	assign reg_we = reg_intf_req[69] & reg_intf_req[68];
	// Trace: design.sv:80945:3
	assign reg_re = reg_intf_req[69] & ~reg_intf_req[68];
	// Trace: design.sv:80946:3
	assign reg_addr = reg_intf_req[63-:32];
	// Trace: design.sv:80947:3
	assign reg_wdata = reg_intf_req[31-:32];
	// Trace: design.sv:80948:3
	assign reg_be = reg_intf_req[67-:4];
	// Trace: design.sv:80949:3
	assign reg_intf_rsp[31-:32] = reg_rdata;
	// Trace: design.sv:80950:3
	assign reg_intf_rsp[33] = reg_error;
	// Trace: design.sv:80951:3
	assign reg_intf_rsp[32] = 1'b1;
	// Trace: design.sv:80953:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:80954:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:80960:3
	wire wakeup_state_qs;
	// Trace: design.sv:80961:3
	wire wakeup_state_wd;
	// Trace: design.sv:80962:3
	wire wakeup_state_we;
	// Trace: design.sv:80963:3
	wire [31:0] restore_address_qs;
	// Trace: design.sv:80964:3
	wire [31:0] restore_address_wd;
	// Trace: design.sv:80965:3
	wire restore_address_we;
	// Trace: design.sv:80966:3
	wire [31:0] en_wait_for_intr_qs;
	// Trace: design.sv:80967:3
	wire [31:0] en_wait_for_intr_wd;
	// Trace: design.sv:80968:3
	wire en_wait_for_intr_we;
	// Trace: design.sv:80969:3
	wire [31:0] intr_state_qs;
	// Trace: design.sv:80970:3
	wire [31:0] intr_state_wd;
	// Trace: design.sv:80971:3
	wire intr_state_we;
	// Trace: design.sv:80972:3
	wire power_gate_core_qs;
	// Trace: design.sv:80973:3
	wire power_gate_core_wd;
	// Trace: design.sv:80974:3
	wire power_gate_core_we;
	// Trace: design.sv:80975:3
	wire power_gate_core_ack_qs;
	// Trace: design.sv:80976:3
	wire [31:0] cpu_reset_assert_counter_qs;
	// Trace: design.sv:80977:3
	wire [31:0] cpu_reset_assert_counter_wd;
	// Trace: design.sv:80978:3
	wire cpu_reset_assert_counter_we;
	// Trace: design.sv:80979:3
	wire [31:0] cpu_reset_deassert_counter_qs;
	// Trace: design.sv:80980:3
	wire [31:0] cpu_reset_deassert_counter_wd;
	// Trace: design.sv:80981:3
	wire cpu_reset_deassert_counter_we;
	// Trace: design.sv:80982:3
	wire [31:0] cpu_switch_off_counter_qs;
	// Trace: design.sv:80983:3
	wire [31:0] cpu_switch_off_counter_wd;
	// Trace: design.sv:80984:3
	wire cpu_switch_off_counter_we;
	// Trace: design.sv:80985:3
	wire [31:0] cpu_switch_on_counter_qs;
	// Trace: design.sv:80986:3
	wire [31:0] cpu_switch_on_counter_wd;
	// Trace: design.sv:80987:3
	wire cpu_switch_on_counter_we;
	// Trace: design.sv:80988:3
	wire cpu_wait_ack_switch_on_counter_qs;
	// Trace: design.sv:80989:3
	wire cpu_wait_ack_switch_on_counter_wd;
	// Trace: design.sv:80990:3
	wire cpu_wait_ack_switch_on_counter_we;
	// Trace: design.sv:80991:3
	wire [31:0] cpu_iso_off_counter_qs;
	// Trace: design.sv:80992:3
	wire [31:0] cpu_iso_off_counter_wd;
	// Trace: design.sv:80993:3
	wire cpu_iso_off_counter_we;
	// Trace: design.sv:80994:3
	wire [31:0] cpu_iso_on_counter_qs;
	// Trace: design.sv:80995:3
	wire [31:0] cpu_iso_on_counter_wd;
	// Trace: design.sv:80996:3
	wire cpu_iso_on_counter_we;
	// Trace: design.sv:80997:3
	wire cpu_counters_stop_cpu_reset_assert_stop_bit_counter_qs;
	// Trace: design.sv:80998:3
	wire cpu_counters_stop_cpu_reset_assert_stop_bit_counter_wd;
	// Trace: design.sv:80999:3
	wire cpu_counters_stop_cpu_reset_assert_stop_bit_counter_we;
	// Trace: design.sv:81000:3
	wire cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_qs;
	// Trace: design.sv:81001:3
	wire cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_wd;
	// Trace: design.sv:81002:3
	wire cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_we;
	// Trace: design.sv:81003:3
	wire cpu_counters_stop_cpu_switch_off_stop_bit_counter_qs;
	// Trace: design.sv:81004:3
	wire cpu_counters_stop_cpu_switch_off_stop_bit_counter_wd;
	// Trace: design.sv:81005:3
	wire cpu_counters_stop_cpu_switch_off_stop_bit_counter_we;
	// Trace: design.sv:81006:3
	wire cpu_counters_stop_cpu_switch_on_stop_bit_counter_qs;
	// Trace: design.sv:81007:3
	wire cpu_counters_stop_cpu_switch_on_stop_bit_counter_wd;
	// Trace: design.sv:81008:3
	wire cpu_counters_stop_cpu_switch_on_stop_bit_counter_we;
	// Trace: design.sv:81009:3
	wire cpu_counters_stop_cpu_iso_off_stop_bit_counter_qs;
	// Trace: design.sv:81010:3
	wire cpu_counters_stop_cpu_iso_off_stop_bit_counter_wd;
	// Trace: design.sv:81011:3
	wire cpu_counters_stop_cpu_iso_off_stop_bit_counter_we;
	// Trace: design.sv:81012:3
	wire cpu_counters_stop_cpu_iso_on_stop_bit_counter_qs;
	// Trace: design.sv:81013:3
	wire cpu_counters_stop_cpu_iso_on_stop_bit_counter_wd;
	// Trace: design.sv:81014:3
	wire cpu_counters_stop_cpu_iso_on_stop_bit_counter_we;
	// Trace: design.sv:81015:3
	wire power_gate_periph_ack_qs;
	// Trace: design.sv:81016:3
	wire periph_reset_qs;
	// Trace: design.sv:81017:3
	wire periph_reset_wd;
	// Trace: design.sv:81018:3
	wire periph_reset_we;
	// Trace: design.sv:81019:3
	wire periph_switch_qs;
	// Trace: design.sv:81020:3
	wire periph_switch_wd;
	// Trace: design.sv:81021:3
	wire periph_switch_we;
	// Trace: design.sv:81022:3
	wire periph_wait_ack_switch_on_qs;
	// Trace: design.sv:81023:3
	wire periph_wait_ack_switch_on_wd;
	// Trace: design.sv:81024:3
	wire periph_wait_ack_switch_on_we;
	// Trace: design.sv:81025:3
	wire periph_iso_qs;
	// Trace: design.sv:81026:3
	wire periph_iso_wd;
	// Trace: design.sv:81027:3
	wire periph_iso_we;
	// Trace: design.sv:81028:3
	wire periph_clk_gate_qs;
	// Trace: design.sv:81029:3
	wire periph_clk_gate_wd;
	// Trace: design.sv:81030:3
	wire periph_clk_gate_we;
	// Trace: design.sv:81031:3
	wire ram_0_clk_gate_qs;
	// Trace: design.sv:81032:3
	wire ram_0_clk_gate_wd;
	// Trace: design.sv:81033:3
	wire ram_0_clk_gate_we;
	// Trace: design.sv:81034:3
	wire power_gate_ram_block_0_ack_qs;
	// Trace: design.sv:81035:3
	wire ram_0_switch_qs;
	// Trace: design.sv:81036:3
	wire ram_0_switch_wd;
	// Trace: design.sv:81037:3
	wire ram_0_switch_we;
	// Trace: design.sv:81038:3
	wire ram_0_wait_ack_switch_on_qs;
	// Trace: design.sv:81039:3
	wire ram_0_wait_ack_switch_on_wd;
	// Trace: design.sv:81040:3
	wire ram_0_wait_ack_switch_on_we;
	// Trace: design.sv:81041:3
	wire ram_0_iso_qs;
	// Trace: design.sv:81042:3
	wire ram_0_iso_wd;
	// Trace: design.sv:81043:3
	wire ram_0_iso_we;
	// Trace: design.sv:81044:3
	wire ram_0_retentive_qs;
	// Trace: design.sv:81045:3
	wire ram_0_retentive_wd;
	// Trace: design.sv:81046:3
	wire ram_0_retentive_we;
	// Trace: design.sv:81047:3
	wire ram_1_clk_gate_qs;
	// Trace: design.sv:81048:3
	wire ram_1_clk_gate_wd;
	// Trace: design.sv:81049:3
	wire ram_1_clk_gate_we;
	// Trace: design.sv:81050:3
	wire power_gate_ram_block_1_ack_qs;
	// Trace: design.sv:81051:3
	wire ram_1_switch_qs;
	// Trace: design.sv:81052:3
	wire ram_1_switch_wd;
	// Trace: design.sv:81053:3
	wire ram_1_switch_we;
	// Trace: design.sv:81054:3
	wire ram_1_wait_ack_switch_on_qs;
	// Trace: design.sv:81055:3
	wire ram_1_wait_ack_switch_on_wd;
	// Trace: design.sv:81056:3
	wire ram_1_wait_ack_switch_on_we;
	// Trace: design.sv:81057:3
	wire ram_1_iso_qs;
	// Trace: design.sv:81058:3
	wire ram_1_iso_wd;
	// Trace: design.sv:81059:3
	wire ram_1_iso_we;
	// Trace: design.sv:81060:3
	wire ram_1_retentive_qs;
	// Trace: design.sv:81061:3
	wire ram_1_retentive_wd;
	// Trace: design.sv:81062:3
	wire ram_1_retentive_we;
	// Trace: design.sv:81063:3
	wire [2:0] monitor_power_gate_core_qs;
	// Trace: design.sv:81064:3
	wire [2:0] monitor_power_gate_periph_qs;
	// Trace: design.sv:81065:3
	wire [1:0] monitor_power_gate_ram_block_0_qs;
	// Trace: design.sv:81066:3
	wire [1:0] monitor_power_gate_ram_block_1_qs;
	// Trace: design.sv:81067:3
	wire master_cpu_force_switch_off_qs;
	// Trace: design.sv:81068:3
	wire master_cpu_force_switch_off_wd;
	// Trace: design.sv:81069:3
	wire master_cpu_force_switch_off_we;
	// Trace: design.sv:81070:3
	wire master_cpu_force_switch_on_qs;
	// Trace: design.sv:81071:3
	wire master_cpu_force_switch_on_wd;
	// Trace: design.sv:81072:3
	wire master_cpu_force_switch_on_we;
	// Trace: design.sv:81073:3
	wire master_cpu_force_reset_assert_qs;
	// Trace: design.sv:81074:3
	wire master_cpu_force_reset_assert_wd;
	// Trace: design.sv:81075:3
	wire master_cpu_force_reset_assert_we;
	// Trace: design.sv:81076:3
	wire master_cpu_force_reset_deassert_qs;
	// Trace: design.sv:81077:3
	wire master_cpu_force_reset_deassert_wd;
	// Trace: design.sv:81078:3
	wire master_cpu_force_reset_deassert_we;
	// Trace: design.sv:81079:3
	wire master_cpu_force_iso_off_qs;
	// Trace: design.sv:81080:3
	wire master_cpu_force_iso_off_wd;
	// Trace: design.sv:81081:3
	wire master_cpu_force_iso_off_we;
	// Trace: design.sv:81082:3
	wire master_cpu_force_iso_on_qs;
	// Trace: design.sv:81083:3
	wire master_cpu_force_iso_on_wd;
	// Trace: design.sv:81084:3
	wire master_cpu_force_iso_on_we;
	// Trace: design.sv:81089:3
	localparam signed [31:0] sv2v_uu_u_wakeup_state_DW = 1;
	// removed localparam type sv2v_uu_u_wakeup_state_d
	localparam [0:0] sv2v_uu_u_wakeup_state_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_wakeup_state(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wakeup_state_we),
		.wd(wakeup_state_wd),
		.de(1'b0),
		.d(sv2v_uu_u_wakeup_state_ext_d_0),
		.qe(),
		.q(reg2hw[321]),
		.qs(wakeup_state_qs)
	);
	// Trace: design.sv:81116:3
	localparam signed [31:0] sv2v_uu_u_restore_address_DW = 32;
	// removed localparam type sv2v_uu_u_restore_address_d
	localparam [31:0] sv2v_uu_u_restore_address_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_restore_address(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(restore_address_we),
		.wd(restore_address_wd),
		.de(1'b0),
		.d(sv2v_uu_u_restore_address_ext_d_0),
		.qe(),
		.q(reg2hw[320-:32]),
		.qs(restore_address_qs)
	);
	// Trace: design.sv:81143:3
	localparam signed [31:0] sv2v_uu_u_en_wait_for_intr_DW = 32;
	// removed localparam type sv2v_uu_u_en_wait_for_intr_d
	localparam [31:0] sv2v_uu_u_en_wait_for_intr_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_en_wait_for_intr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(en_wait_for_intr_we),
		.wd(en_wait_for_intr_wd),
		.de(1'b0),
		.d(sv2v_uu_u_en_wait_for_intr_ext_d_0),
		.qe(),
		.q(reg2hw[288-:32]),
		.qs(en_wait_for_intr_qs)
	);
	// Trace: design.sv:81170:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_intr_state(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_we),
		.wd(intr_state_wd),
		.de(hw2reg[220]),
		.d(hw2reg[252-:32]),
		.qe(),
		.q(reg2hw[256-:32]),
		.qs(intr_state_qs)
	);
	// Trace: design.sv:81197:3
	localparam signed [31:0] sv2v_uu_u_power_gate_core_DW = 1;
	// removed localparam type sv2v_uu_u_power_gate_core_d
	localparam [0:0] sv2v_uu_u_power_gate_core_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_power_gate_core(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(power_gate_core_we),
		.wd(power_gate_core_wd),
		.de(1'b0),
		.d(sv2v_uu_u_power_gate_core_ext_d_0),
		.qe(),
		.q(reg2hw[224]),
		.qs(power_gate_core_qs)
	);
	// Trace: design.sv:81224:3
	localparam signed [31:0] sv2v_uu_u_power_gate_core_ack_DW = 1;
	// removed localparam type sv2v_uu_u_power_gate_core_ack_wd
	localparam [0:0] sv2v_uu_u_power_gate_core_ack_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_power_gate_core_ack(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_power_gate_core_ack_ext_wd_0),
		.de(hw2reg[218]),
		.d(hw2reg[219]),
		.qe(),
		.q(reg2hw[223]),
		.qs(power_gate_core_ack_qs)
	);
	// Trace: design.sv:81250:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_cpu_reset_assert_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_reset_assert_counter_we),
		.wd(cpu_reset_assert_counter_wd),
		.de(hw2reg[185]),
		.d(hw2reg[217-:32]),
		.qe(),
		.q(reg2hw[222-:32]),
		.qs(cpu_reset_assert_counter_qs)
	);
	// Trace: design.sv:81277:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_cpu_reset_deassert_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_reset_deassert_counter_we),
		.wd(cpu_reset_deassert_counter_wd),
		.de(hw2reg[152]),
		.d(hw2reg[184-:32]),
		.qe(),
		.q(reg2hw[190-:32]),
		.qs(cpu_reset_deassert_counter_qs)
	);
	// Trace: design.sv:81304:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_cpu_switch_off_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_switch_off_counter_we),
		.wd(cpu_switch_off_counter_wd),
		.de(hw2reg[119]),
		.d(hw2reg[151-:32]),
		.qe(),
		.q(reg2hw[158-:32]),
		.qs(cpu_switch_off_counter_qs)
	);
	// Trace: design.sv:81331:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_cpu_switch_on_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_switch_on_counter_we),
		.wd(cpu_switch_on_counter_wd),
		.de(hw2reg[86]),
		.d(hw2reg[118-:32]),
		.qe(),
		.q(reg2hw[126-:32]),
		.qs(cpu_switch_on_counter_qs)
	);
	// Trace: design.sv:81358:3
	localparam signed [31:0] sv2v_uu_u_cpu_wait_ack_switch_on_counter_DW = 1;
	// removed localparam type sv2v_uu_u_cpu_wait_ack_switch_on_counter_d
	localparam [0:0] sv2v_uu_u_cpu_wait_ack_switch_on_counter_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cpu_wait_ack_switch_on_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_wait_ack_switch_on_counter_we),
		.wd(cpu_wait_ack_switch_on_counter_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cpu_wait_ack_switch_on_counter_ext_d_0),
		.qe(),
		.q(reg2hw[94]),
		.qs(cpu_wait_ack_switch_on_counter_qs)
	);
	// Trace: design.sv:81385:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_cpu_iso_off_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_iso_off_counter_we),
		.wd(cpu_iso_off_counter_wd),
		.de(hw2reg[53]),
		.d(hw2reg[85-:32]),
		.qe(),
		.q(reg2hw[93-:32]),
		.qs(cpu_iso_off_counter_qs)
	);
	// Trace: design.sv:81412:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_cpu_iso_on_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_iso_on_counter_we),
		.wd(cpu_iso_on_counter_wd),
		.de(hw2reg[20]),
		.d(hw2reg[52-:32]),
		.qe(),
		.q(reg2hw[61-:32]),
		.qs(cpu_iso_on_counter_qs)
	);
	// Trace: design.sv:81440:3
	localparam signed [31:0] sv2v_uu_u_cpu_counters_stop_cpu_reset_assert_stop_bit_counter_DW = 1;
	// removed localparam type sv2v_uu_u_cpu_counters_stop_cpu_reset_assert_stop_bit_counter_d
	localparam [0:0] sv2v_uu_u_cpu_counters_stop_cpu_reset_assert_stop_bit_counter_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cpu_counters_stop_cpu_reset_assert_stop_bit_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_counters_stop_cpu_reset_assert_stop_bit_counter_we),
		.wd(cpu_counters_stop_cpu_reset_assert_stop_bit_counter_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cpu_counters_stop_cpu_reset_assert_stop_bit_counter_ext_d_0),
		.qe(),
		.q(reg2hw[29]),
		.qs(cpu_counters_stop_cpu_reset_assert_stop_bit_counter_qs)
	);
	// Trace: design.sv:81466:3
	localparam signed [31:0] sv2v_uu_u_cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_DW = 1;
	// removed localparam type sv2v_uu_u_cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_d
	localparam [0:0] sv2v_uu_u_cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cpu_counters_stop_cpu_reset_deassert_stop_bit_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_we),
		.wd(cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_ext_d_0),
		.qe(),
		.q(reg2hw[28]),
		.qs(cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_qs)
	);
	// Trace: design.sv:81492:3
	localparam signed [31:0] sv2v_uu_u_cpu_counters_stop_cpu_switch_off_stop_bit_counter_DW = 1;
	// removed localparam type sv2v_uu_u_cpu_counters_stop_cpu_switch_off_stop_bit_counter_d
	localparam [0:0] sv2v_uu_u_cpu_counters_stop_cpu_switch_off_stop_bit_counter_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cpu_counters_stop_cpu_switch_off_stop_bit_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_counters_stop_cpu_switch_off_stop_bit_counter_we),
		.wd(cpu_counters_stop_cpu_switch_off_stop_bit_counter_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cpu_counters_stop_cpu_switch_off_stop_bit_counter_ext_d_0),
		.qe(),
		.q(reg2hw[27]),
		.qs(cpu_counters_stop_cpu_switch_off_stop_bit_counter_qs)
	);
	// Trace: design.sv:81518:3
	localparam signed [31:0] sv2v_uu_u_cpu_counters_stop_cpu_switch_on_stop_bit_counter_DW = 1;
	// removed localparam type sv2v_uu_u_cpu_counters_stop_cpu_switch_on_stop_bit_counter_d
	localparam [0:0] sv2v_uu_u_cpu_counters_stop_cpu_switch_on_stop_bit_counter_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cpu_counters_stop_cpu_switch_on_stop_bit_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_counters_stop_cpu_switch_on_stop_bit_counter_we),
		.wd(cpu_counters_stop_cpu_switch_on_stop_bit_counter_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cpu_counters_stop_cpu_switch_on_stop_bit_counter_ext_d_0),
		.qe(),
		.q(reg2hw[26]),
		.qs(cpu_counters_stop_cpu_switch_on_stop_bit_counter_qs)
	);
	// Trace: design.sv:81544:3
	localparam signed [31:0] sv2v_uu_u_cpu_counters_stop_cpu_iso_off_stop_bit_counter_DW = 1;
	// removed localparam type sv2v_uu_u_cpu_counters_stop_cpu_iso_off_stop_bit_counter_d
	localparam [0:0] sv2v_uu_u_cpu_counters_stop_cpu_iso_off_stop_bit_counter_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cpu_counters_stop_cpu_iso_off_stop_bit_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_counters_stop_cpu_iso_off_stop_bit_counter_we),
		.wd(cpu_counters_stop_cpu_iso_off_stop_bit_counter_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cpu_counters_stop_cpu_iso_off_stop_bit_counter_ext_d_0),
		.qe(),
		.q(reg2hw[25]),
		.qs(cpu_counters_stop_cpu_iso_off_stop_bit_counter_qs)
	);
	// Trace: design.sv:81570:3
	localparam signed [31:0] sv2v_uu_u_cpu_counters_stop_cpu_iso_on_stop_bit_counter_DW = 1;
	// removed localparam type sv2v_uu_u_cpu_counters_stop_cpu_iso_on_stop_bit_counter_d
	localparam [0:0] sv2v_uu_u_cpu_counters_stop_cpu_iso_on_stop_bit_counter_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_cpu_counters_stop_cpu_iso_on_stop_bit_counter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cpu_counters_stop_cpu_iso_on_stop_bit_counter_we),
		.wd(cpu_counters_stop_cpu_iso_on_stop_bit_counter_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cpu_counters_stop_cpu_iso_on_stop_bit_counter_ext_d_0),
		.qe(),
		.q(reg2hw[24]),
		.qs(cpu_counters_stop_cpu_iso_on_stop_bit_counter_qs)
	);
	// Trace: design.sv:81597:3
	localparam signed [31:0] sv2v_uu_u_power_gate_periph_ack_DW = 1;
	// removed localparam type sv2v_uu_u_power_gate_periph_ack_wd
	localparam [0:0] sv2v_uu_u_power_gate_periph_ack_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_power_gate_periph_ack(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_power_gate_periph_ack_ext_wd_0),
		.de(hw2reg[18]),
		.d(hw2reg[19]),
		.qe(),
		.q(reg2hw[23]),
		.qs(power_gate_periph_ack_qs)
	);
	// Trace: design.sv:81623:3
	localparam signed [31:0] sv2v_uu_u_periph_reset_DW = 1;
	// removed localparam type sv2v_uu_u_periph_reset_d
	localparam [0:0] sv2v_uu_u_periph_reset_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_periph_reset(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(periph_reset_we),
		.wd(periph_reset_wd),
		.de(1'b0),
		.d(sv2v_uu_u_periph_reset_ext_d_0),
		.qe(),
		.q(reg2hw[22]),
		.qs(periph_reset_qs)
	);
	// Trace: design.sv:81650:3
	localparam signed [31:0] sv2v_uu_u_periph_switch_DW = 1;
	// removed localparam type sv2v_uu_u_periph_switch_d
	localparam [0:0] sv2v_uu_u_periph_switch_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_periph_switch(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(periph_switch_we),
		.wd(periph_switch_wd),
		.de(1'b0),
		.d(sv2v_uu_u_periph_switch_ext_d_0),
		.qe(),
		.q(reg2hw[21]),
		.qs(periph_switch_qs)
	);
	// Trace: design.sv:81677:3
	localparam signed [31:0] sv2v_uu_u_periph_wait_ack_switch_on_DW = 1;
	// removed localparam type sv2v_uu_u_periph_wait_ack_switch_on_d
	localparam [0:0] sv2v_uu_u_periph_wait_ack_switch_on_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_periph_wait_ack_switch_on(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(periph_wait_ack_switch_on_we),
		.wd(periph_wait_ack_switch_on_wd),
		.de(1'b0),
		.d(sv2v_uu_u_periph_wait_ack_switch_on_ext_d_0),
		.qe(),
		.q(reg2hw[20]),
		.qs(periph_wait_ack_switch_on_qs)
	);
	// Trace: design.sv:81704:3
	localparam signed [31:0] sv2v_uu_u_periph_iso_DW = 1;
	// removed localparam type sv2v_uu_u_periph_iso_d
	localparam [0:0] sv2v_uu_u_periph_iso_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_periph_iso(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(periph_iso_we),
		.wd(periph_iso_wd),
		.de(1'b0),
		.d(sv2v_uu_u_periph_iso_ext_d_0),
		.qe(),
		.q(reg2hw[19]),
		.qs(periph_iso_qs)
	);
	// Trace: design.sv:81731:3
	localparam signed [31:0] sv2v_uu_u_periph_clk_gate_DW = 1;
	// removed localparam type sv2v_uu_u_periph_clk_gate_d
	localparam [0:0] sv2v_uu_u_periph_clk_gate_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_periph_clk_gate(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(periph_clk_gate_we),
		.wd(periph_clk_gate_wd),
		.de(1'b0),
		.d(sv2v_uu_u_periph_clk_gate_ext_d_0),
		.qe(),
		.q(reg2hw[18]),
		.qs(periph_clk_gate_qs)
	);
	// Trace: design.sv:81758:3
	localparam signed [31:0] sv2v_uu_u_ram_0_clk_gate_DW = 1;
	// removed localparam type sv2v_uu_u_ram_0_clk_gate_d
	localparam [0:0] sv2v_uu_u_ram_0_clk_gate_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_0_clk_gate(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_0_clk_gate_we),
		.wd(ram_0_clk_gate_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_0_clk_gate_ext_d_0),
		.qe(),
		.q(reg2hw[17]),
		.qs(ram_0_clk_gate_qs)
	);
	// Trace: design.sv:81785:3
	localparam signed [31:0] sv2v_uu_u_power_gate_ram_block_0_ack_DW = 1;
	// removed localparam type sv2v_uu_u_power_gate_ram_block_0_ack_wd
	localparam [0:0] sv2v_uu_u_power_gate_ram_block_0_ack_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_power_gate_ram_block_0_ack(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_power_gate_ram_block_0_ack_ext_wd_0),
		.de(hw2reg[16]),
		.d(hw2reg[17]),
		.qe(),
		.q(reg2hw[16]),
		.qs(power_gate_ram_block_0_ack_qs)
	);
	// Trace: design.sv:81811:3
	localparam signed [31:0] sv2v_uu_u_ram_0_switch_DW = 1;
	// removed localparam type sv2v_uu_u_ram_0_switch_d
	localparam [0:0] sv2v_uu_u_ram_0_switch_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_0_switch(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_0_switch_we),
		.wd(ram_0_switch_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_0_switch_ext_d_0),
		.qe(),
		.q(reg2hw[15]),
		.qs(ram_0_switch_qs)
	);
	// Trace: design.sv:81838:3
	localparam signed [31:0] sv2v_uu_u_ram_0_wait_ack_switch_on_DW = 1;
	// removed localparam type sv2v_uu_u_ram_0_wait_ack_switch_on_d
	localparam [0:0] sv2v_uu_u_ram_0_wait_ack_switch_on_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_0_wait_ack_switch_on(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_0_wait_ack_switch_on_we),
		.wd(ram_0_wait_ack_switch_on_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_0_wait_ack_switch_on_ext_d_0),
		.qe(),
		.q(reg2hw[14]),
		.qs(ram_0_wait_ack_switch_on_qs)
	);
	// Trace: design.sv:81865:3
	localparam signed [31:0] sv2v_uu_u_ram_0_iso_DW = 1;
	// removed localparam type sv2v_uu_u_ram_0_iso_d
	localparam [0:0] sv2v_uu_u_ram_0_iso_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_0_iso(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_0_iso_we),
		.wd(ram_0_iso_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_0_iso_ext_d_0),
		.qe(),
		.q(reg2hw[13]),
		.qs(ram_0_iso_qs)
	);
	// Trace: design.sv:81892:3
	localparam signed [31:0] sv2v_uu_u_ram_0_retentive_DW = 1;
	// removed localparam type sv2v_uu_u_ram_0_retentive_d
	localparam [0:0] sv2v_uu_u_ram_0_retentive_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_0_retentive(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_0_retentive_we),
		.wd(ram_0_retentive_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_0_retentive_ext_d_0),
		.qe(),
		.q(reg2hw[12]),
		.qs(ram_0_retentive_qs)
	);
	// Trace: design.sv:81919:3
	localparam signed [31:0] sv2v_uu_u_ram_1_clk_gate_DW = 1;
	// removed localparam type sv2v_uu_u_ram_1_clk_gate_d
	localparam [0:0] sv2v_uu_u_ram_1_clk_gate_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_1_clk_gate(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_1_clk_gate_we),
		.wd(ram_1_clk_gate_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_1_clk_gate_ext_d_0),
		.qe(),
		.q(reg2hw[11]),
		.qs(ram_1_clk_gate_qs)
	);
	// Trace: design.sv:81946:3
	localparam signed [31:0] sv2v_uu_u_power_gate_ram_block_1_ack_DW = 1;
	// removed localparam type sv2v_uu_u_power_gate_ram_block_1_ack_wd
	localparam [0:0] sv2v_uu_u_power_gate_ram_block_1_ack_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_power_gate_ram_block_1_ack(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_power_gate_ram_block_1_ack_ext_wd_0),
		.de(hw2reg[14]),
		.d(hw2reg[15]),
		.qe(),
		.q(reg2hw[10]),
		.qs(power_gate_ram_block_1_ack_qs)
	);
	// Trace: design.sv:81972:3
	localparam signed [31:0] sv2v_uu_u_ram_1_switch_DW = 1;
	// removed localparam type sv2v_uu_u_ram_1_switch_d
	localparam [0:0] sv2v_uu_u_ram_1_switch_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_1_switch(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_1_switch_we),
		.wd(ram_1_switch_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_1_switch_ext_d_0),
		.qe(),
		.q(reg2hw[9]),
		.qs(ram_1_switch_qs)
	);
	// Trace: design.sv:81999:3
	localparam signed [31:0] sv2v_uu_u_ram_1_wait_ack_switch_on_DW = 1;
	// removed localparam type sv2v_uu_u_ram_1_wait_ack_switch_on_d
	localparam [0:0] sv2v_uu_u_ram_1_wait_ack_switch_on_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_1_wait_ack_switch_on(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_1_wait_ack_switch_on_we),
		.wd(ram_1_wait_ack_switch_on_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_1_wait_ack_switch_on_ext_d_0),
		.qe(),
		.q(reg2hw[8]),
		.qs(ram_1_wait_ack_switch_on_qs)
	);
	// Trace: design.sv:82026:3
	localparam signed [31:0] sv2v_uu_u_ram_1_iso_DW = 1;
	// removed localparam type sv2v_uu_u_ram_1_iso_d
	localparam [0:0] sv2v_uu_u_ram_1_iso_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_1_iso(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_1_iso_we),
		.wd(ram_1_iso_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_1_iso_ext_d_0),
		.qe(),
		.q(reg2hw[7]),
		.qs(ram_1_iso_qs)
	);
	// Trace: design.sv:82053:3
	localparam signed [31:0] sv2v_uu_u_ram_1_retentive_DW = 1;
	// removed localparam type sv2v_uu_u_ram_1_retentive_d
	localparam [0:0] sv2v_uu_u_ram_1_retentive_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ram_1_retentive(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ram_1_retentive_we),
		.wd(ram_1_retentive_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ram_1_retentive_ext_d_0),
		.qe(),
		.q(reg2hw[6]),
		.qs(ram_1_retentive_qs)
	);
	// Trace: design.sv:82080:3
	localparam signed [31:0] sv2v_uu_u_monitor_power_gate_core_DW = 3;
	// removed localparam type sv2v_uu_u_monitor_power_gate_core_wd
	localparam [2:0] sv2v_uu_u_monitor_power_gate_core_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RO"),
		.RESVAL(3'h0)
	) u_monitor_power_gate_core(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_monitor_power_gate_core_ext_wd_0),
		.de(hw2reg[10]),
		.d(hw2reg[13-:3]),
		.qe(),
		.q(),
		.qs(monitor_power_gate_core_qs)
	);
	// Trace: design.sv:82106:3
	localparam signed [31:0] sv2v_uu_u_monitor_power_gate_periph_DW = 3;
	// removed localparam type sv2v_uu_u_monitor_power_gate_periph_wd
	localparam [2:0] sv2v_uu_u_monitor_power_gate_periph_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RO"),
		.RESVAL(3'h0)
	) u_monitor_power_gate_periph(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_monitor_power_gate_periph_ext_wd_0),
		.de(hw2reg[6]),
		.d(hw2reg[9-:3]),
		.qe(),
		.q(),
		.qs(monitor_power_gate_periph_qs)
	);
	// Trace: design.sv:82132:3
	localparam signed [31:0] sv2v_uu_u_monitor_power_gate_ram_block_0_DW = 2;
	// removed localparam type sv2v_uu_u_monitor_power_gate_ram_block_0_wd
	localparam [1:0] sv2v_uu_u_monitor_power_gate_ram_block_0_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RO"),
		.RESVAL(2'h0)
	) u_monitor_power_gate_ram_block_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_monitor_power_gate_ram_block_0_ext_wd_0),
		.de(hw2reg[3]),
		.d(hw2reg[5-:2]),
		.qe(),
		.q(),
		.qs(monitor_power_gate_ram_block_0_qs)
	);
	// Trace: design.sv:82158:3
	localparam signed [31:0] sv2v_uu_u_monitor_power_gate_ram_block_1_DW = 2;
	// removed localparam type sv2v_uu_u_monitor_power_gate_ram_block_1_wd
	localparam [1:0] sv2v_uu_u_monitor_power_gate_ram_block_1_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RO"),
		.RESVAL(2'h0)
	) u_monitor_power_gate_ram_block_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_monitor_power_gate_ram_block_1_ext_wd_0),
		.de(hw2reg[0]),
		.d(hw2reg[2-:2]),
		.qe(),
		.q(),
		.qs(monitor_power_gate_ram_block_1_qs)
	);
	// Trace: design.sv:82184:3
	localparam signed [31:0] sv2v_uu_u_master_cpu_force_switch_off_DW = 1;
	// removed localparam type sv2v_uu_u_master_cpu_force_switch_off_d
	localparam [0:0] sv2v_uu_u_master_cpu_force_switch_off_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_master_cpu_force_switch_off(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(master_cpu_force_switch_off_we),
		.wd(master_cpu_force_switch_off_wd),
		.de(1'b0),
		.d(sv2v_uu_u_master_cpu_force_switch_off_ext_d_0),
		.qe(),
		.q(reg2hw[5]),
		.qs(master_cpu_force_switch_off_qs)
	);
	// Trace: design.sv:82211:3
	localparam signed [31:0] sv2v_uu_u_master_cpu_force_switch_on_DW = 1;
	// removed localparam type sv2v_uu_u_master_cpu_force_switch_on_d
	localparam [0:0] sv2v_uu_u_master_cpu_force_switch_on_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_master_cpu_force_switch_on(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(master_cpu_force_switch_on_we),
		.wd(master_cpu_force_switch_on_wd),
		.de(1'b0),
		.d(sv2v_uu_u_master_cpu_force_switch_on_ext_d_0),
		.qe(),
		.q(reg2hw[4]),
		.qs(master_cpu_force_switch_on_qs)
	);
	// Trace: design.sv:82238:3
	localparam signed [31:0] sv2v_uu_u_master_cpu_force_reset_assert_DW = 1;
	// removed localparam type sv2v_uu_u_master_cpu_force_reset_assert_d
	localparam [0:0] sv2v_uu_u_master_cpu_force_reset_assert_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_master_cpu_force_reset_assert(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(master_cpu_force_reset_assert_we),
		.wd(master_cpu_force_reset_assert_wd),
		.de(1'b0),
		.d(sv2v_uu_u_master_cpu_force_reset_assert_ext_d_0),
		.qe(),
		.q(reg2hw[3]),
		.qs(master_cpu_force_reset_assert_qs)
	);
	// Trace: design.sv:82265:3
	localparam signed [31:0] sv2v_uu_u_master_cpu_force_reset_deassert_DW = 1;
	// removed localparam type sv2v_uu_u_master_cpu_force_reset_deassert_d
	localparam [0:0] sv2v_uu_u_master_cpu_force_reset_deassert_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_master_cpu_force_reset_deassert(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(master_cpu_force_reset_deassert_we),
		.wd(master_cpu_force_reset_deassert_wd),
		.de(1'b0),
		.d(sv2v_uu_u_master_cpu_force_reset_deassert_ext_d_0),
		.qe(),
		.q(reg2hw[2]),
		.qs(master_cpu_force_reset_deassert_qs)
	);
	// Trace: design.sv:82292:3
	localparam signed [31:0] sv2v_uu_u_master_cpu_force_iso_off_DW = 1;
	// removed localparam type sv2v_uu_u_master_cpu_force_iso_off_d
	localparam [0:0] sv2v_uu_u_master_cpu_force_iso_off_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_master_cpu_force_iso_off(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(master_cpu_force_iso_off_we),
		.wd(master_cpu_force_iso_off_wd),
		.de(1'b0),
		.d(sv2v_uu_u_master_cpu_force_iso_off_ext_d_0),
		.qe(),
		.q(reg2hw[1]),
		.qs(master_cpu_force_iso_off_qs)
	);
	// Trace: design.sv:82319:3
	localparam signed [31:0] sv2v_uu_u_master_cpu_force_iso_on_DW = 1;
	// removed localparam type sv2v_uu_u_master_cpu_force_iso_on_d
	localparam [0:0] sv2v_uu_u_master_cpu_force_iso_on_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_master_cpu_force_iso_on(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(master_cpu_force_iso_on_we),
		.wd(master_cpu_force_iso_on_wd),
		.de(1'b0),
		.d(sv2v_uu_u_master_cpu_force_iso_on_ext_d_0),
		.qe(),
		.q(reg2hw[-0]),
		.qs(master_cpu_force_iso_on_qs)
	);
	// Trace: design.sv:82346:3
	reg [41:0] addr_hit;
	// Trace: design.sv:82347:3
	localparam signed [31:0] power_manager_reg_pkg_BlockAw = 8;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_CPU_COUNTERS_STOP_OFFSET = 8'h34;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_CPU_ISO_OFF_COUNTER_OFFSET = 8'h2c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_CPU_ISO_ON_COUNTER_OFFSET = 8'h30;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_CPU_RESET_ASSERT_COUNTER_OFFSET = 8'h18;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_CPU_RESET_DEASSERT_COUNTER_OFFSET = 8'h1c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_CPU_SWITCH_OFF_COUNTER_OFFSET = 8'h20;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_CPU_SWITCH_ON_COUNTER_OFFSET = 8'h24;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_CPU_WAIT_ACK_SWITCH_ON_COUNTER_OFFSET = 8'h28;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_EN_WAIT_FOR_INTR_OFFSET = 8'h08;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_INTR_STATE_OFFSET = 8'h0c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_ISO_OFF_OFFSET = 8'ha0;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_ISO_ON_OFFSET = 8'ha4;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_RESET_ASSERT_OFFSET = 8'h98;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_RESET_DEASSERT_OFFSET = 8'h9c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_SWITCH_OFF_OFFSET = 8'h90;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_SWITCH_ON_OFFSET = 8'h94;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MONITOR_POWER_GATE_CORE_OFFSET = 8'h80;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MONITOR_POWER_GATE_PERIPH_OFFSET = 8'h84;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MONITOR_POWER_GATE_RAM_BLOCK_0_OFFSET = 8'h88;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_MONITOR_POWER_GATE_RAM_BLOCK_1_OFFSET = 8'h8c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_PERIPH_CLK_GATE_OFFSET = 8'h4c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_PERIPH_ISO_OFFSET = 8'h48;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_PERIPH_RESET_OFFSET = 8'h3c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_PERIPH_SWITCH_OFFSET = 8'h40;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_PERIPH_WAIT_ACK_SWITCH_ON_OFFSET = 8'h44;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_CORE_ACK_OFFSET = 8'h14;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_CORE_OFFSET = 8'h10;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_PERIPH_ACK_OFFSET = 8'h38;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_RAM_BLOCK_0_ACK_OFFSET = 8'h54;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_RAM_BLOCK_1_ACK_OFFSET = 8'h6c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_0_CLK_GATE_OFFSET = 8'h50;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_0_ISO_OFFSET = 8'h60;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_0_RETENTIVE_OFFSET = 8'h64;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_0_SWITCH_OFFSET = 8'h58;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_0_WAIT_ACK_SWITCH_ON_OFFSET = 8'h5c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_1_CLK_GATE_OFFSET = 8'h68;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_1_ISO_OFFSET = 8'h78;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_1_RETENTIVE_OFFSET = 8'h7c;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_1_SWITCH_OFFSET = 8'h70;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RAM_1_WAIT_ACK_SWITCH_ON_OFFSET = 8'h74;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_RESTORE_ADDRESS_OFFSET = 8'h04;
	localparam [7:0] power_manager_reg_pkg_POWER_MANAGER_WAKEUP_STATE_OFFSET = 8'h00;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:82348:5
		addr_hit = 1'sb0;
		// Trace: design.sv:82349:5
		addr_hit[0] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_WAKEUP_STATE_OFFSET;
		// Trace: design.sv:82350:5
		addr_hit[1] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RESTORE_ADDRESS_OFFSET;
		// Trace: design.sv:82351:5
		addr_hit[2] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_EN_WAIT_FOR_INTR_OFFSET;
		// Trace: design.sv:82352:5
		addr_hit[3] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_INTR_STATE_OFFSET;
		// Trace: design.sv:82353:5
		addr_hit[4] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_CORE_OFFSET;
		// Trace: design.sv:82354:5
		addr_hit[5] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_CORE_ACK_OFFSET;
		// Trace: design.sv:82355:5
		addr_hit[6] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_CPU_RESET_ASSERT_COUNTER_OFFSET;
		// Trace: design.sv:82356:5
		addr_hit[7] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_CPU_RESET_DEASSERT_COUNTER_OFFSET;
		// Trace: design.sv:82357:5
		addr_hit[8] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_CPU_SWITCH_OFF_COUNTER_OFFSET;
		// Trace: design.sv:82358:5
		addr_hit[9] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_CPU_SWITCH_ON_COUNTER_OFFSET;
		// Trace: design.sv:82359:5
		addr_hit[10] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_CPU_WAIT_ACK_SWITCH_ON_COUNTER_OFFSET;
		// Trace: design.sv:82360:5
		addr_hit[11] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_CPU_ISO_OFF_COUNTER_OFFSET;
		// Trace: design.sv:82361:5
		addr_hit[12] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_CPU_ISO_ON_COUNTER_OFFSET;
		// Trace: design.sv:82362:5
		addr_hit[13] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_CPU_COUNTERS_STOP_OFFSET;
		// Trace: design.sv:82363:5
		addr_hit[14] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_PERIPH_ACK_OFFSET;
		// Trace: design.sv:82364:5
		addr_hit[15] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_PERIPH_RESET_OFFSET;
		// Trace: design.sv:82365:5
		addr_hit[16] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_PERIPH_SWITCH_OFFSET;
		// Trace: design.sv:82366:5
		addr_hit[17] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_PERIPH_WAIT_ACK_SWITCH_ON_OFFSET;
		// Trace: design.sv:82367:5
		addr_hit[18] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_PERIPH_ISO_OFFSET;
		// Trace: design.sv:82368:5
		addr_hit[19] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_PERIPH_CLK_GATE_OFFSET;
		// Trace: design.sv:82369:5
		addr_hit[20] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_0_CLK_GATE_OFFSET;
		// Trace: design.sv:82370:5
		addr_hit[21] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_RAM_BLOCK_0_ACK_OFFSET;
		// Trace: design.sv:82371:5
		addr_hit[22] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_0_SWITCH_OFFSET;
		// Trace: design.sv:82372:5
		addr_hit[23] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_0_WAIT_ACK_SWITCH_ON_OFFSET;
		// Trace: design.sv:82373:5
		addr_hit[24] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_0_ISO_OFFSET;
		// Trace: design.sv:82374:5
		addr_hit[25] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_0_RETENTIVE_OFFSET;
		// Trace: design.sv:82375:5
		addr_hit[26] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_1_CLK_GATE_OFFSET;
		// Trace: design.sv:82376:5
		addr_hit[27] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_POWER_GATE_RAM_BLOCK_1_ACK_OFFSET;
		// Trace: design.sv:82377:5
		addr_hit[28] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_1_SWITCH_OFFSET;
		// Trace: design.sv:82378:5
		addr_hit[29] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_1_WAIT_ACK_SWITCH_ON_OFFSET;
		// Trace: design.sv:82379:5
		addr_hit[30] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_1_ISO_OFFSET;
		// Trace: design.sv:82380:5
		addr_hit[31] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_RAM_1_RETENTIVE_OFFSET;
		// Trace: design.sv:82381:5
		addr_hit[32] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MONITOR_POWER_GATE_CORE_OFFSET;
		// Trace: design.sv:82382:5
		addr_hit[33] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MONITOR_POWER_GATE_PERIPH_OFFSET;
		// Trace: design.sv:82383:5
		addr_hit[34] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MONITOR_POWER_GATE_RAM_BLOCK_0_OFFSET;
		// Trace: design.sv:82384:5
		addr_hit[35] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MONITOR_POWER_GATE_RAM_BLOCK_1_OFFSET;
		// Trace: design.sv:82385:5
		addr_hit[36] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_SWITCH_OFF_OFFSET;
		// Trace: design.sv:82386:5
		addr_hit[37] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_SWITCH_ON_OFFSET;
		// Trace: design.sv:82387:5
		addr_hit[38] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_RESET_ASSERT_OFFSET;
		// Trace: design.sv:82388:5
		addr_hit[39] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_RESET_DEASSERT_OFFSET;
		// Trace: design.sv:82389:5
		addr_hit[40] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_ISO_OFF_OFFSET;
		// Trace: design.sv:82390:5
		addr_hit[41] = reg_addr == power_manager_reg_pkg_POWER_MANAGER_MASTER_CPU_FORCE_ISO_ON_OFFSET;
	end
	// Trace: design.sv:82393:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:82396:3
	localparam [167:0] power_manager_reg_pkg_POWER_MANAGER_PERMIT = 168'b000111111111111100010001111111111111111100011111111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:82397:5
		wr_err = reg_we & ((((((((((((((((((((((((((((((((((((((((((addr_hit[0] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[164+:4] & ~reg_be)) | (addr_hit[1] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[160+:4] & ~reg_be))) | (addr_hit[2] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[156+:4] & ~reg_be))) | (addr_hit[3] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[152+:4] & ~reg_be))) | (addr_hit[4] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[148+:4] & ~reg_be))) | (addr_hit[5] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[144+:4] & ~reg_be))) | (addr_hit[6] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[140+:4] & ~reg_be))) | (addr_hit[7] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[136+:4] & ~reg_be))) | (addr_hit[8] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[132+:4] & ~reg_be))) | (addr_hit[9] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[128+:4] & ~reg_be))) | (addr_hit[10] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[124+:4] & ~reg_be))) | (addr_hit[11] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[120+:4] & ~reg_be))) | (addr_hit[12] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[116+:4] & ~reg_be))) | (addr_hit[13] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[112+:4] & ~reg_be))) | (addr_hit[14] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[108+:4] & ~reg_be))) | (addr_hit[15] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[104+:4] & ~reg_be))) | (addr_hit[16] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[100+:4] & ~reg_be))) | (addr_hit[17] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[96+:4] & ~reg_be))) | (addr_hit[18] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[92+:4] & ~reg_be))) | (addr_hit[19] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[88+:4] & ~reg_be))) | (addr_hit[20] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[84+:4] & ~reg_be))) | (addr_hit[21] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[80+:4] & ~reg_be))) | (addr_hit[22] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[76+:4] & ~reg_be))) | (addr_hit[23] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[72+:4] & ~reg_be))) | (addr_hit[24] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[68+:4] & ~reg_be))) | (addr_hit[25] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[64+:4] & ~reg_be))) | (addr_hit[26] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[60+:4] & ~reg_be))) | (addr_hit[27] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[56+:4] & ~reg_be))) | (addr_hit[28] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[52+:4] & ~reg_be))) | (addr_hit[29] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[48+:4] & ~reg_be))) | (addr_hit[30] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[44+:4] & ~reg_be))) | (addr_hit[31] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[40+:4] & ~reg_be))) | (addr_hit[32] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[36+:4] & ~reg_be))) | (addr_hit[33] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[32+:4] & ~reg_be))) | (addr_hit[34] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[28+:4] & ~reg_be))) | (addr_hit[35] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[24+:4] & ~reg_be))) | (addr_hit[36] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[20+:4] & ~reg_be))) | (addr_hit[37] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[16+:4] & ~reg_be))) | (addr_hit[38] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[12+:4] & ~reg_be))) | (addr_hit[39] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[8+:4] & ~reg_be))) | (addr_hit[40] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[4+:4] & ~reg_be))) | (addr_hit[41] & |(power_manager_reg_pkg_POWER_MANAGER_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:82442:3
	assign wakeup_state_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:82443:3
	assign wakeup_state_wd = reg_wdata[0];
	// Trace: design.sv:82445:3
	assign restore_address_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:82446:3
	assign restore_address_wd = reg_wdata[31:0];
	// Trace: design.sv:82448:3
	assign en_wait_for_intr_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:82449:3
	assign en_wait_for_intr_wd = reg_wdata[31:0];
	// Trace: design.sv:82451:3
	assign intr_state_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:82452:3
	assign intr_state_wd = reg_wdata[31:0];
	// Trace: design.sv:82454:3
	assign power_gate_core_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:82455:3
	assign power_gate_core_wd = reg_wdata[0];
	// Trace: design.sv:82457:3
	assign cpu_reset_assert_counter_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:82458:3
	assign cpu_reset_assert_counter_wd = reg_wdata[31:0];
	// Trace: design.sv:82460:3
	assign cpu_reset_deassert_counter_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:82461:3
	assign cpu_reset_deassert_counter_wd = reg_wdata[31:0];
	// Trace: design.sv:82463:3
	assign cpu_switch_off_counter_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:82464:3
	assign cpu_switch_off_counter_wd = reg_wdata[31:0];
	// Trace: design.sv:82466:3
	assign cpu_switch_on_counter_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:82467:3
	assign cpu_switch_on_counter_wd = reg_wdata[31:0];
	// Trace: design.sv:82469:3
	assign cpu_wait_ack_switch_on_counter_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:82470:3
	assign cpu_wait_ack_switch_on_counter_wd = reg_wdata[0];
	// Trace: design.sv:82472:3
	assign cpu_iso_off_counter_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:82473:3
	assign cpu_iso_off_counter_wd = reg_wdata[31:0];
	// Trace: design.sv:82475:3
	assign cpu_iso_on_counter_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:82476:3
	assign cpu_iso_on_counter_wd = reg_wdata[31:0];
	// Trace: design.sv:82478:3
	assign cpu_counters_stop_cpu_reset_assert_stop_bit_counter_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:82479:3
	assign cpu_counters_stop_cpu_reset_assert_stop_bit_counter_wd = reg_wdata[0];
	// Trace: design.sv:82481:3
	assign cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:82482:3
	assign cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_wd = reg_wdata[1];
	// Trace: design.sv:82484:3
	assign cpu_counters_stop_cpu_switch_off_stop_bit_counter_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:82485:3
	assign cpu_counters_stop_cpu_switch_off_stop_bit_counter_wd = reg_wdata[2];
	// Trace: design.sv:82487:3
	assign cpu_counters_stop_cpu_switch_on_stop_bit_counter_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:82488:3
	assign cpu_counters_stop_cpu_switch_on_stop_bit_counter_wd = reg_wdata[3];
	// Trace: design.sv:82490:3
	assign cpu_counters_stop_cpu_iso_off_stop_bit_counter_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:82491:3
	assign cpu_counters_stop_cpu_iso_off_stop_bit_counter_wd = reg_wdata[4];
	// Trace: design.sv:82493:3
	assign cpu_counters_stop_cpu_iso_on_stop_bit_counter_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:82494:3
	assign cpu_counters_stop_cpu_iso_on_stop_bit_counter_wd = reg_wdata[5];
	// Trace: design.sv:82496:3
	assign periph_reset_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:82497:3
	assign periph_reset_wd = reg_wdata[0];
	// Trace: design.sv:82499:3
	assign periph_switch_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:82500:3
	assign periph_switch_wd = reg_wdata[0];
	// Trace: design.sv:82502:3
	assign periph_wait_ack_switch_on_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:82503:3
	assign periph_wait_ack_switch_on_wd = reg_wdata[0];
	// Trace: design.sv:82505:3
	assign periph_iso_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:82506:3
	assign periph_iso_wd = reg_wdata[0];
	// Trace: design.sv:82508:3
	assign periph_clk_gate_we = (addr_hit[19] & reg_we) & !reg_error;
	// Trace: design.sv:82509:3
	assign periph_clk_gate_wd = reg_wdata[0];
	// Trace: design.sv:82511:3
	assign ram_0_clk_gate_we = (addr_hit[20] & reg_we) & !reg_error;
	// Trace: design.sv:82512:3
	assign ram_0_clk_gate_wd = reg_wdata[0];
	// Trace: design.sv:82514:3
	assign ram_0_switch_we = (addr_hit[22] & reg_we) & !reg_error;
	// Trace: design.sv:82515:3
	assign ram_0_switch_wd = reg_wdata[0];
	// Trace: design.sv:82517:3
	assign ram_0_wait_ack_switch_on_we = (addr_hit[23] & reg_we) & !reg_error;
	// Trace: design.sv:82518:3
	assign ram_0_wait_ack_switch_on_wd = reg_wdata[0];
	// Trace: design.sv:82520:3
	assign ram_0_iso_we = (addr_hit[24] & reg_we) & !reg_error;
	// Trace: design.sv:82521:3
	assign ram_0_iso_wd = reg_wdata[0];
	// Trace: design.sv:82523:3
	assign ram_0_retentive_we = (addr_hit[25] & reg_we) & !reg_error;
	// Trace: design.sv:82524:3
	assign ram_0_retentive_wd = reg_wdata[0];
	// Trace: design.sv:82526:3
	assign ram_1_clk_gate_we = (addr_hit[26] & reg_we) & !reg_error;
	// Trace: design.sv:82527:3
	assign ram_1_clk_gate_wd = reg_wdata[0];
	// Trace: design.sv:82529:3
	assign ram_1_switch_we = (addr_hit[28] & reg_we) & !reg_error;
	// Trace: design.sv:82530:3
	assign ram_1_switch_wd = reg_wdata[0];
	// Trace: design.sv:82532:3
	assign ram_1_wait_ack_switch_on_we = (addr_hit[29] & reg_we) & !reg_error;
	// Trace: design.sv:82533:3
	assign ram_1_wait_ack_switch_on_wd = reg_wdata[0];
	// Trace: design.sv:82535:3
	assign ram_1_iso_we = (addr_hit[30] & reg_we) & !reg_error;
	// Trace: design.sv:82536:3
	assign ram_1_iso_wd = reg_wdata[0];
	// Trace: design.sv:82538:3
	assign ram_1_retentive_we = (addr_hit[31] & reg_we) & !reg_error;
	// Trace: design.sv:82539:3
	assign ram_1_retentive_wd = reg_wdata[0];
	// Trace: design.sv:82541:3
	assign master_cpu_force_switch_off_we = (addr_hit[36] & reg_we) & !reg_error;
	// Trace: design.sv:82542:3
	assign master_cpu_force_switch_off_wd = reg_wdata[0];
	// Trace: design.sv:82544:3
	assign master_cpu_force_switch_on_we = (addr_hit[37] & reg_we) & !reg_error;
	// Trace: design.sv:82545:3
	assign master_cpu_force_switch_on_wd = reg_wdata[0];
	// Trace: design.sv:82547:3
	assign master_cpu_force_reset_assert_we = (addr_hit[38] & reg_we) & !reg_error;
	// Trace: design.sv:82548:3
	assign master_cpu_force_reset_assert_wd = reg_wdata[0];
	// Trace: design.sv:82550:3
	assign master_cpu_force_reset_deassert_we = (addr_hit[39] & reg_we) & !reg_error;
	// Trace: design.sv:82551:3
	assign master_cpu_force_reset_deassert_wd = reg_wdata[0];
	// Trace: design.sv:82553:3
	assign master_cpu_force_iso_off_we = (addr_hit[40] & reg_we) & !reg_error;
	// Trace: design.sv:82554:3
	assign master_cpu_force_iso_off_wd = reg_wdata[0];
	// Trace: design.sv:82556:3
	assign master_cpu_force_iso_on_we = (addr_hit[41] & reg_we) & !reg_error;
	// Trace: design.sv:82557:3
	assign master_cpu_force_iso_on_wd = reg_wdata[0];
	// Trace: design.sv:82560:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:82561:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:82562:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]:
				// Trace: design.sv:82564:9
				reg_rdata_next[0] = wakeup_state_qs;
			addr_hit[1]:
				// Trace: design.sv:82568:9
				reg_rdata_next[31:0] = restore_address_qs;
			addr_hit[2]:
				// Trace: design.sv:82572:9
				reg_rdata_next[31:0] = en_wait_for_intr_qs;
			addr_hit[3]:
				// Trace: design.sv:82576:9
				reg_rdata_next[31:0] = intr_state_qs;
			addr_hit[4]:
				// Trace: design.sv:82580:9
				reg_rdata_next[0] = power_gate_core_qs;
			addr_hit[5]:
				// Trace: design.sv:82584:9
				reg_rdata_next[0] = power_gate_core_ack_qs;
			addr_hit[6]:
				// Trace: design.sv:82588:9
				reg_rdata_next[31:0] = cpu_reset_assert_counter_qs;
			addr_hit[7]:
				// Trace: design.sv:82592:9
				reg_rdata_next[31:0] = cpu_reset_deassert_counter_qs;
			addr_hit[8]:
				// Trace: design.sv:82596:9
				reg_rdata_next[31:0] = cpu_switch_off_counter_qs;
			addr_hit[9]:
				// Trace: design.sv:82600:9
				reg_rdata_next[31:0] = cpu_switch_on_counter_qs;
			addr_hit[10]:
				// Trace: design.sv:82604:9
				reg_rdata_next[0] = cpu_wait_ack_switch_on_counter_qs;
			addr_hit[11]:
				// Trace: design.sv:82608:9
				reg_rdata_next[31:0] = cpu_iso_off_counter_qs;
			addr_hit[12]:
				// Trace: design.sv:82612:9
				reg_rdata_next[31:0] = cpu_iso_on_counter_qs;
			addr_hit[13]: begin
				// Trace: design.sv:82616:9
				reg_rdata_next[0] = cpu_counters_stop_cpu_reset_assert_stop_bit_counter_qs;
				// Trace: design.sv:82617:9
				reg_rdata_next[1] = cpu_counters_stop_cpu_reset_deassert_stop_bit_counter_qs;
				// Trace: design.sv:82618:9
				reg_rdata_next[2] = cpu_counters_stop_cpu_switch_off_stop_bit_counter_qs;
				// Trace: design.sv:82619:9
				reg_rdata_next[3] = cpu_counters_stop_cpu_switch_on_stop_bit_counter_qs;
				// Trace: design.sv:82620:9
				reg_rdata_next[4] = cpu_counters_stop_cpu_iso_off_stop_bit_counter_qs;
				// Trace: design.sv:82621:9
				reg_rdata_next[5] = cpu_counters_stop_cpu_iso_on_stop_bit_counter_qs;
			end
			addr_hit[14]:
				// Trace: design.sv:82625:9
				reg_rdata_next[0] = power_gate_periph_ack_qs;
			addr_hit[15]:
				// Trace: design.sv:82629:9
				reg_rdata_next[0] = periph_reset_qs;
			addr_hit[16]:
				// Trace: design.sv:82633:9
				reg_rdata_next[0] = periph_switch_qs;
			addr_hit[17]:
				// Trace: design.sv:82637:9
				reg_rdata_next[0] = periph_wait_ack_switch_on_qs;
			addr_hit[18]:
				// Trace: design.sv:82641:9
				reg_rdata_next[0] = periph_iso_qs;
			addr_hit[19]:
				// Trace: design.sv:82645:9
				reg_rdata_next[0] = periph_clk_gate_qs;
			addr_hit[20]:
				// Trace: design.sv:82649:9
				reg_rdata_next[0] = ram_0_clk_gate_qs;
			addr_hit[21]:
				// Trace: design.sv:82653:9
				reg_rdata_next[0] = power_gate_ram_block_0_ack_qs;
			addr_hit[22]:
				// Trace: design.sv:82657:9
				reg_rdata_next[0] = ram_0_switch_qs;
			addr_hit[23]:
				// Trace: design.sv:82661:9
				reg_rdata_next[0] = ram_0_wait_ack_switch_on_qs;
			addr_hit[24]:
				// Trace: design.sv:82665:9
				reg_rdata_next[0] = ram_0_iso_qs;
			addr_hit[25]:
				// Trace: design.sv:82669:9
				reg_rdata_next[0] = ram_0_retentive_qs;
			addr_hit[26]:
				// Trace: design.sv:82673:9
				reg_rdata_next[0] = ram_1_clk_gate_qs;
			addr_hit[27]:
				// Trace: design.sv:82677:9
				reg_rdata_next[0] = power_gate_ram_block_1_ack_qs;
			addr_hit[28]:
				// Trace: design.sv:82681:9
				reg_rdata_next[0] = ram_1_switch_qs;
			addr_hit[29]:
				// Trace: design.sv:82685:9
				reg_rdata_next[0] = ram_1_wait_ack_switch_on_qs;
			addr_hit[30]:
				// Trace: design.sv:82689:9
				reg_rdata_next[0] = ram_1_iso_qs;
			addr_hit[31]:
				// Trace: design.sv:82693:9
				reg_rdata_next[0] = ram_1_retentive_qs;
			addr_hit[32]:
				// Trace: design.sv:82697:9
				reg_rdata_next[2:0] = monitor_power_gate_core_qs;
			addr_hit[33]:
				// Trace: design.sv:82701:9
				reg_rdata_next[2:0] = monitor_power_gate_periph_qs;
			addr_hit[34]:
				// Trace: design.sv:82705:9
				reg_rdata_next[1:0] = monitor_power_gate_ram_block_0_qs;
			addr_hit[35]:
				// Trace: design.sv:82709:9
				reg_rdata_next[1:0] = monitor_power_gate_ram_block_1_qs;
			addr_hit[36]:
				// Trace: design.sv:82713:9
				reg_rdata_next[0] = master_cpu_force_switch_off_qs;
			addr_hit[37]:
				// Trace: design.sv:82717:9
				reg_rdata_next[0] = master_cpu_force_switch_on_qs;
			addr_hit[38]:
				// Trace: design.sv:82721:9
				reg_rdata_next[0] = master_cpu_force_reset_assert_qs;
			addr_hit[39]:
				// Trace: design.sv:82725:9
				reg_rdata_next[0] = master_cpu_force_reset_deassert_qs;
			addr_hit[40]:
				// Trace: design.sv:82729:9
				reg_rdata_next[0] = master_cpu_force_iso_off_qs;
			addr_hit[41]:
				// Trace: design.sv:82733:9
				reg_rdata_next[0] = master_cpu_force_iso_on_qs;
			default:
				// Trace: design.sv:82737:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:82746:3
	wire unused_wdata;
	// Trace: design.sv:82747:3
	wire unused_be;
	// Trace: design.sv:82748:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:82749:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
// removed module with interface ports: power_manager_reg_top_intf
module power_manager_counter_sequence (
	clk_i,
	rst_ni,
	start_off_sequence_i,
	start_on_sequence_i,
	switch_ack_i,
	counter_expired_switch_off_i,
	counter_expired_switch_on_i,
	counter_start_switch_off_o,
	counter_start_switch_on_o,
	switch_onoff_signal_o
);
	reg _sv2v_0;
	// Trace: design.sv:82813:15
	parameter [0:0] IDLE_VALUE = 1'b1;
	// Trace: design.sv:82815:15
	parameter [0:0] ONOFF_AT_RESET = 1'b1;
	// Trace: design.sv:82817:5
	input wire clk_i;
	// Trace: design.sv:82818:5
	input wire rst_ni;
	// Trace: design.sv:82821:5
	input wire start_off_sequence_i;
	// Trace: design.sv:82822:5
	input wire start_on_sequence_i;
	// Trace: design.sv:82824:5
	input wire switch_ack_i;
	// Trace: design.sv:82827:5
	input wire counter_expired_switch_off_i;
	// Trace: design.sv:82828:5
	input wire counter_expired_switch_on_i;
	// Trace: design.sv:82830:5
	output reg counter_start_switch_off_o;
	// Trace: design.sv:82831:5
	output reg counter_start_switch_on_o;
	// Trace: design.sv:82834:5
	output wire switch_onoff_signal_o;
	// Trace: design.sv:82838:3
	// removed localparam type sequence_fsm_state
	// Trace: design.sv:82848:3
	reg [2:0] sequence_curr_state;
	reg [2:0] sequence_next_state;
	// Trace: design.sv:82850:3
	reg switch_onoff_signal_d;
	reg switch_onoff_signal_q;
	// Trace: design.sv:82853:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_
		// Trace: design.sv:82854:5
		if (~rst_ni) begin
			// Trace: design.sv:82855:7
			sequence_curr_state <= 3'd0;
			// Trace: design.sv:82856:7
			switch_onoff_signal_q <= ONOFF_AT_RESET;
		end
		else begin
			// Trace: design.sv:82858:7
			sequence_curr_state <= sequence_next_state;
			// Trace: design.sv:82859:7
			switch_onoff_signal_q <= switch_onoff_signal_d;
		end
	end
	// Trace: design.sv:82863:3
	assign switch_onoff_signal_o = switch_onoff_signal_q;
	// Trace: design.sv:82866:3
	always @(*) begin : power_manager_counter_sequence_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:82868:5
		sequence_next_state = sequence_curr_state;
		// Trace: design.sv:82869:5
		counter_start_switch_off_o = 1'b0;
		// Trace: design.sv:82870:5
		counter_start_switch_on_o = 1'b0;
		// Trace: design.sv:82871:5
		switch_onoff_signal_d = switch_onoff_signal_q;
		// Trace: design.sv:82873:5
		(* full_case, parallel_case *)
		case (sequence_curr_state)
			3'd0: begin
				// Trace: design.sv:82876:9
				switch_onoff_signal_d = ONOFF_AT_RESET;
				// Trace: design.sv:82877:9
				sequence_next_state = 3'd1;
			end
			3'd1: begin
				// Trace: design.sv:82881:9
				switch_onoff_signal_d = IDLE_VALUE;
				// Trace: design.sv:82882:9
				if (start_off_sequence_i) begin
					// Trace: design.sv:82883:11
					counter_start_switch_off_o = 1'b1;
					// Trace: design.sv:82884:11
					sequence_next_state = 3'd2;
				end
			end
			3'd2: begin
				// Trace: design.sv:82889:9
				switch_onoff_signal_d = IDLE_VALUE;
				// Trace: design.sv:82890:9
				sequence_next_state = (counter_expired_switch_off_i ? 3'd3 : 3'd2);
				// Trace: design.sv:82891:9
				sequence_next_state = (counter_expired_switch_off_i ? 3'd3 : 3'd2);
			end
			3'd3: begin
				// Trace: design.sv:82895:9
				switch_onoff_signal_d = ~IDLE_VALUE;
				// Trace: design.sv:82896:9
				if (start_on_sequence_i) begin
					// Trace: design.sv:82897:11
					counter_start_switch_on_o = 1'b1;
					// Trace: design.sv:82898:11
					sequence_next_state = 3'd4;
				end
			end
			3'd4: begin
				// Trace: design.sv:82903:9
				switch_onoff_signal_d = ~IDLE_VALUE;
				// Trace: design.sv:82904:9
				if (counter_expired_switch_on_i)
					// Trace: design.sv:82905:11
					sequence_next_state = (switch_ack_i ? 3'd6 : 3'd5);
				else
					// Trace: design.sv:82907:11
					sequence_next_state = 3'd4;
			end
			3'd5: begin
				// Trace: design.sv:82912:9
				switch_onoff_signal_d = ~IDLE_VALUE;
				// Trace: design.sv:82913:9
				sequence_next_state = (switch_ack_i ? 3'd6 : 3'd5);
			end
			3'd6: begin
				// Trace: design.sv:82917:9
				switch_onoff_signal_d = IDLE_VALUE;
				// Trace: design.sv:82918:9
				sequence_next_state = 3'd1;
			end
			default:
				// Trace: design.sv:82923:9
				sequence_next_state = 3'd1;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module power_manager_sequence (
	clk_i,
	rst_ni,
	start_off_sequence_i,
	start_on_sequence_i,
	switch_ack_i,
	switch_onoff_signal_o
);
	reg _sv2v_0;
	// Trace: design.sv:82937:15
	parameter [0:0] IDLE_VALUE = 1'b1;
	// Trace: design.sv:82939:15
	parameter [0:0] ONOFF_AT_RESET = 1'b1;
	// Trace: design.sv:82941:5
	input wire clk_i;
	// Trace: design.sv:82942:5
	input wire rst_ni;
	// Trace: design.sv:82945:5
	input wire start_off_sequence_i;
	// Trace: design.sv:82946:5
	input wire start_on_sequence_i;
	// Trace: design.sv:82948:5
	input wire switch_ack_i;
	// Trace: design.sv:82951:5
	output wire switch_onoff_signal_o;
	// Trace: design.sv:82954:3
	// removed localparam type sequence_fsm_state
	// Trace: design.sv:82962:3
	reg [2:0] sequence_curr_state;
	reg [2:0] sequence_next_state;
	// Trace: design.sv:82964:3
	reg switch_onoff_signal_d;
	reg switch_onoff_signal_q;
	// Trace: design.sv:82967:3
	always @(posedge clk_i or negedge rst_ni) begin : proc_
		// Trace: design.sv:82968:5
		if (~rst_ni) begin
			// Trace: design.sv:82969:7
			sequence_curr_state <= 3'd0;
			// Trace: design.sv:82970:7
			switch_onoff_signal_q <= ONOFF_AT_RESET;
		end
		else begin
			// Trace: design.sv:82972:7
			sequence_curr_state <= sequence_next_state;
			// Trace: design.sv:82973:7
			switch_onoff_signal_q <= switch_onoff_signal_d;
		end
	end
	// Trace: design.sv:82977:3
	assign switch_onoff_signal_o = switch_onoff_signal_q;
	// Trace: design.sv:82980:3
	always @(*) begin : power_manager_sequence_fsm
		if (_sv2v_0)
			;
		// Trace: design.sv:82982:5
		sequence_next_state = sequence_curr_state;
		// Trace: design.sv:82983:5
		switch_onoff_signal_d = switch_onoff_signal_q;
		// Trace: design.sv:82985:5
		(* full_case, parallel_case *)
		case (sequence_curr_state)
			3'd0: begin
				// Trace: design.sv:82988:9
				switch_onoff_signal_d = ONOFF_AT_RESET;
				// Trace: design.sv:82989:9
				sequence_next_state = 3'd1;
			end
			3'd1: begin
				// Trace: design.sv:82993:9
				switch_onoff_signal_d = IDLE_VALUE;
				// Trace: design.sv:82994:9
				if (start_off_sequence_i)
					// Trace: design.sv:82995:11
					sequence_next_state = 3'd2;
			end
			3'd2: begin
				// Trace: design.sv:83000:9
				switch_onoff_signal_d = ~IDLE_VALUE;
				// Trace: design.sv:83001:9
				if (start_on_sequence_i)
					// Trace: design.sv:83002:11
					sequence_next_state = 3'd3;
			end
			3'd3: begin
				// Trace: design.sv:83007:9
				switch_onoff_signal_d = ~IDLE_VALUE;
				// Trace: design.sv:83008:9
				if (switch_ack_i)
					// Trace: design.sv:83009:11
					sequence_next_state = 3'd4;
			end
			3'd4: begin
				// Trace: design.sv:83014:9
				switch_onoff_signal_d = IDLE_VALUE;
				// Trace: design.sv:83015:9
				sequence_next_state = 3'd1;
			end
			default:
				// Trace: design.sv:83019:9
				sequence_next_state = 3'd1;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module power_manager_2EE6F (
	clk_i,
	rst_ni,
	reg_req_i,
	reg_rsp_o,
	core_sleep_i,
	intr_i,
	ext_irq_i,
	peripheral_subsystem_clkgate_en_o,
	memory_subsystem_clkgate_en_o,
	cpu_subsystem_powergate_switch_o,
	cpu_subsystem_powergate_switch_ack_i,
	cpu_subsystem_powergate_iso_o,
	cpu_subsystem_rst_no,
	peripheral_subsystem_powergate_switch_o,
	peripheral_subsystem_powergate_switch_ack_i,
	peripheral_subsystem_powergate_iso_o,
	peripheral_subsystem_rst_no,
	memory_subsystem_banks_powergate_switch_o,
	memory_subsystem_banks_powergate_switch_ack_i,
	memory_subsystem_banks_powergate_iso_o,
	memory_subsystem_banks_set_retentive_o,
	external_subsystem_powergate_switch_o,
	external_subsystem_powergate_switch_ack_i,
	external_subsystem_powergate_iso_o,
	external_subsystem_rst_no,
	external_ram_banks_set_retentive_o
);
	reg _sv2v_0;
	// Trace: design.sv:83034:20
	// removed localparam type reg_req_t
	// Trace: design.sv:83035:20
	// removed localparam type reg_rsp_t
	// Trace: design.sv:83036:15
	parameter [0:0] SWITCH_IDLE_VALUE = 1'b1;
	// Trace: design.sv:83037:15
	parameter [0:0] ISO_IDLE_VALUE = 1'b1;
	// Trace: design.sv:83038:15
	parameter [0:0] RESET_IDLE_VALUE = 1'b1;
	// Trace: design.sv:83050:15
	parameter [0:0] SWITCH_VALUE_AT_RESET = SWITCH_IDLE_VALUE;
	// Trace: design.sv:83051:15
	parameter [0:0] ISO_VALUE_AT_RESET = ISO_IDLE_VALUE;
	// Trace: design.sv:83052:15
	parameter [0:0] RESET_VALUE_AT_RESET = ~RESET_IDLE_VALUE;
	// Trace: design.sv:83054:5
	input wire clk_i;
	// Trace: design.sv:83055:5
	input wire rst_ni;
	// Trace: design.sv:83058:5
	input wire [69:0] reg_req_i;
	// Trace: design.sv:83059:5
	output wire [33:0] reg_rsp_o;
	// Trace: design.sv:83062:5
	input wire core_sleep_i;
	// Trace: design.sv:83065:5
	input wire [31:0] intr_i;
	// Trace: design.sv:83068:5
	localparam core_v_mini_mcu_pkg_PLIC_NINT = 64;
	localparam core_v_mini_mcu_pkg_PLIC_USED_NINT = 50;
	localparam core_v_mini_mcu_pkg_NEXT_INT = 14;
	input wire [13:0] ext_irq_i;
	// Trace: design.sv:83071:5
	output wire peripheral_subsystem_clkgate_en_o;
	// Trace: design.sv:83072:5
	localparam [31:0] core_v_mini_mcu_pkg_NUM_BANKS = 2;
	output wire [1:0] memory_subsystem_clkgate_en_o;
	// Trace: design.sv:83075:5
	output wire cpu_subsystem_powergate_switch_o;
	// Trace: design.sv:83076:5
	input wire cpu_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:83077:5
	output wire cpu_subsystem_powergate_iso_o;
	// Trace: design.sv:83078:5
	output wire cpu_subsystem_rst_no;
	// Trace: design.sv:83079:5
	output wire peripheral_subsystem_powergate_switch_o;
	// Trace: design.sv:83080:5
	input wire peripheral_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:83081:5
	output wire peripheral_subsystem_powergate_iso_o;
	// Trace: design.sv:83082:5
	output wire peripheral_subsystem_rst_no;
	// Trace: design.sv:83083:5
	output wire [1:0] memory_subsystem_banks_powergate_switch_o;
	// Trace: design.sv:83084:5
	input wire [1:0] memory_subsystem_banks_powergate_switch_ack_i;
	// Trace: design.sv:83085:5
	output wire [1:0] memory_subsystem_banks_powergate_iso_o;
	// Trace: design.sv:83086:5
	output wire [1:0] memory_subsystem_banks_set_retentive_o;
	// Trace: design.sv:83087:5
	localparam [31:0] core_v_mini_mcu_pkg_EXTERNAL_DOMAINS = 0;
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_switch_o;
	// Trace: design.sv:83088:5
	input wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:83089:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_iso_o;
	// Trace: design.sv:83090:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_rst_no;
	// Trace: design.sv:83091:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_ram_banks_set_retentive_o;
	// Trace: design.sv:83094:3
	// removed import power_manager_reg_pkg::*;
	// Trace: design.sv:83096:3
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_counters_stop_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_iso_off_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_iso_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_reset_assert_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_reset_deassert_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_switch_off_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_switch_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_cpu_wait_ack_switch_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_en_wait_for_intr_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_intr_state_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_iso_off_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_iso_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_reset_assert_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_reset_deassert_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_switch_off_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_master_cpu_force_switch_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_clk_gate_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_iso_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_reset_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_switch_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_periph_wait_ack_switch_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_core_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_core_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_periph_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_ram_block_0_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_power_gate_ram_block_1_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_clk_gate_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_iso_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_retentive_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_switch_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_0_wait_ack_switch_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_clk_gate_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_iso_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_retentive_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_switch_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_ram_1_wait_ack_switch_on_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_restore_address_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_wakeup_state_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_reg2hw_t
	wire [321:0] reg2hw;
	// Trace: design.sv:83097:3
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_iso_off_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_iso_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_reset_assert_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_reset_deassert_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_switch_off_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_cpu_switch_on_counter_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_intr_state_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_monitor_power_gate_core_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_monitor_power_gate_periph_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_monitor_power_gate_ram_block_0_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_monitor_power_gate_ram_block_1_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_power_gate_core_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_power_gate_periph_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_power_gate_ram_block_0_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_power_gate_ram_block_1_ack_reg_t
	// removed localparam type power_manager_reg_pkg_power_manager_hw2reg_t
	wire [252:0] hw2reg;
	// Trace: design.sv:83099:3
	reg start_on_sequence;
	// Trace: design.sv:83101:3
	assign hw2reg[236:221] = {intr_i[29:22], intr_i[21], intr_i[20], intr_i[19], intr_i[18], intr_i[17], intr_i[16], intr_i[11], intr_i[7]};
	// Trace: design.sv:83113:3
	generate
		if (1) begin : genblk1
			// Trace: design.sv:83116:5
			assign hw2reg[252:237] = $unsigned(ext_irq_i);
		end
	endgenerate
	// Trace: design.sv:83119:3
	assign hw2reg[220] = 1'b1;
	// Trace: design.sv:83121:3
	power_manager_reg_top_E039C power_manager_reg_top_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(reg_req_i),
		.reg_rsp_o(reg_rsp_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:83134:3
	wire cpu_subsystem_powergate_switch;
	// Trace: design.sv:83135:3
	wire cpu_subsystem_powergate_iso;
	// Trace: design.sv:83136:3
	wire cpu_subsystem_rst_n;
	// Trace: design.sv:83137:3
	wire peripheral_subsystem_powergate_switch;
	// Trace: design.sv:83138:3
	wire peripheral_subsystem_powergate_iso;
	// Trace: design.sv:83139:3
	wire peripheral_subsystem_rst_n;
	// Trace: design.sv:83140:3
	wire [1:0] memory_subsystem_banks_powergate_switch;
	// Trace: design.sv:83141:3
	wire [1:0] memory_subsystem_banks_powergate_iso;
	// Trace: design.sv:83142:3
	wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_switch;
	// Trace: design.sv:83143:3
	wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_iso;
	// Trace: design.sv:83144:3
	wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_rst_n;
	// Trace: design.sv:83146:3
	assign cpu_subsystem_powergate_switch_o = cpu_subsystem_powergate_switch;
	// Trace: design.sv:83147:3
	assign cpu_subsystem_powergate_iso_o = cpu_subsystem_powergate_iso;
	// Trace: design.sv:83148:3
	assign cpu_subsystem_rst_no = cpu_subsystem_rst_n;
	// Trace: design.sv:83149:3
	assign peripheral_subsystem_powergate_switch_o = peripheral_subsystem_powergate_switch;
	// Trace: design.sv:83150:3
	assign peripheral_subsystem_powergate_iso_o = peripheral_subsystem_powergate_iso;
	// Trace: design.sv:83151:3
	assign peripheral_subsystem_rst_no = peripheral_subsystem_rst_n;
	// Trace: design.sv:83152:3
	assign memory_subsystem_banks_powergate_switch_o = memory_subsystem_banks_powergate_switch;
	// Trace: design.sv:83153:3
	assign memory_subsystem_banks_powergate_iso_o = memory_subsystem_banks_powergate_iso;
	// Trace: design.sv:83154:3
	assign external_subsystem_powergate_switch_o = external_subsystem_powergate_switch;
	// Trace: design.sv:83155:3
	assign external_subsystem_powergate_iso_o = external_subsystem_powergate_iso;
	// Trace: design.sv:83156:3
	assign external_subsystem_rst_no = external_subsystem_rst_n;
	// Trace: design.sv:83162:5
	assign peripheral_subsystem_clkgate_en_o = reg2hw[18];
	// Trace: design.sv:83164:5
	assign memory_subsystem_clkgate_en_o[0] = reg2hw[17];
	// Trace: design.sv:83165:5
	assign memory_subsystem_clkgate_en_o[1] = reg2hw[11];
	// Trace: design.sv:83171:3
	wire cpu_subsystem_powergate_switch_ack_sync;
	// Trace: design.sv:83173:3
	sync #(.ResetValue(1'b0)) sync_cpu_ack_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(cpu_subsystem_powergate_switch_ack_i),
		.serial_o(cpu_subsystem_powergate_switch_ack_sync)
	);
	// Trace: design.sv:83182:3
	assign hw2reg[218] = 1'b1;
	// Trace: design.sv:83183:3
	assign hw2reg[219] = cpu_subsystem_powergate_switch_ack_sync;
	// Trace: design.sv:83186:3
	wire cpu_switch_wait_ack;
	// Trace: design.sv:83187:3
	assign cpu_switch_wait_ack = (reg2hw[94] ? reg2hw[223] == SWITCH_IDLE_VALUE : 1'b1);
	// Trace: design.sv:83189:3
	always @(*) begin : power_manager_start_on_sequence_gen
		if (_sv2v_0)
			;
		// Trace: design.sv:83190:5
		if ((reg2hw[288-:32] & reg2hw[256-:32]) != {32 {1'sb0}})
			// Trace: design.sv:83191:7
			start_on_sequence = 1'b1;
		else
			// Trace: design.sv:83193:7
			start_on_sequence = 1'b0;
	end
	// Trace: design.sv:83197:3
	wire cpu_powergate_counter_start_reset_assert;
	wire cpu_powergate_counter_expired_reset_assert;
	// Trace: design.sv:83198:3
	wire cpu_powergate_counter_start_reset_deassert;
	wire cpu_powergate_counter_expired_reset_deassert;
	// Trace: design.sv:83200:3
	reg_to_counter #(
		.DW(32),
		.ExpireValue(1'sb0)
	) reg_to_counter_cpu_reset_assert_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.stop_i(reg2hw[29]),
		.start_i(cpu_powergate_counter_start_reset_assert),
		.done_o(cpu_powergate_counter_expired_reset_assert),
		.hw2reg_d_o(hw2reg[217-:32]),
		.hw2reg_de_o(hw2reg[185]),
		.hw2reg_q_i(reg2hw[222-:32])
	);
	// Trace: design.sv:83214:3
	reg_to_counter #(
		.DW(32),
		.ExpireValue(1'sb0)
	) reg_to_counter_cpu_reset_deassert_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.stop_i(reg2hw[28]),
		.start_i(cpu_powergate_counter_start_reset_deassert),
		.done_o(cpu_powergate_counter_expired_reset_deassert),
		.hw2reg_d_o(hw2reg[184-:32]),
		.hw2reg_de_o(hw2reg[152]),
		.hw2reg_q_i(reg2hw[190-:32])
	);
	// Trace: design.sv:83228:3
	power_manager_counter_sequence #(
		.IDLE_VALUE(RESET_IDLE_VALUE),
		.ONOFF_AT_RESET(RESET_VALUE_AT_RESET)
	) power_manager_counter_sequence_cpu_reset_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i((reg2hw[224] && core_sleep_i) || reg2hw[3]),
		.start_on_sequence_i(start_on_sequence || reg2hw[2]),
		.switch_ack_i(cpu_switch_wait_ack),
		.counter_expired_switch_off_i(cpu_powergate_counter_expired_reset_assert),
		.counter_expired_switch_on_i(cpu_powergate_counter_expired_reset_deassert),
		.counter_start_switch_off_o(cpu_powergate_counter_start_reset_assert),
		.counter_start_switch_on_o(cpu_powergate_counter_start_reset_deassert),
		.switch_onoff_signal_o(cpu_subsystem_rst_n)
	);
	// Trace: design.sv:83251:3
	wire cpu_powergate_counter_start_switch_off;
	wire cpu_powergate_counter_expired_switch_off;
	// Trace: design.sv:83252:3
	wire cpu_powergate_counter_start_switch_on;
	wire cpu_powergate_counter_expired_switch_on;
	// Trace: design.sv:83254:3
	reg_to_counter #(
		.DW(32),
		.ExpireValue(1'sb0)
	) reg_to_counter_cpu_powergate_switch_off_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.stop_i(reg2hw[27]),
		.start_i(cpu_powergate_counter_start_switch_off),
		.done_o(cpu_powergate_counter_expired_switch_off),
		.hw2reg_d_o(hw2reg[151-:32]),
		.hw2reg_de_o(hw2reg[119]),
		.hw2reg_q_i(reg2hw[158-:32])
	);
	// Trace: design.sv:83268:3
	reg_to_counter #(
		.DW(32),
		.ExpireValue(1'sb0)
	) reg_to_counter_cpu_powergate_switch_on_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.stop_i(reg2hw[26]),
		.start_i(cpu_powergate_counter_start_switch_on),
		.done_o(cpu_powergate_counter_expired_switch_on),
		.hw2reg_d_o(hw2reg[118-:32]),
		.hw2reg_de_o(hw2reg[86]),
		.hw2reg_q_i(reg2hw[126-:32])
	);
	// Trace: design.sv:83282:3
	power_manager_counter_sequence #(
		.IDLE_VALUE(SWITCH_IDLE_VALUE),
		.ONOFF_AT_RESET(SWITCH_VALUE_AT_RESET)
	) power_manager_counter_sequence_cpu_switch_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i((reg2hw[224] && core_sleep_i) || reg2hw[5]),
		.start_on_sequence_i(start_on_sequence || reg2hw[4]),
		.switch_ack_i(1'b1),
		.counter_expired_switch_off_i(cpu_powergate_counter_expired_switch_off),
		.counter_expired_switch_on_i(cpu_powergate_counter_expired_switch_on),
		.counter_start_switch_off_o(cpu_powergate_counter_start_switch_off),
		.counter_start_switch_on_o(cpu_powergate_counter_start_switch_on),
		.switch_onoff_signal_o(cpu_subsystem_powergate_switch)
	);
	// Trace: design.sv:83305:3
	wire cpu_powergate_counter_start_iso_off;
	wire cpu_powergate_counter_expired_iso_off;
	// Trace: design.sv:83306:3
	wire cpu_powergate_counter_start_iso_on;
	wire cpu_powergate_counter_expired_iso_on;
	// Trace: design.sv:83308:3
	reg_to_counter #(
		.DW(32),
		.ExpireValue(1'sb0)
	) reg_to_counter_cpu_powergate_iso_off_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.stop_i(reg2hw[25]),
		.start_i(cpu_powergate_counter_start_iso_off),
		.done_o(cpu_powergate_counter_expired_iso_off),
		.hw2reg_d_o(hw2reg[85-:32]),
		.hw2reg_de_o(hw2reg[53]),
		.hw2reg_q_i(reg2hw[93-:32])
	);
	// Trace: design.sv:83322:3
	reg_to_counter #(
		.DW(32),
		.ExpireValue(1'sb0)
	) reg_to_counter_cpu_powergate_iso_on_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.stop_i(reg2hw[24]),
		.start_i(cpu_powergate_counter_start_iso_on),
		.done_o(cpu_powergate_counter_expired_iso_on),
		.hw2reg_d_o(hw2reg[52-:32]),
		.hw2reg_de_o(hw2reg[20]),
		.hw2reg_q_i(reg2hw[61-:32])
	);
	// Trace: design.sv:83336:3
	power_manager_counter_sequence #(
		.IDLE_VALUE(ISO_IDLE_VALUE),
		.ONOFF_AT_RESET(ISO_VALUE_AT_RESET)
	) power_manager_counter_sequence_cpu_iso_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i((reg2hw[224] && core_sleep_i) || reg2hw[1]),
		.start_on_sequence_i(start_on_sequence || reg2hw[-0]),
		.switch_ack_i(cpu_switch_wait_ack),
		.counter_expired_switch_off_i(cpu_powergate_counter_expired_iso_off),
		.counter_expired_switch_on_i(cpu_powergate_counter_expired_iso_on),
		.counter_start_switch_off_o(cpu_powergate_counter_start_iso_off),
		.counter_start_switch_on_o(cpu_powergate_counter_start_iso_on),
		.switch_onoff_signal_o(cpu_subsystem_powergate_iso)
	);
	// Trace: design.sv:83363:3
	wire peripheral_subsystem_powergate_switch_ack_sync;
	// Trace: design.sv:83365:3
	sync #(.ResetValue(1'b0)) sync_periph_ack_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(peripheral_subsystem_powergate_switch_ack_i),
		.serial_o(peripheral_subsystem_powergate_switch_ack_sync)
	);
	// Trace: design.sv:83374:3
	assign hw2reg[18] = 1'b1;
	// Trace: design.sv:83375:3
	assign hw2reg[19] = peripheral_subsystem_powergate_switch_ack_sync;
	// Trace: design.sv:83378:3
	wire periph_switch_wait_ack;
	// Trace: design.sv:83379:3
	assign periph_switch_wait_ack = (reg2hw[20] ? reg2hw[23] == SWITCH_IDLE_VALUE : 1'b1);
	// Trace: design.sv:83381:3
	power_manager_sequence #(
		.IDLE_VALUE(RESET_IDLE_VALUE),
		.ONOFF_AT_RESET(RESET_VALUE_AT_RESET)
	) power_manager_sequence_periph_reset_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[22]),
		.start_on_sequence_i(~reg2hw[22]),
		.switch_ack_i(periph_switch_wait_ack),
		.switch_onoff_signal_o(peripheral_subsystem_rst_n)
	);
	// Trace: design.sv:83397:3
	power_manager_sequence #(
		.IDLE_VALUE(SWITCH_IDLE_VALUE),
		.ONOFF_AT_RESET(SWITCH_VALUE_AT_RESET)
	) power_manager_sequence_periph_switch_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[21]),
		.start_on_sequence_i(~reg2hw[21]),
		.switch_ack_i(1'b1),
		.switch_onoff_signal_o(peripheral_subsystem_powergate_switch)
	);
	// Trace: design.sv:83413:3
	power_manager_sequence #(
		.IDLE_VALUE(ISO_IDLE_VALUE),
		.ONOFF_AT_RESET(ISO_VALUE_AT_RESET)
	) power_manager_sequence_periph_iso_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[19]),
		.start_on_sequence_i(~reg2hw[19]),
		.switch_ack_i(periph_switch_wait_ack),
		.switch_onoff_signal_o(peripheral_subsystem_powergate_iso)
	);
	// Trace: design.sv:83433:3
	wire ram_0_subsystem_powergate_switch_ack_sync;
	// Trace: design.sv:83435:3
	sync #(.ResetValue(1'b0)) sync_ram_0_ack_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(memory_subsystem_banks_powergate_switch_ack_i[0]),
		.serial_o(ram_0_subsystem_powergate_switch_ack_sync)
	);
	// Trace: design.sv:83444:3
	assign hw2reg[16] = 1'b1;
	// Trace: design.sv:83445:3
	assign hw2reg[17] = ram_0_subsystem_powergate_switch_ack_sync;
	// Trace: design.sv:83448:3
	wire ram_0_switch_wait_ack;
	// Trace: design.sv:83449:3
	assign ram_0_switch_wait_ack = (reg2hw[14] ? reg2hw[16] == SWITCH_IDLE_VALUE : 1'b1);
	// Trace: design.sv:83451:3
	power_manager_sequence #(
		.IDLE_VALUE(SWITCH_IDLE_VALUE),
		.ONOFF_AT_RESET(SWITCH_VALUE_AT_RESET)
	) power_manager_sequence_ram_0_switch_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[15]),
		.start_on_sequence_i(~reg2hw[15]),
		.switch_ack_i(1'b1),
		.switch_onoff_signal_o(memory_subsystem_banks_powergate_switch[0])
	);
	// Trace: design.sv:83467:3
	power_manager_sequence #(
		.IDLE_VALUE(ISO_IDLE_VALUE),
		.ONOFF_AT_RESET(ISO_VALUE_AT_RESET)
	) power_manager_sequence_ram_0_iso_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[13]),
		.start_on_sequence_i(~reg2hw[13]),
		.switch_ack_i(ram_0_switch_wait_ack),
		.switch_onoff_signal_o(memory_subsystem_banks_powergate_iso[0])
	);
	// Trace: design.sv:83483:3
	power_manager_sequence #(
		.IDLE_VALUE(ISO_IDLE_VALUE),
		.ONOFF_AT_RESET(ISO_VALUE_AT_RESET)
	) power_manager_sequence_ram_0_retentive_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[12]),
		.start_on_sequence_i(~reg2hw[12]),
		.switch_ack_i(1'b1),
		.switch_onoff_signal_o(memory_subsystem_banks_set_retentive_o[0])
	);
	// Trace: design.sv:83503:3
	wire ram_1_subsystem_powergate_switch_ack_sync;
	// Trace: design.sv:83505:3
	sync #(.ResetValue(1'b0)) sync_ram_1_ack_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.serial_i(memory_subsystem_banks_powergate_switch_ack_i[1]),
		.serial_o(ram_1_subsystem_powergate_switch_ack_sync)
	);
	// Trace: design.sv:83514:3
	assign hw2reg[14] = 1'b1;
	// Trace: design.sv:83515:3
	assign hw2reg[15] = ram_1_subsystem_powergate_switch_ack_sync;
	// Trace: design.sv:83518:3
	wire ram_1_switch_wait_ack;
	// Trace: design.sv:83519:3
	assign ram_1_switch_wait_ack = (reg2hw[8] ? reg2hw[10] == SWITCH_IDLE_VALUE : 1'b1);
	// Trace: design.sv:83521:3
	power_manager_sequence #(
		.IDLE_VALUE(SWITCH_IDLE_VALUE),
		.ONOFF_AT_RESET(SWITCH_VALUE_AT_RESET)
	) power_manager_sequence_ram_1_switch_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[9]),
		.start_on_sequence_i(~reg2hw[9]),
		.switch_ack_i(1'b1),
		.switch_onoff_signal_o(memory_subsystem_banks_powergate_switch[1])
	);
	// Trace: design.sv:83537:3
	power_manager_sequence #(
		.IDLE_VALUE(ISO_IDLE_VALUE),
		.ONOFF_AT_RESET(ISO_VALUE_AT_RESET)
	) power_manager_sequence_ram_1_iso_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[7]),
		.start_on_sequence_i(~reg2hw[7]),
		.switch_ack_i(ram_1_switch_wait_ack),
		.switch_onoff_signal_o(memory_subsystem_banks_powergate_iso[1])
	);
	// Trace: design.sv:83553:3
	power_manager_sequence #(
		.IDLE_VALUE(ISO_IDLE_VALUE),
		.ONOFF_AT_RESET(ISO_VALUE_AT_RESET)
	) power_manager_sequence_ram_1_retentive_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.start_off_sequence_i(reg2hw[6]),
		.start_on_sequence_i(~reg2hw[6]),
		.switch_ack_i(1'b1),
		.switch_onoff_signal_o(memory_subsystem_banks_set_retentive_o[1])
	);
	// Trace: design.sv:83573:3
	assign hw2reg[10] = 1'b1;
	// Trace: design.sv:83574:3
	assign hw2reg[13-:3] = {cpu_subsystem_rst_n, cpu_subsystem_powergate_iso, cpu_subsystem_powergate_switch};
	// Trace: design.sv:83576:3
	assign hw2reg[6] = 1'b1;
	// Trace: design.sv:83577:3
	assign hw2reg[9-:3] = {peripheral_subsystem_rst_n, peripheral_subsystem_powergate_iso, peripheral_subsystem_powergate_switch};
	// Trace: design.sv:83579:3
	assign hw2reg[3] = 1'b1;
	// Trace: design.sv:83580:3
	assign hw2reg[5-:2] = {memory_subsystem_banks_powergate_iso[0], memory_subsystem_banks_powergate_switch[0]};
	// Trace: design.sv:83582:3
	assign hw2reg[0] = 1'b1;
	// Trace: design.sv:83583:3
	assign hw2reg[2-:2] = {memory_subsystem_banks_powergate_iso[1], memory_subsystem_banks_powergate_switch[1]};
	initial _sv2v_0 = 0;
endmodule
module reg_to_counter (
	clk_i,
	rst_ni,
	stop_i,
	start_i,
	done_o,
	hw2reg_d_o,
	hw2reg_de_o,
	hw2reg_q_i
);
	reg _sv2v_0;
	// Trace: design.sv:83597:15
	parameter signed [31:0] DW = 8;
	// Trace: design.sv:83598:15
	parameter [DW - 1:0] ExpireValue = 1'sb0;
	// Trace: design.sv:83600:5
	input wire clk_i;
	// Trace: design.sv:83601:5
	input wire rst_ni;
	// Trace: design.sv:83603:5
	input wire stop_i;
	// Trace: design.sv:83604:5
	input wire start_i;
	// Trace: design.sv:83605:5
	output reg done_o;
	// Trace: design.sv:83607:5
	output reg [DW - 1:0] hw2reg_d_o;
	// Trace: design.sv:83608:5
	output reg hw2reg_de_o;
	// Trace: design.sv:83610:5
	input wire [DW - 1:0] hw2reg_q_i;
	// Trace: design.sv:83614:3
	// removed localparam type cnt_fsm_state
	// Trace: design.sv:83620:3
	reg [1:0] counter_curr_state;
	reg [1:0] counter_next_state;
	// Trace: design.sv:83622:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:83623:5
		if (~rst_ni)
			// Trace: design.sv:83624:7
			counter_curr_state <= 2'd0;
		else
			// Trace: design.sv:83626:7
			counter_curr_state <= counter_next_state;
	// Trace: design.sv:83631:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:83633:5
		hw2reg_d_o = hw2reg_q_i - 1;
		// Trace: design.sv:83634:5
		hw2reg_de_o = 1'b0;
		// Trace: design.sv:83635:5
		done_o = 1'b0;
		// Trace: design.sv:83636:5
		counter_next_state = counter_curr_state;
		// Trace: design.sv:83638:5
		(* full_case, parallel_case *)
		case (counter_curr_state)
			2'd0: begin
				// Trace: design.sv:83641:9
				hw2reg_de_o = start_i;
				// Trace: design.sv:83642:9
				counter_next_state = (start_i ? 2'd1 : 2'd0);
			end
			2'd1: begin
				// Trace: design.sv:83646:9
				hw2reg_de_o = 1'b1;
				// Trace: design.sv:83647:9
				counter_next_state = (hw2reg_d_o == ExpireValue ? 2'd2 : 2'd1);
			end
			2'd2: begin
				// Trace: design.sv:83651:9
				done_o = 1'b1;
				// Trace: design.sv:83652:9
				counter_next_state = (stop_i ? 2'd0 : 2'd2);
			end
			default:
				// Trace: design.sv:83656:9
				counter_next_state = counter_curr_state;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
module tlul_adapter_reg (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	re_o,
	we_o,
	addr_o,
	wdata_o,
	be_o,
	rdata_i,
	error_i
);
	reg _sv2v_0;
	// removed import tlul_pkg::*;
	// Trace: design.sv:83674:14
	parameter [0:0] EnableDataIntgGen = 1'b0;
	// Trace: design.sv:83675:14
	parameter signed [31:0] RegAw = 8;
	// Trace: design.sv:83676:14
	parameter signed [31:0] RegDw = 32;
	// Trace: design.sv:83677:14
	localparam signed [31:0] RegBw = RegDw / 8;
	// Trace: design.sv:83679:3
	input clk_i;
	// Trace: design.sv:83680:3
	input rst_ni;
	// Trace: design.sv:83683:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:83684:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:83687:3
	output wire re_o;
	// Trace: design.sv:83688:3
	output wire we_o;
	// Trace: design.sv:83689:3
	output wire [RegAw - 1:0] addr_o;
	// Trace: design.sv:83690:3
	output wire [RegDw - 1:0] wdata_o;
	// Trace: design.sv:83691:3
	output wire [RegBw - 1:0] be_o;
	// Trace: design.sv:83692:3
	input [RegDw - 1:0] rdata_i;
	// Trace: design.sv:83693:3
	input error_i;
	// Trace: design.sv:83696:3
	localparam signed [31:0] IW = top_pkg_TL_AIW;
	// Trace: design.sv:83697:3
	localparam signed [31:0] SZW = top_pkg_TL_SZW;
	// Trace: design.sv:83699:3
	reg outstanding;
	// Trace: design.sv:83700:3
	wire a_ack;
	wire d_ack;
	// Trace: design.sv:83702:3
	reg [RegDw - 1:0] rdata;
	// Trace: design.sv:83703:3
	reg error;
	wire err_internal;
	// Trace: design.sv:83705:3
	reg addr_align_err;
	// Trace: design.sv:83706:3
	wire malformed_meta_err;
	// Trace: design.sv:83707:3
	wire tl_err;
	// Trace: design.sv:83709:3
	reg [7:0] reqid;
	// Trace: design.sv:83710:3
	reg [SZW - 1:0] reqsz;
	// Trace: design.sv:83711:3
	reg [2:0] rspop;
	// Trace: design.sv:83713:3
	wire rd_req;
	wire wr_req;
	// Trace: design.sv:83715:3
	assign a_ack = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))] & tl_o[0];
	// Trace: design.sv:83716:3
	assign d_ack = tl_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & tl_i[0];
	// Trace: design.sv:83718:3
	assign wr_req = a_ack & ((tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h0) | (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h1));
	// Trace: design.sv:83719:3
	assign rd_req = a_ack & (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))))) + 1)] == 3'h4);
	// Trace: design.sv:83721:3
	assign we_o = wr_req & ~err_internal;
	// Trace: design.sv:83722:3
	assign re_o = rd_req & ~err_internal;
	// Trace: design.sv:83723:3
	assign wdata_o = tl_i[53-:32];
	// Trace: design.sv:83724:3
	assign be_o = tl_i[top_pkg_TL_DBW + 53-:((top_pkg_TL_DBW + 53) >= 54 ? top_pkg_TL_DBW : 55 - (top_pkg_TL_DBW + 53))];
	// Trace: design.sv:83726:3
	generate
		if (RegAw <= 2) begin : gen_only_one_reg
			// Trace: design.sv:83727:5
			assign addr_o = 1'sb0;
		end
		else begin : gen_more_regs
			// Trace: design.sv:83729:5
			assign addr_o = {tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - (32 - RegAw):(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 29], 2'b00};
		end
	endgenerate
	// Trace: design.sv:83732:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:83733:5
		if (!rst_ni)
			// Trace: design.sv:83733:21
			outstanding <= 1'b0;
		else if (a_ack)
			// Trace: design.sv:83734:21
			outstanding <= 1'b1;
		else if (d_ack)
			// Trace: design.sv:83735:21
			outstanding <= 1'b0;
	// Trace: design.sv:83738:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:83739:5
		if (!rst_ni) begin
			// Trace: design.sv:83740:7
			reqid <= 1'sb0;
			// Trace: design.sv:83741:7
			reqsz <= 1'sb0;
			// Trace: design.sv:83742:7
			rspop <= 3'h0;
		end
		else if (a_ack) begin
			// Trace: design.sv:83744:7
			reqid <= tl_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53)) >= (32'sd32 + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) + 1)];
			// Trace: design.sv:83745:7
			reqsz <= tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 53))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 53))))) + 1)];
			// Trace: design.sv:83747:7
			rspop <= (rd_req ? 3'h1 : 3'h0);
		end
	// Trace: design.sv:83751:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:83752:5
		if (!rst_ni) begin
			// Trace: design.sv:83753:7
			rdata <= 1'sb0;
			// Trace: design.sv:83754:7
			error <= 1'b0;
		end
		else if (a_ack) begin
			// Trace: design.sv:83756:7
			rdata <= ((error_i || err_internal) || wr_req ? {RegDw {1'sb1}} : rdata_i);
			// Trace: design.sv:83757:7
			error <= error_i | err_internal;
		end
	// Trace: design.sv:83761:3
	wire [6:0] data_intg;
	// Trace: design.sv:83762:3
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 57;
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	generate
		if (EnableDataIntgGen) begin : gen_data_intg
			// Trace: design.sv:83763:5
			wire [56:0] unused_data;
			// Trace: design.sv:83765:5
			prim_secded_64_57_enc u_data_gen(
				.in(sv2v_cast_57(rdata)),
				.out({data_intg, unused_data})
			);
		end
		else begin : gen_tieoff_data_intg
			// Trace: design.sv:83770:5
			assign data_intg = 1'sb0;
		end
	endgenerate
	// Trace: design.sv:83773:3
	function automatic [6:0] sv2v_cast_338F4;
		input reg [6:0] inp;
		sv2v_cast_338F4 = inp;
	endfunction
	function automatic [6:0] sv2v_cast_83AAC;
		input reg [6:0] inp;
		sv2v_cast_83AAC = inp;
	endfunction
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_FDEB5;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_FDEB5 = inp;
	endfunction
	function automatic [7:0] sv2v_cast_15E34;
		input reg [7:0] inp;
		sv2v_cast_15E34 = inp;
	endfunction
	function automatic [0:0] sv2v_cast_17D81;
		input reg [0:0] inp;
		sv2v_cast_17D81 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_9783B;
		input reg [31:0] inp;
		sv2v_cast_9783B = inp;
	endfunction
	function automatic [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] sv2v_cast_11E70;
		input reg [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] inp;
		sv2v_cast_11E70 = inp;
	endfunction
	assign tl_o = {outstanding, rspop, 3'b000, sv2v_cast_FDEB5(reqsz), sv2v_cast_15E34(reqid), sv2v_cast_17D81(1'sb0), sv2v_cast_9783B(rdata), sv2v_cast_11E70({sv2v_cast_338F4(1'sb0), sv2v_cast_83AAC(data_intg)}), error, ~outstanding};
	// Trace: design.sv:83789:3
	assign err_internal = (addr_align_err | malformed_meta_err) | tl_err;
	// Trace: design.sv:83792:3
	function automatic tlul_pkg_tl_a_user_chk;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:136:42
		input reg [20:0] user;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:137:5
		reg malformed_err;
		// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:138:5
		reg unused_user;
		begin
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:139:5
			unused_user = |user;
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:140:5
			malformed_err = ~(|{user[15-:2] == 2'b01, user[15-:2] == 2'b10});
			// Trace: ../src/lowrisc_tlul_headers_0.1/rtl/tlul_pkg.sv:141:5
			tlul_pkg_tl_a_user_chk = malformed_err;
		end
	endfunction
	assign malformed_meta_err = tlul_pkg_tl_a_user_chk(tl_i[21-:21]);
	// Trace: design.sv:83798:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:83799:5
		if (wr_req)
			// Trace: design.sv:83801:7
			addr_align_err = |tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 30:(top_pkg_TL_AW + (top_pkg_TL_DBW + 53)) - 31];
		else
			// Trace: design.sv:83804:7
			addr_align_err = 1'b0;
	end
	// Trace: design.sv:83809:3
	tlul_err u_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.err_o(tl_err)
	);
	initial _sv2v_0 = 0;
endmodule
// removed package "i2c_reg_pkg"
module i2c_reg_top (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	reg2hw,
	hw2reg,
	intg_err_o,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:84474:3
	input clk_i;
	// Trace: design.sv:84475:3
	input rst_ni;
	// Trace: design.sv:84477:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:84478:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:84480:3
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_acqdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_fdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_fifo_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_host_timeout_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_enable_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_state_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_test_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_ovrd_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_rdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_stretch_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_target_id_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timeout_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing0_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing1_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing2_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing3_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing4_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_txdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_t
	output wire [388:0] reg2hw;
	// Trace: design.sv:84481:3
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_acqdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_fifo_status_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_intr_state_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_rdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_status_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_val_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_t
	input wire [115:0] hw2reg;
	// Trace: design.sv:84484:3
	output wire intg_err_o;
	// Trace: design.sv:84487:3
	input devmode_i;
	// Trace: design.sv:84490:3
	// removed import i2c_reg_pkg::*;
	// Trace: design.sv:84492:3
	localparam signed [31:0] AW = 7;
	// Trace: design.sv:84493:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:84494:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:84497:3
	wire reg_we;
	// Trace: design.sv:84498:3
	wire reg_re;
	// Trace: design.sv:84499:3
	wire [6:0] reg_addr;
	// Trace: design.sv:84500:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:84501:3
	wire [3:0] reg_be;
	// Trace: design.sv:84502:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:84503:3
	wire reg_error;
	// Trace: design.sv:84505:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:84507:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:84509:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_reg_h2d;
	// Trace: design.sv:84510:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_reg_d2h;
	// Trace: design.sv:84512:3
	assign intg_err_o = 1'sb0;
	// Trace: design.sv:84514:3
	assign tl_reg_h2d = tl_i;
	// Trace: design.sv:84515:3
	assign tl_o = tl_reg_d2h;
	// Trace: design.sv:84517:3
	tlul_adapter_reg #(
		.RegAw(AW),
		.RegDw(DW),
		.EnableDataIntgGen(0)
	) u_reg_if(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_reg_h2d),
		.tl_o(tl_reg_d2h),
		.we_o(reg_we),
		.re_o(reg_re),
		.addr_o(reg_addr),
		.wdata_o(reg_wdata),
		.be_o(reg_be),
		.rdata_i(reg_rdata),
		.error_i(reg_error)
	);
	// Trace: design.sv:84537:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:84538:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:84543:3
	wire intr_state_fmt_watermark_qs;
	// Trace: design.sv:84544:3
	wire intr_state_fmt_watermark_wd;
	// Trace: design.sv:84545:3
	wire intr_state_fmt_watermark_we;
	// Trace: design.sv:84546:3
	wire intr_state_rx_watermark_qs;
	// Trace: design.sv:84547:3
	wire intr_state_rx_watermark_wd;
	// Trace: design.sv:84548:3
	wire intr_state_rx_watermark_we;
	// Trace: design.sv:84549:3
	wire intr_state_fmt_overflow_qs;
	// Trace: design.sv:84550:3
	wire intr_state_fmt_overflow_wd;
	// Trace: design.sv:84551:3
	wire intr_state_fmt_overflow_we;
	// Trace: design.sv:84552:3
	wire intr_state_rx_overflow_qs;
	// Trace: design.sv:84553:3
	wire intr_state_rx_overflow_wd;
	// Trace: design.sv:84554:3
	wire intr_state_rx_overflow_we;
	// Trace: design.sv:84555:3
	wire intr_state_nak_qs;
	// Trace: design.sv:84556:3
	wire intr_state_nak_wd;
	// Trace: design.sv:84557:3
	wire intr_state_nak_we;
	// Trace: design.sv:84558:3
	wire intr_state_scl_interference_qs;
	// Trace: design.sv:84559:3
	wire intr_state_scl_interference_wd;
	// Trace: design.sv:84560:3
	wire intr_state_scl_interference_we;
	// Trace: design.sv:84561:3
	wire intr_state_sda_interference_qs;
	// Trace: design.sv:84562:3
	wire intr_state_sda_interference_wd;
	// Trace: design.sv:84563:3
	wire intr_state_sda_interference_we;
	// Trace: design.sv:84564:3
	wire intr_state_stretch_timeout_qs;
	// Trace: design.sv:84565:3
	wire intr_state_stretch_timeout_wd;
	// Trace: design.sv:84566:3
	wire intr_state_stretch_timeout_we;
	// Trace: design.sv:84567:3
	wire intr_state_sda_unstable_qs;
	// Trace: design.sv:84568:3
	wire intr_state_sda_unstable_wd;
	// Trace: design.sv:84569:3
	wire intr_state_sda_unstable_we;
	// Trace: design.sv:84570:3
	wire intr_state_trans_complete_qs;
	// Trace: design.sv:84571:3
	wire intr_state_trans_complete_wd;
	// Trace: design.sv:84572:3
	wire intr_state_trans_complete_we;
	// Trace: design.sv:84573:3
	wire intr_state_tx_empty_qs;
	// Trace: design.sv:84574:3
	wire intr_state_tx_empty_wd;
	// Trace: design.sv:84575:3
	wire intr_state_tx_empty_we;
	// Trace: design.sv:84576:3
	wire intr_state_tx_nonempty_qs;
	// Trace: design.sv:84577:3
	wire intr_state_tx_nonempty_wd;
	// Trace: design.sv:84578:3
	wire intr_state_tx_nonempty_we;
	// Trace: design.sv:84579:3
	wire intr_state_tx_overflow_qs;
	// Trace: design.sv:84580:3
	wire intr_state_tx_overflow_wd;
	// Trace: design.sv:84581:3
	wire intr_state_tx_overflow_we;
	// Trace: design.sv:84582:3
	wire intr_state_acq_overflow_qs;
	// Trace: design.sv:84583:3
	wire intr_state_acq_overflow_wd;
	// Trace: design.sv:84584:3
	wire intr_state_acq_overflow_we;
	// Trace: design.sv:84585:3
	wire intr_state_ack_stop_qs;
	// Trace: design.sv:84586:3
	wire intr_state_ack_stop_wd;
	// Trace: design.sv:84587:3
	wire intr_state_ack_stop_we;
	// Trace: design.sv:84588:3
	wire intr_state_host_timeout_qs;
	// Trace: design.sv:84589:3
	wire intr_state_host_timeout_wd;
	// Trace: design.sv:84590:3
	wire intr_state_host_timeout_we;
	// Trace: design.sv:84591:3
	wire intr_enable_fmt_watermark_qs;
	// Trace: design.sv:84592:3
	wire intr_enable_fmt_watermark_wd;
	// Trace: design.sv:84593:3
	wire intr_enable_fmt_watermark_we;
	// Trace: design.sv:84594:3
	wire intr_enable_rx_watermark_qs;
	// Trace: design.sv:84595:3
	wire intr_enable_rx_watermark_wd;
	// Trace: design.sv:84596:3
	wire intr_enable_rx_watermark_we;
	// Trace: design.sv:84597:3
	wire intr_enable_fmt_overflow_qs;
	// Trace: design.sv:84598:3
	wire intr_enable_fmt_overflow_wd;
	// Trace: design.sv:84599:3
	wire intr_enable_fmt_overflow_we;
	// Trace: design.sv:84600:3
	wire intr_enable_rx_overflow_qs;
	// Trace: design.sv:84601:3
	wire intr_enable_rx_overflow_wd;
	// Trace: design.sv:84602:3
	wire intr_enable_rx_overflow_we;
	// Trace: design.sv:84603:3
	wire intr_enable_nak_qs;
	// Trace: design.sv:84604:3
	wire intr_enable_nak_wd;
	// Trace: design.sv:84605:3
	wire intr_enable_nak_we;
	// Trace: design.sv:84606:3
	wire intr_enable_scl_interference_qs;
	// Trace: design.sv:84607:3
	wire intr_enable_scl_interference_wd;
	// Trace: design.sv:84608:3
	wire intr_enable_scl_interference_we;
	// Trace: design.sv:84609:3
	wire intr_enable_sda_interference_qs;
	// Trace: design.sv:84610:3
	wire intr_enable_sda_interference_wd;
	// Trace: design.sv:84611:3
	wire intr_enable_sda_interference_we;
	// Trace: design.sv:84612:3
	wire intr_enable_stretch_timeout_qs;
	// Trace: design.sv:84613:3
	wire intr_enable_stretch_timeout_wd;
	// Trace: design.sv:84614:3
	wire intr_enable_stretch_timeout_we;
	// Trace: design.sv:84615:3
	wire intr_enable_sda_unstable_qs;
	// Trace: design.sv:84616:3
	wire intr_enable_sda_unstable_wd;
	// Trace: design.sv:84617:3
	wire intr_enable_sda_unstable_we;
	// Trace: design.sv:84618:3
	wire intr_enable_trans_complete_qs;
	// Trace: design.sv:84619:3
	wire intr_enable_trans_complete_wd;
	// Trace: design.sv:84620:3
	wire intr_enable_trans_complete_we;
	// Trace: design.sv:84621:3
	wire intr_enable_tx_empty_qs;
	// Trace: design.sv:84622:3
	wire intr_enable_tx_empty_wd;
	// Trace: design.sv:84623:3
	wire intr_enable_tx_empty_we;
	// Trace: design.sv:84624:3
	wire intr_enable_tx_nonempty_qs;
	// Trace: design.sv:84625:3
	wire intr_enable_tx_nonempty_wd;
	// Trace: design.sv:84626:3
	wire intr_enable_tx_nonempty_we;
	// Trace: design.sv:84627:3
	wire intr_enable_tx_overflow_qs;
	// Trace: design.sv:84628:3
	wire intr_enable_tx_overflow_wd;
	// Trace: design.sv:84629:3
	wire intr_enable_tx_overflow_we;
	// Trace: design.sv:84630:3
	wire intr_enable_acq_overflow_qs;
	// Trace: design.sv:84631:3
	wire intr_enable_acq_overflow_wd;
	// Trace: design.sv:84632:3
	wire intr_enable_acq_overflow_we;
	// Trace: design.sv:84633:3
	wire intr_enable_ack_stop_qs;
	// Trace: design.sv:84634:3
	wire intr_enable_ack_stop_wd;
	// Trace: design.sv:84635:3
	wire intr_enable_ack_stop_we;
	// Trace: design.sv:84636:3
	wire intr_enable_host_timeout_qs;
	// Trace: design.sv:84637:3
	wire intr_enable_host_timeout_wd;
	// Trace: design.sv:84638:3
	wire intr_enable_host_timeout_we;
	// Trace: design.sv:84639:3
	wire intr_test_fmt_watermark_wd;
	// Trace: design.sv:84640:3
	wire intr_test_fmt_watermark_we;
	// Trace: design.sv:84641:3
	wire intr_test_rx_watermark_wd;
	// Trace: design.sv:84642:3
	wire intr_test_rx_watermark_we;
	// Trace: design.sv:84643:3
	wire intr_test_fmt_overflow_wd;
	// Trace: design.sv:84644:3
	wire intr_test_fmt_overflow_we;
	// Trace: design.sv:84645:3
	wire intr_test_rx_overflow_wd;
	// Trace: design.sv:84646:3
	wire intr_test_rx_overflow_we;
	// Trace: design.sv:84647:3
	wire intr_test_nak_wd;
	// Trace: design.sv:84648:3
	wire intr_test_nak_we;
	// Trace: design.sv:84649:3
	wire intr_test_scl_interference_wd;
	// Trace: design.sv:84650:3
	wire intr_test_scl_interference_we;
	// Trace: design.sv:84651:3
	wire intr_test_sda_interference_wd;
	// Trace: design.sv:84652:3
	wire intr_test_sda_interference_we;
	// Trace: design.sv:84653:3
	wire intr_test_stretch_timeout_wd;
	// Trace: design.sv:84654:3
	wire intr_test_stretch_timeout_we;
	// Trace: design.sv:84655:3
	wire intr_test_sda_unstable_wd;
	// Trace: design.sv:84656:3
	wire intr_test_sda_unstable_we;
	// Trace: design.sv:84657:3
	wire intr_test_trans_complete_wd;
	// Trace: design.sv:84658:3
	wire intr_test_trans_complete_we;
	// Trace: design.sv:84659:3
	wire intr_test_tx_empty_wd;
	// Trace: design.sv:84660:3
	wire intr_test_tx_empty_we;
	// Trace: design.sv:84661:3
	wire intr_test_tx_nonempty_wd;
	// Trace: design.sv:84662:3
	wire intr_test_tx_nonempty_we;
	// Trace: design.sv:84663:3
	wire intr_test_tx_overflow_wd;
	// Trace: design.sv:84664:3
	wire intr_test_tx_overflow_we;
	// Trace: design.sv:84665:3
	wire intr_test_acq_overflow_wd;
	// Trace: design.sv:84666:3
	wire intr_test_acq_overflow_we;
	// Trace: design.sv:84667:3
	wire intr_test_ack_stop_wd;
	// Trace: design.sv:84668:3
	wire intr_test_ack_stop_we;
	// Trace: design.sv:84669:3
	wire intr_test_host_timeout_wd;
	// Trace: design.sv:84670:3
	wire intr_test_host_timeout_we;
	// Trace: design.sv:84671:3
	wire ctrl_enablehost_qs;
	// Trace: design.sv:84672:3
	wire ctrl_enablehost_wd;
	// Trace: design.sv:84673:3
	wire ctrl_enablehost_we;
	// Trace: design.sv:84674:3
	wire ctrl_enabletarget_qs;
	// Trace: design.sv:84675:3
	wire ctrl_enabletarget_wd;
	// Trace: design.sv:84676:3
	wire ctrl_enabletarget_we;
	// Trace: design.sv:84677:3
	wire status_fmtfull_qs;
	// Trace: design.sv:84678:3
	wire status_fmtfull_re;
	// Trace: design.sv:84679:3
	wire status_rxfull_qs;
	// Trace: design.sv:84680:3
	wire status_rxfull_re;
	// Trace: design.sv:84681:3
	wire status_fmtempty_qs;
	// Trace: design.sv:84682:3
	wire status_fmtempty_re;
	// Trace: design.sv:84683:3
	wire status_hostidle_qs;
	// Trace: design.sv:84684:3
	wire status_hostidle_re;
	// Trace: design.sv:84685:3
	wire status_targetidle_qs;
	// Trace: design.sv:84686:3
	wire status_targetidle_re;
	// Trace: design.sv:84687:3
	wire status_rxempty_qs;
	// Trace: design.sv:84688:3
	wire status_rxempty_re;
	// Trace: design.sv:84689:3
	wire status_txfull_qs;
	// Trace: design.sv:84690:3
	wire status_txfull_re;
	// Trace: design.sv:84691:3
	wire status_acqfull_qs;
	// Trace: design.sv:84692:3
	wire status_acqfull_re;
	// Trace: design.sv:84693:3
	wire status_txempty_qs;
	// Trace: design.sv:84694:3
	wire status_txempty_re;
	// Trace: design.sv:84695:3
	wire status_acqempty_qs;
	// Trace: design.sv:84696:3
	wire status_acqempty_re;
	// Trace: design.sv:84697:3
	wire [7:0] rdata_qs;
	// Trace: design.sv:84698:3
	wire rdata_re;
	// Trace: design.sv:84699:3
	wire [7:0] fdata_fbyte_wd;
	// Trace: design.sv:84700:3
	wire fdata_fbyte_we;
	// Trace: design.sv:84701:3
	wire fdata_start_wd;
	// Trace: design.sv:84702:3
	wire fdata_start_we;
	// Trace: design.sv:84703:3
	wire fdata_stop_wd;
	// Trace: design.sv:84704:3
	wire fdata_stop_we;
	// Trace: design.sv:84705:3
	wire fdata_read_wd;
	// Trace: design.sv:84706:3
	wire fdata_read_we;
	// Trace: design.sv:84707:3
	wire fdata_rcont_wd;
	// Trace: design.sv:84708:3
	wire fdata_rcont_we;
	// Trace: design.sv:84709:3
	wire fdata_nakok_wd;
	// Trace: design.sv:84710:3
	wire fdata_nakok_we;
	// Trace: design.sv:84711:3
	wire fifo_ctrl_rxrst_wd;
	// Trace: design.sv:84712:3
	wire fifo_ctrl_rxrst_we;
	// Trace: design.sv:84713:3
	wire fifo_ctrl_fmtrst_wd;
	// Trace: design.sv:84714:3
	wire fifo_ctrl_fmtrst_we;
	// Trace: design.sv:84715:3
	wire [2:0] fifo_ctrl_rxilvl_qs;
	// Trace: design.sv:84716:3
	wire [2:0] fifo_ctrl_rxilvl_wd;
	// Trace: design.sv:84717:3
	wire fifo_ctrl_rxilvl_we;
	// Trace: design.sv:84718:3
	wire [1:0] fifo_ctrl_fmtilvl_qs;
	// Trace: design.sv:84719:3
	wire [1:0] fifo_ctrl_fmtilvl_wd;
	// Trace: design.sv:84720:3
	wire fifo_ctrl_fmtilvl_we;
	// Trace: design.sv:84721:3
	wire fifo_ctrl_acqrst_wd;
	// Trace: design.sv:84722:3
	wire fifo_ctrl_acqrst_we;
	// Trace: design.sv:84723:3
	wire fifo_ctrl_txrst_wd;
	// Trace: design.sv:84724:3
	wire fifo_ctrl_txrst_we;
	// Trace: design.sv:84725:3
	wire [5:0] fifo_status_fmtlvl_qs;
	// Trace: design.sv:84726:3
	wire fifo_status_fmtlvl_re;
	// Trace: design.sv:84727:3
	wire [5:0] fifo_status_txlvl_qs;
	// Trace: design.sv:84728:3
	wire fifo_status_txlvl_re;
	// Trace: design.sv:84729:3
	wire [5:0] fifo_status_rxlvl_qs;
	// Trace: design.sv:84730:3
	wire fifo_status_rxlvl_re;
	// Trace: design.sv:84731:3
	wire [5:0] fifo_status_acqlvl_qs;
	// Trace: design.sv:84732:3
	wire fifo_status_acqlvl_re;
	// Trace: design.sv:84733:3
	wire ovrd_txovrden_qs;
	// Trace: design.sv:84734:3
	wire ovrd_txovrden_wd;
	// Trace: design.sv:84735:3
	wire ovrd_txovrden_we;
	// Trace: design.sv:84736:3
	wire ovrd_sclval_qs;
	// Trace: design.sv:84737:3
	wire ovrd_sclval_wd;
	// Trace: design.sv:84738:3
	wire ovrd_sclval_we;
	// Trace: design.sv:84739:3
	wire ovrd_sdaval_qs;
	// Trace: design.sv:84740:3
	wire ovrd_sdaval_wd;
	// Trace: design.sv:84741:3
	wire ovrd_sdaval_we;
	// Trace: design.sv:84742:3
	wire [15:0] val_scl_rx_qs;
	// Trace: design.sv:84743:3
	wire val_scl_rx_re;
	// Trace: design.sv:84744:3
	wire [15:0] val_sda_rx_qs;
	// Trace: design.sv:84745:3
	wire val_sda_rx_re;
	// Trace: design.sv:84746:3
	wire [15:0] timing0_thigh_qs;
	// Trace: design.sv:84747:3
	wire [15:0] timing0_thigh_wd;
	// Trace: design.sv:84748:3
	wire timing0_thigh_we;
	// Trace: design.sv:84749:3
	wire [15:0] timing0_tlow_qs;
	// Trace: design.sv:84750:3
	wire [15:0] timing0_tlow_wd;
	// Trace: design.sv:84751:3
	wire timing0_tlow_we;
	// Trace: design.sv:84752:3
	wire [15:0] timing1_t_r_qs;
	// Trace: design.sv:84753:3
	wire [15:0] timing1_t_r_wd;
	// Trace: design.sv:84754:3
	wire timing1_t_r_we;
	// Trace: design.sv:84755:3
	wire [15:0] timing1_t_f_qs;
	// Trace: design.sv:84756:3
	wire [15:0] timing1_t_f_wd;
	// Trace: design.sv:84757:3
	wire timing1_t_f_we;
	// Trace: design.sv:84758:3
	wire [15:0] timing2_tsu_sta_qs;
	// Trace: design.sv:84759:3
	wire [15:0] timing2_tsu_sta_wd;
	// Trace: design.sv:84760:3
	wire timing2_tsu_sta_we;
	// Trace: design.sv:84761:3
	wire [15:0] timing2_thd_sta_qs;
	// Trace: design.sv:84762:3
	wire [15:0] timing2_thd_sta_wd;
	// Trace: design.sv:84763:3
	wire timing2_thd_sta_we;
	// Trace: design.sv:84764:3
	wire [15:0] timing3_tsu_dat_qs;
	// Trace: design.sv:84765:3
	wire [15:0] timing3_tsu_dat_wd;
	// Trace: design.sv:84766:3
	wire timing3_tsu_dat_we;
	// Trace: design.sv:84767:3
	wire [15:0] timing3_thd_dat_qs;
	// Trace: design.sv:84768:3
	wire [15:0] timing3_thd_dat_wd;
	// Trace: design.sv:84769:3
	wire timing3_thd_dat_we;
	// Trace: design.sv:84770:3
	wire [15:0] timing4_tsu_sto_qs;
	// Trace: design.sv:84771:3
	wire [15:0] timing4_tsu_sto_wd;
	// Trace: design.sv:84772:3
	wire timing4_tsu_sto_we;
	// Trace: design.sv:84773:3
	wire [15:0] timing4_t_buf_qs;
	// Trace: design.sv:84774:3
	wire [15:0] timing4_t_buf_wd;
	// Trace: design.sv:84775:3
	wire timing4_t_buf_we;
	// Trace: design.sv:84776:3
	wire [30:0] timeout_ctrl_val_qs;
	// Trace: design.sv:84777:3
	wire [30:0] timeout_ctrl_val_wd;
	// Trace: design.sv:84778:3
	wire timeout_ctrl_val_we;
	// Trace: design.sv:84779:3
	wire timeout_ctrl_en_qs;
	// Trace: design.sv:84780:3
	wire timeout_ctrl_en_wd;
	// Trace: design.sv:84781:3
	wire timeout_ctrl_en_we;
	// Trace: design.sv:84782:3
	wire [6:0] target_id_address0_qs;
	// Trace: design.sv:84783:3
	wire [6:0] target_id_address0_wd;
	// Trace: design.sv:84784:3
	wire target_id_address0_we;
	// Trace: design.sv:84785:3
	wire [6:0] target_id_mask0_qs;
	// Trace: design.sv:84786:3
	wire [6:0] target_id_mask0_wd;
	// Trace: design.sv:84787:3
	wire target_id_mask0_we;
	// Trace: design.sv:84788:3
	wire [6:0] target_id_address1_qs;
	// Trace: design.sv:84789:3
	wire [6:0] target_id_address1_wd;
	// Trace: design.sv:84790:3
	wire target_id_address1_we;
	// Trace: design.sv:84791:3
	wire [6:0] target_id_mask1_qs;
	// Trace: design.sv:84792:3
	wire [6:0] target_id_mask1_wd;
	// Trace: design.sv:84793:3
	wire target_id_mask1_we;
	// Trace: design.sv:84794:3
	wire [7:0] acqdata_abyte_qs;
	// Trace: design.sv:84795:3
	wire acqdata_abyte_re;
	// Trace: design.sv:84796:3
	wire [1:0] acqdata_signal_qs;
	// Trace: design.sv:84797:3
	wire acqdata_signal_re;
	// Trace: design.sv:84798:3
	wire [7:0] txdata_wd;
	// Trace: design.sv:84799:3
	wire txdata_we;
	// Trace: design.sv:84800:3
	wire stretch_ctrl_enableaddr_qs;
	// Trace: design.sv:84801:3
	wire stretch_ctrl_enableaddr_wd;
	// Trace: design.sv:84802:3
	wire stretch_ctrl_enableaddr_we;
	// Trace: design.sv:84803:3
	wire stretch_ctrl_enabletx_qs;
	// Trace: design.sv:84804:3
	wire stretch_ctrl_enabletx_wd;
	// Trace: design.sv:84805:3
	wire stretch_ctrl_enabletx_we;
	// Trace: design.sv:84806:3
	wire stretch_ctrl_enableacq_qs;
	// Trace: design.sv:84807:3
	wire stretch_ctrl_enableacq_wd;
	// Trace: design.sv:84808:3
	wire stretch_ctrl_enableacq_we;
	// Trace: design.sv:84809:3
	wire stretch_ctrl_stop_qs;
	// Trace: design.sv:84810:3
	wire stretch_ctrl_stop_wd;
	// Trace: design.sv:84811:3
	wire stretch_ctrl_stop_we;
	// Trace: design.sv:84812:3
	wire [31:0] host_timeout_ctrl_qs;
	// Trace: design.sv:84813:3
	wire [31:0] host_timeout_ctrl_wd;
	// Trace: design.sv:84814:3
	wire host_timeout_ctrl_we;
	// Trace: design.sv:84820:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_fmt_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_fmt_watermark_we),
		.wd(intr_state_fmt_watermark_wd),
		.de(hw2reg[114]),
		.d(hw2reg[115]),
		.qe(),
		.q(reg2hw[388]),
		.qs(intr_state_fmt_watermark_qs)
	);
	// Trace: design.sv:84846:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_rx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_rx_watermark_we),
		.wd(intr_state_rx_watermark_wd),
		.de(hw2reg[112]),
		.d(hw2reg[113]),
		.qe(),
		.q(reg2hw[387]),
		.qs(intr_state_rx_watermark_qs)
	);
	// Trace: design.sv:84872:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_fmt_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_fmt_overflow_we),
		.wd(intr_state_fmt_overflow_wd),
		.de(hw2reg[110]),
		.d(hw2reg[111]),
		.qe(),
		.q(reg2hw[386]),
		.qs(intr_state_fmt_overflow_qs)
	);
	// Trace: design.sv:84898:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_rx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_rx_overflow_we),
		.wd(intr_state_rx_overflow_wd),
		.de(hw2reg[108]),
		.d(hw2reg[109]),
		.qe(),
		.q(reg2hw[385]),
		.qs(intr_state_rx_overflow_qs)
	);
	// Trace: design.sv:84924:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_nak(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_nak_we),
		.wd(intr_state_nak_wd),
		.de(hw2reg[106]),
		.d(hw2reg[107]),
		.qe(),
		.q(reg2hw[384]),
		.qs(intr_state_nak_qs)
	);
	// Trace: design.sv:84950:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_scl_interference(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_scl_interference_we),
		.wd(intr_state_scl_interference_wd),
		.de(hw2reg[104]),
		.d(hw2reg[105]),
		.qe(),
		.q(reg2hw[383]),
		.qs(intr_state_scl_interference_qs)
	);
	// Trace: design.sv:84976:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_sda_interference(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_sda_interference_we),
		.wd(intr_state_sda_interference_wd),
		.de(hw2reg[102]),
		.d(hw2reg[103]),
		.qe(),
		.q(reg2hw[382]),
		.qs(intr_state_sda_interference_qs)
	);
	// Trace: design.sv:85002:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_stretch_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_stretch_timeout_we),
		.wd(intr_state_stretch_timeout_wd),
		.de(hw2reg[100]),
		.d(hw2reg[101]),
		.qe(),
		.q(reg2hw[381]),
		.qs(intr_state_stretch_timeout_qs)
	);
	// Trace: design.sv:85028:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_sda_unstable(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_sda_unstable_we),
		.wd(intr_state_sda_unstable_wd),
		.de(hw2reg[98]),
		.d(hw2reg[99]),
		.qe(),
		.q(reg2hw[380]),
		.qs(intr_state_sda_unstable_qs)
	);
	// Trace: design.sv:85054:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_trans_complete(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_trans_complete_we),
		.wd(intr_state_trans_complete_wd),
		.de(hw2reg[96]),
		.d(hw2reg[97]),
		.qe(),
		.q(reg2hw[379]),
		.qs(intr_state_trans_complete_qs)
	);
	// Trace: design.sv:85080:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_tx_empty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_tx_empty_we),
		.wd(intr_state_tx_empty_wd),
		.de(hw2reg[94]),
		.d(hw2reg[95]),
		.qe(),
		.q(reg2hw[378]),
		.qs(intr_state_tx_empty_qs)
	);
	// Trace: design.sv:85106:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_tx_nonempty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_tx_nonempty_we),
		.wd(intr_state_tx_nonempty_wd),
		.de(hw2reg[92]),
		.d(hw2reg[93]),
		.qe(),
		.q(reg2hw[377]),
		.qs(intr_state_tx_nonempty_qs)
	);
	// Trace: design.sv:85132:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_tx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_tx_overflow_we),
		.wd(intr_state_tx_overflow_wd),
		.de(hw2reg[90]),
		.d(hw2reg[91]),
		.qe(),
		.q(reg2hw[376]),
		.qs(intr_state_tx_overflow_qs)
	);
	// Trace: design.sv:85158:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_acq_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_acq_overflow_we),
		.wd(intr_state_acq_overflow_wd),
		.de(hw2reg[88]),
		.d(hw2reg[89]),
		.qe(),
		.q(reg2hw[375]),
		.qs(intr_state_acq_overflow_qs)
	);
	// Trace: design.sv:85184:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_ack_stop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_ack_stop_we),
		.wd(intr_state_ack_stop_wd),
		.de(hw2reg[86]),
		.d(hw2reg[87]),
		.qe(),
		.q(reg2hw[374]),
		.qs(intr_state_ack_stop_qs)
	);
	// Trace: design.sv:85210:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_host_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_host_timeout_we),
		.wd(intr_state_host_timeout_wd),
		.de(hw2reg[84]),
		.d(hw2reg[85]),
		.qe(),
		.q(reg2hw[373]),
		.qs(intr_state_host_timeout_qs)
	);
	// Trace: design.sv:85238:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_fmt_watermark_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_fmt_watermark_d
	localparam [0:0] sv2v_uu_u_intr_enable_fmt_watermark_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_fmt_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_fmt_watermark_we),
		.wd(intr_enable_fmt_watermark_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_fmt_watermark_ext_d_0),
		.qe(),
		.q(reg2hw[372]),
		.qs(intr_enable_fmt_watermark_qs)
	);
	// Trace: design.sv:85264:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_rx_watermark_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_rx_watermark_d
	localparam [0:0] sv2v_uu_u_intr_enable_rx_watermark_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_rx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_rx_watermark_we),
		.wd(intr_enable_rx_watermark_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_rx_watermark_ext_d_0),
		.qe(),
		.q(reg2hw[371]),
		.qs(intr_enable_rx_watermark_qs)
	);
	// Trace: design.sv:85290:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_fmt_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_fmt_overflow_d
	localparam [0:0] sv2v_uu_u_intr_enable_fmt_overflow_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_fmt_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_fmt_overflow_we),
		.wd(intr_enable_fmt_overflow_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_fmt_overflow_ext_d_0),
		.qe(),
		.q(reg2hw[370]),
		.qs(intr_enable_fmt_overflow_qs)
	);
	// Trace: design.sv:85316:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_rx_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_rx_overflow_d
	localparam [0:0] sv2v_uu_u_intr_enable_rx_overflow_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_rx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_rx_overflow_we),
		.wd(intr_enable_rx_overflow_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_rx_overflow_ext_d_0),
		.qe(),
		.q(reg2hw[369]),
		.qs(intr_enable_rx_overflow_qs)
	);
	// Trace: design.sv:85342:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_nak_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_nak_d
	localparam [0:0] sv2v_uu_u_intr_enable_nak_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_nak(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_nak_we),
		.wd(intr_enable_nak_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_nak_ext_d_0),
		.qe(),
		.q(reg2hw[368]),
		.qs(intr_enable_nak_qs)
	);
	// Trace: design.sv:85368:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_scl_interference_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_scl_interference_d
	localparam [0:0] sv2v_uu_u_intr_enable_scl_interference_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_scl_interference(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_scl_interference_we),
		.wd(intr_enable_scl_interference_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_scl_interference_ext_d_0),
		.qe(),
		.q(reg2hw[367]),
		.qs(intr_enable_scl_interference_qs)
	);
	// Trace: design.sv:85394:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_sda_interference_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_sda_interference_d
	localparam [0:0] sv2v_uu_u_intr_enable_sda_interference_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_sda_interference(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_sda_interference_we),
		.wd(intr_enable_sda_interference_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_sda_interference_ext_d_0),
		.qe(),
		.q(reg2hw[366]),
		.qs(intr_enable_sda_interference_qs)
	);
	// Trace: design.sv:85420:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_stretch_timeout_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_stretch_timeout_d
	localparam [0:0] sv2v_uu_u_intr_enable_stretch_timeout_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_stretch_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_stretch_timeout_we),
		.wd(intr_enable_stretch_timeout_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_stretch_timeout_ext_d_0),
		.qe(),
		.q(reg2hw[365]),
		.qs(intr_enable_stretch_timeout_qs)
	);
	// Trace: design.sv:85446:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_sda_unstable_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_sda_unstable_d
	localparam [0:0] sv2v_uu_u_intr_enable_sda_unstable_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_sda_unstable(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_sda_unstable_we),
		.wd(intr_enable_sda_unstable_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_sda_unstable_ext_d_0),
		.qe(),
		.q(reg2hw[364]),
		.qs(intr_enable_sda_unstable_qs)
	);
	// Trace: design.sv:85472:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_trans_complete_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_trans_complete_d
	localparam [0:0] sv2v_uu_u_intr_enable_trans_complete_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_trans_complete(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_trans_complete_we),
		.wd(intr_enable_trans_complete_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_trans_complete_ext_d_0),
		.qe(),
		.q(reg2hw[363]),
		.qs(intr_enable_trans_complete_qs)
	);
	// Trace: design.sv:85498:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_tx_empty_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_tx_empty_d
	localparam [0:0] sv2v_uu_u_intr_enable_tx_empty_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_tx_empty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_tx_empty_we),
		.wd(intr_enable_tx_empty_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_tx_empty_ext_d_0),
		.qe(),
		.q(reg2hw[362]),
		.qs(intr_enable_tx_empty_qs)
	);
	// Trace: design.sv:85524:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_tx_nonempty_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_tx_nonempty_d
	localparam [0:0] sv2v_uu_u_intr_enable_tx_nonempty_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_tx_nonempty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_tx_nonempty_we),
		.wd(intr_enable_tx_nonempty_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_tx_nonempty_ext_d_0),
		.qe(),
		.q(reg2hw[361]),
		.qs(intr_enable_tx_nonempty_qs)
	);
	// Trace: design.sv:85550:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_tx_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_tx_overflow_d
	localparam [0:0] sv2v_uu_u_intr_enable_tx_overflow_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_tx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_tx_overflow_we),
		.wd(intr_enable_tx_overflow_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_tx_overflow_ext_d_0),
		.qe(),
		.q(reg2hw[360]),
		.qs(intr_enable_tx_overflow_qs)
	);
	// Trace: design.sv:85576:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_acq_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_acq_overflow_d
	localparam [0:0] sv2v_uu_u_intr_enable_acq_overflow_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_acq_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_acq_overflow_we),
		.wd(intr_enable_acq_overflow_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_acq_overflow_ext_d_0),
		.qe(),
		.q(reg2hw[359]),
		.qs(intr_enable_acq_overflow_qs)
	);
	// Trace: design.sv:85602:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_ack_stop_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_ack_stop_d
	localparam [0:0] sv2v_uu_u_intr_enable_ack_stop_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_ack_stop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_ack_stop_we),
		.wd(intr_enable_ack_stop_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_ack_stop_ext_d_0),
		.qe(),
		.q(reg2hw[358]),
		.qs(intr_enable_ack_stop_qs)
	);
	// Trace: design.sv:85628:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_host_timeout_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_host_timeout_d
	localparam [0:0] sv2v_uu_u_intr_enable_host_timeout_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_host_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_host_timeout_we),
		.wd(intr_enable_host_timeout_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_host_timeout_ext_d_0),
		.qe(),
		.q(reg2hw[357]),
		.qs(intr_enable_host_timeout_qs)
	);
	// Trace: design.sv:85656:3
	localparam [31:0] sv2v_uu_u_intr_test_fmt_watermark_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_fmt_watermark_d
	localparam [0:0] sv2v_uu_u_intr_test_fmt_watermark_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_fmt_watermark(
		.re(1'b0),
		.we(intr_test_fmt_watermark_we),
		.wd(intr_test_fmt_watermark_wd),
		.d(sv2v_uu_u_intr_test_fmt_watermark_ext_d_0),
		.qre(),
		.qe(reg2hw[355]),
		.q(reg2hw[356]),
		.qs()
	);
	// Trace: design.sv:85671:3
	localparam [31:0] sv2v_uu_u_intr_test_rx_watermark_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_rx_watermark_d
	localparam [0:0] sv2v_uu_u_intr_test_rx_watermark_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_rx_watermark(
		.re(1'b0),
		.we(intr_test_rx_watermark_we),
		.wd(intr_test_rx_watermark_wd),
		.d(sv2v_uu_u_intr_test_rx_watermark_ext_d_0),
		.qre(),
		.qe(reg2hw[353]),
		.q(reg2hw[354]),
		.qs()
	);
	// Trace: design.sv:85686:3
	localparam [31:0] sv2v_uu_u_intr_test_fmt_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_fmt_overflow_d
	localparam [0:0] sv2v_uu_u_intr_test_fmt_overflow_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_fmt_overflow(
		.re(1'b0),
		.we(intr_test_fmt_overflow_we),
		.wd(intr_test_fmt_overflow_wd),
		.d(sv2v_uu_u_intr_test_fmt_overflow_ext_d_0),
		.qre(),
		.qe(reg2hw[351]),
		.q(reg2hw[352]),
		.qs()
	);
	// Trace: design.sv:85701:3
	localparam [31:0] sv2v_uu_u_intr_test_rx_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_rx_overflow_d
	localparam [0:0] sv2v_uu_u_intr_test_rx_overflow_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_rx_overflow(
		.re(1'b0),
		.we(intr_test_rx_overflow_we),
		.wd(intr_test_rx_overflow_wd),
		.d(sv2v_uu_u_intr_test_rx_overflow_ext_d_0),
		.qre(),
		.qe(reg2hw[349]),
		.q(reg2hw[350]),
		.qs()
	);
	// Trace: design.sv:85716:3
	localparam [31:0] sv2v_uu_u_intr_test_nak_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_nak_d
	localparam [0:0] sv2v_uu_u_intr_test_nak_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_nak(
		.re(1'b0),
		.we(intr_test_nak_we),
		.wd(intr_test_nak_wd),
		.d(sv2v_uu_u_intr_test_nak_ext_d_0),
		.qre(),
		.qe(reg2hw[347]),
		.q(reg2hw[348]),
		.qs()
	);
	// Trace: design.sv:85731:3
	localparam [31:0] sv2v_uu_u_intr_test_scl_interference_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_scl_interference_d
	localparam [0:0] sv2v_uu_u_intr_test_scl_interference_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_scl_interference(
		.re(1'b0),
		.we(intr_test_scl_interference_we),
		.wd(intr_test_scl_interference_wd),
		.d(sv2v_uu_u_intr_test_scl_interference_ext_d_0),
		.qre(),
		.qe(reg2hw[345]),
		.q(reg2hw[346]),
		.qs()
	);
	// Trace: design.sv:85746:3
	localparam [31:0] sv2v_uu_u_intr_test_sda_interference_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_sda_interference_d
	localparam [0:0] sv2v_uu_u_intr_test_sda_interference_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_sda_interference(
		.re(1'b0),
		.we(intr_test_sda_interference_we),
		.wd(intr_test_sda_interference_wd),
		.d(sv2v_uu_u_intr_test_sda_interference_ext_d_0),
		.qre(),
		.qe(reg2hw[343]),
		.q(reg2hw[344]),
		.qs()
	);
	// Trace: design.sv:85761:3
	localparam [31:0] sv2v_uu_u_intr_test_stretch_timeout_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_stretch_timeout_d
	localparam [0:0] sv2v_uu_u_intr_test_stretch_timeout_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_stretch_timeout(
		.re(1'b0),
		.we(intr_test_stretch_timeout_we),
		.wd(intr_test_stretch_timeout_wd),
		.d(sv2v_uu_u_intr_test_stretch_timeout_ext_d_0),
		.qre(),
		.qe(reg2hw[341]),
		.q(reg2hw[342]),
		.qs()
	);
	// Trace: design.sv:85776:3
	localparam [31:0] sv2v_uu_u_intr_test_sda_unstable_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_sda_unstable_d
	localparam [0:0] sv2v_uu_u_intr_test_sda_unstable_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_sda_unstable(
		.re(1'b0),
		.we(intr_test_sda_unstable_we),
		.wd(intr_test_sda_unstable_wd),
		.d(sv2v_uu_u_intr_test_sda_unstable_ext_d_0),
		.qre(),
		.qe(reg2hw[339]),
		.q(reg2hw[340]),
		.qs()
	);
	// Trace: design.sv:85791:3
	localparam [31:0] sv2v_uu_u_intr_test_trans_complete_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_trans_complete_d
	localparam [0:0] sv2v_uu_u_intr_test_trans_complete_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_trans_complete(
		.re(1'b0),
		.we(intr_test_trans_complete_we),
		.wd(intr_test_trans_complete_wd),
		.d(sv2v_uu_u_intr_test_trans_complete_ext_d_0),
		.qre(),
		.qe(reg2hw[337]),
		.q(reg2hw[338]),
		.qs()
	);
	// Trace: design.sv:85806:3
	localparam [31:0] sv2v_uu_u_intr_test_tx_empty_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_tx_empty_d
	localparam [0:0] sv2v_uu_u_intr_test_tx_empty_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_tx_empty(
		.re(1'b0),
		.we(intr_test_tx_empty_we),
		.wd(intr_test_tx_empty_wd),
		.d(sv2v_uu_u_intr_test_tx_empty_ext_d_0),
		.qre(),
		.qe(reg2hw[335]),
		.q(reg2hw[336]),
		.qs()
	);
	// Trace: design.sv:85821:3
	localparam [31:0] sv2v_uu_u_intr_test_tx_nonempty_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_tx_nonempty_d
	localparam [0:0] sv2v_uu_u_intr_test_tx_nonempty_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_tx_nonempty(
		.re(1'b0),
		.we(intr_test_tx_nonempty_we),
		.wd(intr_test_tx_nonempty_wd),
		.d(sv2v_uu_u_intr_test_tx_nonempty_ext_d_0),
		.qre(),
		.qe(reg2hw[333]),
		.q(reg2hw[334]),
		.qs()
	);
	// Trace: design.sv:85836:3
	localparam [31:0] sv2v_uu_u_intr_test_tx_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_tx_overflow_d
	localparam [0:0] sv2v_uu_u_intr_test_tx_overflow_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_tx_overflow(
		.re(1'b0),
		.we(intr_test_tx_overflow_we),
		.wd(intr_test_tx_overflow_wd),
		.d(sv2v_uu_u_intr_test_tx_overflow_ext_d_0),
		.qre(),
		.qe(reg2hw[331]),
		.q(reg2hw[332]),
		.qs()
	);
	// Trace: design.sv:85851:3
	localparam [31:0] sv2v_uu_u_intr_test_acq_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_acq_overflow_d
	localparam [0:0] sv2v_uu_u_intr_test_acq_overflow_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_acq_overflow(
		.re(1'b0),
		.we(intr_test_acq_overflow_we),
		.wd(intr_test_acq_overflow_wd),
		.d(sv2v_uu_u_intr_test_acq_overflow_ext_d_0),
		.qre(),
		.qe(reg2hw[329]),
		.q(reg2hw[330]),
		.qs()
	);
	// Trace: design.sv:85866:3
	localparam [31:0] sv2v_uu_u_intr_test_ack_stop_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_ack_stop_d
	localparam [0:0] sv2v_uu_u_intr_test_ack_stop_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_ack_stop(
		.re(1'b0),
		.we(intr_test_ack_stop_we),
		.wd(intr_test_ack_stop_wd),
		.d(sv2v_uu_u_intr_test_ack_stop_ext_d_0),
		.qre(),
		.qe(reg2hw[327]),
		.q(reg2hw[328]),
		.qs()
	);
	// Trace: design.sv:85881:3
	localparam [31:0] sv2v_uu_u_intr_test_host_timeout_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_host_timeout_d
	localparam [0:0] sv2v_uu_u_intr_test_host_timeout_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_host_timeout(
		.re(1'b0),
		.we(intr_test_host_timeout_we),
		.wd(intr_test_host_timeout_wd),
		.d(sv2v_uu_u_intr_test_host_timeout_ext_d_0),
		.qre(),
		.qe(reg2hw[325]),
		.q(reg2hw[326]),
		.qs()
	);
	// Trace: design.sv:85898:3
	localparam signed [31:0] sv2v_uu_u_ctrl_enablehost_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_enablehost_d
	localparam [0:0] sv2v_uu_u_ctrl_enablehost_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_enablehost(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_enablehost_we),
		.wd(ctrl_enablehost_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_enablehost_ext_d_0),
		.qe(),
		.q(reg2hw[324]),
		.qs(ctrl_enablehost_qs)
	);
	// Trace: design.sv:85924:3
	localparam signed [31:0] sv2v_uu_u_ctrl_enabletarget_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_enabletarget_d
	localparam [0:0] sv2v_uu_u_ctrl_enabletarget_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_enabletarget(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_enabletarget_we),
		.wd(ctrl_enabletarget_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_enabletarget_ext_d_0),
		.qe(),
		.q(reg2hw[323]),
		.qs(ctrl_enabletarget_qs)
	);
	// Trace: design.sv:85952:3
	localparam [31:0] sv2v_uu_u_status_fmtfull_DW = 1;
	// removed localparam type sv2v_uu_u_status_fmtfull_wd
	localparam [0:0] sv2v_uu_u_status_fmtfull_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_fmtfull(
		.re(status_fmtfull_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_fmtfull_ext_wd_0),
		.d(hw2reg[83]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_fmtfull_qs)
	);
	// Trace: design.sv:85967:3
	localparam [31:0] sv2v_uu_u_status_rxfull_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxfull_wd
	localparam [0:0] sv2v_uu_u_status_rxfull_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_rxfull(
		.re(status_rxfull_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxfull_ext_wd_0),
		.d(hw2reg[82]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_rxfull_qs)
	);
	// Trace: design.sv:85982:3
	localparam [31:0] sv2v_uu_u_status_fmtempty_DW = 1;
	// removed localparam type sv2v_uu_u_status_fmtempty_wd
	localparam [0:0] sv2v_uu_u_status_fmtempty_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_fmtempty(
		.re(status_fmtempty_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_fmtempty_ext_wd_0),
		.d(hw2reg[81]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_fmtempty_qs)
	);
	// Trace: design.sv:85997:3
	localparam [31:0] sv2v_uu_u_status_hostidle_DW = 1;
	// removed localparam type sv2v_uu_u_status_hostidle_wd
	localparam [0:0] sv2v_uu_u_status_hostidle_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_hostidle(
		.re(status_hostidle_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_hostidle_ext_wd_0),
		.d(hw2reg[80]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_hostidle_qs)
	);
	// Trace: design.sv:86012:3
	localparam [31:0] sv2v_uu_u_status_targetidle_DW = 1;
	// removed localparam type sv2v_uu_u_status_targetidle_wd
	localparam [0:0] sv2v_uu_u_status_targetidle_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_targetidle(
		.re(status_targetidle_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_targetidle_ext_wd_0),
		.d(hw2reg[79]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_targetidle_qs)
	);
	// Trace: design.sv:86027:3
	localparam [31:0] sv2v_uu_u_status_rxempty_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxempty_wd
	localparam [0:0] sv2v_uu_u_status_rxempty_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_rxempty(
		.re(status_rxempty_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxempty_ext_wd_0),
		.d(hw2reg[78]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_rxempty_qs)
	);
	// Trace: design.sv:86042:3
	localparam [31:0] sv2v_uu_u_status_txfull_DW = 1;
	// removed localparam type sv2v_uu_u_status_txfull_wd
	localparam [0:0] sv2v_uu_u_status_txfull_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_txfull(
		.re(status_txfull_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txfull_ext_wd_0),
		.d(hw2reg[77]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_txfull_qs)
	);
	// Trace: design.sv:86057:3
	localparam [31:0] sv2v_uu_u_status_acqfull_DW = 1;
	// removed localparam type sv2v_uu_u_status_acqfull_wd
	localparam [0:0] sv2v_uu_u_status_acqfull_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_acqfull(
		.re(status_acqfull_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_acqfull_ext_wd_0),
		.d(hw2reg[76]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_acqfull_qs)
	);
	// Trace: design.sv:86072:3
	localparam [31:0] sv2v_uu_u_status_txempty_DW = 1;
	// removed localparam type sv2v_uu_u_status_txempty_wd
	localparam [0:0] sv2v_uu_u_status_txempty_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_txempty(
		.re(status_txempty_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txempty_ext_wd_0),
		.d(hw2reg[75]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_txempty_qs)
	);
	// Trace: design.sv:86087:3
	localparam [31:0] sv2v_uu_u_status_acqempty_DW = 1;
	// removed localparam type sv2v_uu_u_status_acqempty_wd
	localparam [0:0] sv2v_uu_u_status_acqempty_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_acqempty(
		.re(status_acqempty_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_acqempty_ext_wd_0),
		.d(hw2reg[74]),
		.qre(),
		.qe(),
		.q(),
		.qs(status_acqempty_qs)
	);
	// Trace: design.sv:86103:3
	localparam [31:0] sv2v_uu_u_rdata_DW = 8;
	// removed localparam type sv2v_uu_u_rdata_wd
	localparam [7:0] sv2v_uu_u_rdata_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(8)) u_rdata(
		.re(rdata_re),
		.we(1'b0),
		.wd(sv2v_uu_u_rdata_ext_wd_0),
		.d(hw2reg[73-:8]),
		.qre(reg2hw[314]),
		.qe(),
		.q(reg2hw[322-:8]),
		.qs(rdata_qs)
	);
	// Trace: design.sv:86120:3
	localparam signed [31:0] sv2v_uu_u_fdata_fbyte_DW = 8;
	// removed localparam type sv2v_uu_u_fdata_fbyte_d
	localparam [7:0] sv2v_uu_u_fdata_fbyte_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("WO"),
		.RESVAL(8'h00)
	) u_fdata_fbyte(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fdata_fbyte_we),
		.wd(fdata_fbyte_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fdata_fbyte_ext_d_0),
		.qe(reg2hw[305]),
		.q(reg2hw[313-:8]),
		.qs()
	);
	// Trace: design.sv:86145:3
	localparam signed [31:0] sv2v_uu_u_fdata_start_DW = 1;
	// removed localparam type sv2v_uu_u_fdata_start_d
	localparam [0:0] sv2v_uu_u_fdata_start_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fdata_start(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fdata_start_we),
		.wd(fdata_start_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fdata_start_ext_d_0),
		.qe(reg2hw[303]),
		.q(reg2hw[304]),
		.qs()
	);
	// Trace: design.sv:86170:3
	localparam signed [31:0] sv2v_uu_u_fdata_stop_DW = 1;
	// removed localparam type sv2v_uu_u_fdata_stop_d
	localparam [0:0] sv2v_uu_u_fdata_stop_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fdata_stop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fdata_stop_we),
		.wd(fdata_stop_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fdata_stop_ext_d_0),
		.qe(reg2hw[301]),
		.q(reg2hw[302]),
		.qs()
	);
	// Trace: design.sv:86195:3
	localparam signed [31:0] sv2v_uu_u_fdata_read_DW = 1;
	// removed localparam type sv2v_uu_u_fdata_read_d
	localparam [0:0] sv2v_uu_u_fdata_read_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fdata_read(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fdata_read_we),
		.wd(fdata_read_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fdata_read_ext_d_0),
		.qe(reg2hw[299]),
		.q(reg2hw[300]),
		.qs()
	);
	// Trace: design.sv:86220:3
	localparam signed [31:0] sv2v_uu_u_fdata_rcont_DW = 1;
	// removed localparam type sv2v_uu_u_fdata_rcont_d
	localparam [0:0] sv2v_uu_u_fdata_rcont_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fdata_rcont(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fdata_rcont_we),
		.wd(fdata_rcont_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fdata_rcont_ext_d_0),
		.qe(reg2hw[297]),
		.q(reg2hw[298]),
		.qs()
	);
	// Trace: design.sv:86245:3
	localparam signed [31:0] sv2v_uu_u_fdata_nakok_DW = 1;
	// removed localparam type sv2v_uu_u_fdata_nakok_d
	localparam [0:0] sv2v_uu_u_fdata_nakok_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fdata_nakok(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fdata_nakok_we),
		.wd(fdata_nakok_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fdata_nakok_ext_d_0),
		.qe(reg2hw[295]),
		.q(reg2hw[296]),
		.qs()
	);
	// Trace: design.sv:86272:3
	localparam signed [31:0] sv2v_uu_u_fifo_ctrl_rxrst_DW = 1;
	// removed localparam type sv2v_uu_u_fifo_ctrl_rxrst_d
	localparam [0:0] sv2v_uu_u_fifo_ctrl_rxrst_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fifo_ctrl_rxrst(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_rxrst_we),
		.wd(fifo_ctrl_rxrst_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fifo_ctrl_rxrst_ext_d_0),
		.qe(reg2hw[293]),
		.q(reg2hw[294]),
		.qs()
	);
	// Trace: design.sv:86297:3
	localparam signed [31:0] sv2v_uu_u_fifo_ctrl_fmtrst_DW = 1;
	// removed localparam type sv2v_uu_u_fifo_ctrl_fmtrst_d
	localparam [0:0] sv2v_uu_u_fifo_ctrl_fmtrst_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fifo_ctrl_fmtrst(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_fmtrst_we),
		.wd(fifo_ctrl_fmtrst_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fifo_ctrl_fmtrst_ext_d_0),
		.qe(reg2hw[291]),
		.q(reg2hw[292]),
		.qs()
	);
	// Trace: design.sv:86322:3
	localparam signed [31:0] sv2v_uu_u_fifo_ctrl_rxilvl_DW = 3;
	// removed localparam type sv2v_uu_u_fifo_ctrl_rxilvl_d
	localparam [2:0] sv2v_uu_u_fifo_ctrl_rxilvl_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_fifo_ctrl_rxilvl(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_rxilvl_we),
		.wd(fifo_ctrl_rxilvl_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fifo_ctrl_rxilvl_ext_d_0),
		.qe(reg2hw[287]),
		.q(reg2hw[290-:3]),
		.qs(fifo_ctrl_rxilvl_qs)
	);
	// Trace: design.sv:86348:3
	localparam signed [31:0] sv2v_uu_u_fifo_ctrl_fmtilvl_DW = 2;
	// removed localparam type sv2v_uu_u_fifo_ctrl_fmtilvl_d
	localparam [1:0] sv2v_uu_u_fifo_ctrl_fmtilvl_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_fifo_ctrl_fmtilvl(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_fmtilvl_we),
		.wd(fifo_ctrl_fmtilvl_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fifo_ctrl_fmtilvl_ext_d_0),
		.qe(reg2hw[284]),
		.q(reg2hw[286-:2]),
		.qs(fifo_ctrl_fmtilvl_qs)
	);
	// Trace: design.sv:86374:3
	localparam signed [31:0] sv2v_uu_u_fifo_ctrl_acqrst_DW = 1;
	// removed localparam type sv2v_uu_u_fifo_ctrl_acqrst_d
	localparam [0:0] sv2v_uu_u_fifo_ctrl_acqrst_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fifo_ctrl_acqrst(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_acqrst_we),
		.wd(fifo_ctrl_acqrst_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fifo_ctrl_acqrst_ext_d_0),
		.qe(reg2hw[282]),
		.q(reg2hw[283]),
		.qs()
	);
	// Trace: design.sv:86399:3
	localparam signed [31:0] sv2v_uu_u_fifo_ctrl_txrst_DW = 1;
	// removed localparam type sv2v_uu_u_fifo_ctrl_txrst_d
	localparam [0:0] sv2v_uu_u_fifo_ctrl_txrst_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fifo_ctrl_txrst(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_txrst_we),
		.wd(fifo_ctrl_txrst_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fifo_ctrl_txrst_ext_d_0),
		.qe(reg2hw[280]),
		.q(reg2hw[281]),
		.qs()
	);
	// Trace: design.sv:86426:3
	localparam [31:0] sv2v_uu_u_fifo_status_fmtlvl_DW = 6;
	// removed localparam type sv2v_uu_u_fifo_status_fmtlvl_wd
	localparam [5:0] sv2v_uu_u_fifo_status_fmtlvl_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(6)) u_fifo_status_fmtlvl(
		.re(fifo_status_fmtlvl_re),
		.we(1'b0),
		.wd(sv2v_uu_u_fifo_status_fmtlvl_ext_wd_0),
		.d(hw2reg[65-:6]),
		.qre(),
		.qe(),
		.q(),
		.qs(fifo_status_fmtlvl_qs)
	);
	// Trace: design.sv:86441:3
	localparam [31:0] sv2v_uu_u_fifo_status_txlvl_DW = 6;
	// removed localparam type sv2v_uu_u_fifo_status_txlvl_wd
	localparam [5:0] sv2v_uu_u_fifo_status_txlvl_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(6)) u_fifo_status_txlvl(
		.re(fifo_status_txlvl_re),
		.we(1'b0),
		.wd(sv2v_uu_u_fifo_status_txlvl_ext_wd_0),
		.d(hw2reg[59-:6]),
		.qre(),
		.qe(),
		.q(),
		.qs(fifo_status_txlvl_qs)
	);
	// Trace: design.sv:86456:3
	localparam [31:0] sv2v_uu_u_fifo_status_rxlvl_DW = 6;
	// removed localparam type sv2v_uu_u_fifo_status_rxlvl_wd
	localparam [5:0] sv2v_uu_u_fifo_status_rxlvl_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(6)) u_fifo_status_rxlvl(
		.re(fifo_status_rxlvl_re),
		.we(1'b0),
		.wd(sv2v_uu_u_fifo_status_rxlvl_ext_wd_0),
		.d(hw2reg[53-:6]),
		.qre(),
		.qe(),
		.q(),
		.qs(fifo_status_rxlvl_qs)
	);
	// Trace: design.sv:86471:3
	localparam [31:0] sv2v_uu_u_fifo_status_acqlvl_DW = 6;
	// removed localparam type sv2v_uu_u_fifo_status_acqlvl_wd
	localparam [5:0] sv2v_uu_u_fifo_status_acqlvl_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(6)) u_fifo_status_acqlvl(
		.re(fifo_status_acqlvl_re),
		.we(1'b0),
		.wd(sv2v_uu_u_fifo_status_acqlvl_ext_wd_0),
		.d(hw2reg[47-:6]),
		.qre(),
		.qe(),
		.q(),
		.qs(fifo_status_acqlvl_qs)
	);
	// Trace: design.sv:86488:3
	localparam signed [31:0] sv2v_uu_u_ovrd_txovrden_DW = 1;
	// removed localparam type sv2v_uu_u_ovrd_txovrden_d
	localparam [0:0] sv2v_uu_u_ovrd_txovrden_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ovrd_txovrden(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ovrd_txovrden_we),
		.wd(ovrd_txovrden_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ovrd_txovrden_ext_d_0),
		.qe(),
		.q(reg2hw[279]),
		.qs(ovrd_txovrden_qs)
	);
	// Trace: design.sv:86514:3
	localparam signed [31:0] sv2v_uu_u_ovrd_sclval_DW = 1;
	// removed localparam type sv2v_uu_u_ovrd_sclval_d
	localparam [0:0] sv2v_uu_u_ovrd_sclval_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ovrd_sclval(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ovrd_sclval_we),
		.wd(ovrd_sclval_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ovrd_sclval_ext_d_0),
		.qe(),
		.q(reg2hw[278]),
		.qs(ovrd_sclval_qs)
	);
	// Trace: design.sv:86540:3
	localparam signed [31:0] sv2v_uu_u_ovrd_sdaval_DW = 1;
	// removed localparam type sv2v_uu_u_ovrd_sdaval_d
	localparam [0:0] sv2v_uu_u_ovrd_sdaval_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ovrd_sdaval(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ovrd_sdaval_we),
		.wd(ovrd_sdaval_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ovrd_sdaval_ext_d_0),
		.qe(),
		.q(reg2hw[277]),
		.qs(ovrd_sdaval_qs)
	);
	// Trace: design.sv:86568:3
	localparam [31:0] sv2v_uu_u_val_scl_rx_DW = 16;
	// removed localparam type sv2v_uu_u_val_scl_rx_wd
	localparam [15:0] sv2v_uu_u_val_scl_rx_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(16)) u_val_scl_rx(
		.re(val_scl_rx_re),
		.we(1'b0),
		.wd(sv2v_uu_u_val_scl_rx_ext_wd_0),
		.d(hw2reg[41-:16]),
		.qre(),
		.qe(),
		.q(),
		.qs(val_scl_rx_qs)
	);
	// Trace: design.sv:86583:3
	localparam [31:0] sv2v_uu_u_val_sda_rx_DW = 16;
	// removed localparam type sv2v_uu_u_val_sda_rx_wd
	localparam [15:0] sv2v_uu_u_val_sda_rx_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(16)) u_val_sda_rx(
		.re(val_sda_rx_re),
		.we(1'b0),
		.wd(sv2v_uu_u_val_sda_rx_ext_wd_0),
		.d(hw2reg[25-:16]),
		.qre(),
		.qe(),
		.q(),
		.qs(val_sda_rx_qs)
	);
	// Trace: design.sv:86600:3
	localparam signed [31:0] sv2v_uu_u_timing0_thigh_DW = 16;
	// removed localparam type sv2v_uu_u_timing0_thigh_d
	localparam [15:0] sv2v_uu_u_timing0_thigh_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing0_thigh(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing0_thigh_we),
		.wd(timing0_thigh_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing0_thigh_ext_d_0),
		.qe(),
		.q(reg2hw[276-:16]),
		.qs(timing0_thigh_qs)
	);
	// Trace: design.sv:86626:3
	localparam signed [31:0] sv2v_uu_u_timing0_tlow_DW = 16;
	// removed localparam type sv2v_uu_u_timing0_tlow_d
	localparam [15:0] sv2v_uu_u_timing0_tlow_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing0_tlow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing0_tlow_we),
		.wd(timing0_tlow_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing0_tlow_ext_d_0),
		.qe(),
		.q(reg2hw[260-:16]),
		.qs(timing0_tlow_qs)
	);
	// Trace: design.sv:86654:3
	localparam signed [31:0] sv2v_uu_u_timing1_t_r_DW = 16;
	// removed localparam type sv2v_uu_u_timing1_t_r_d
	localparam [15:0] sv2v_uu_u_timing1_t_r_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing1_t_r(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing1_t_r_we),
		.wd(timing1_t_r_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing1_t_r_ext_d_0),
		.qe(),
		.q(reg2hw[244-:16]),
		.qs(timing1_t_r_qs)
	);
	// Trace: design.sv:86680:3
	localparam signed [31:0] sv2v_uu_u_timing1_t_f_DW = 16;
	// removed localparam type sv2v_uu_u_timing1_t_f_d
	localparam [15:0] sv2v_uu_u_timing1_t_f_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing1_t_f(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing1_t_f_we),
		.wd(timing1_t_f_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing1_t_f_ext_d_0),
		.qe(),
		.q(reg2hw[228-:16]),
		.qs(timing1_t_f_qs)
	);
	// Trace: design.sv:86708:3
	localparam signed [31:0] sv2v_uu_u_timing2_tsu_sta_DW = 16;
	// removed localparam type sv2v_uu_u_timing2_tsu_sta_d
	localparam [15:0] sv2v_uu_u_timing2_tsu_sta_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing2_tsu_sta(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing2_tsu_sta_we),
		.wd(timing2_tsu_sta_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing2_tsu_sta_ext_d_0),
		.qe(),
		.q(reg2hw[212-:16]),
		.qs(timing2_tsu_sta_qs)
	);
	// Trace: design.sv:86734:3
	localparam signed [31:0] sv2v_uu_u_timing2_thd_sta_DW = 16;
	// removed localparam type sv2v_uu_u_timing2_thd_sta_d
	localparam [15:0] sv2v_uu_u_timing2_thd_sta_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing2_thd_sta(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing2_thd_sta_we),
		.wd(timing2_thd_sta_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing2_thd_sta_ext_d_0),
		.qe(),
		.q(reg2hw[196-:16]),
		.qs(timing2_thd_sta_qs)
	);
	// Trace: design.sv:86762:3
	localparam signed [31:0] sv2v_uu_u_timing3_tsu_dat_DW = 16;
	// removed localparam type sv2v_uu_u_timing3_tsu_dat_d
	localparam [15:0] sv2v_uu_u_timing3_tsu_dat_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing3_tsu_dat(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing3_tsu_dat_we),
		.wd(timing3_tsu_dat_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing3_tsu_dat_ext_d_0),
		.qe(),
		.q(reg2hw[180-:16]),
		.qs(timing3_tsu_dat_qs)
	);
	// Trace: design.sv:86788:3
	localparam signed [31:0] sv2v_uu_u_timing3_thd_dat_DW = 16;
	// removed localparam type sv2v_uu_u_timing3_thd_dat_d
	localparam [15:0] sv2v_uu_u_timing3_thd_dat_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing3_thd_dat(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing3_thd_dat_we),
		.wd(timing3_thd_dat_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing3_thd_dat_ext_d_0),
		.qe(),
		.q(reg2hw[164-:16]),
		.qs(timing3_thd_dat_qs)
	);
	// Trace: design.sv:86816:3
	localparam signed [31:0] sv2v_uu_u_timing4_tsu_sto_DW = 16;
	// removed localparam type sv2v_uu_u_timing4_tsu_sto_d
	localparam [15:0] sv2v_uu_u_timing4_tsu_sto_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing4_tsu_sto(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing4_tsu_sto_we),
		.wd(timing4_tsu_sto_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing4_tsu_sto_ext_d_0),
		.qe(),
		.q(reg2hw[148-:16]),
		.qs(timing4_tsu_sto_qs)
	);
	// Trace: design.sv:86842:3
	localparam signed [31:0] sv2v_uu_u_timing4_t_buf_DW = 16;
	// removed localparam type sv2v_uu_u_timing4_t_buf_d
	localparam [15:0] sv2v_uu_u_timing4_t_buf_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_timing4_t_buf(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timing4_t_buf_we),
		.wd(timing4_t_buf_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timing4_t_buf_ext_d_0),
		.qe(),
		.q(reg2hw[132-:16]),
		.qs(timing4_t_buf_qs)
	);
	// Trace: design.sv:86870:3
	localparam signed [31:0] sv2v_uu_u_timeout_ctrl_val_DW = 31;
	// removed localparam type sv2v_uu_u_timeout_ctrl_val_d
	localparam [30:0] sv2v_uu_u_timeout_ctrl_val_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(31),
		.SWACCESS("RW"),
		.RESVAL(31'h00000000)
	) u_timeout_ctrl_val(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timeout_ctrl_val_we),
		.wd(timeout_ctrl_val_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timeout_ctrl_val_ext_d_0),
		.qe(),
		.q(reg2hw[116-:31]),
		.qs(timeout_ctrl_val_qs)
	);
	// Trace: design.sv:86896:3
	localparam signed [31:0] sv2v_uu_u_timeout_ctrl_en_DW = 1;
	// removed localparam type sv2v_uu_u_timeout_ctrl_en_d
	localparam [0:0] sv2v_uu_u_timeout_ctrl_en_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_timeout_ctrl_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timeout_ctrl_en_we),
		.wd(timeout_ctrl_en_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timeout_ctrl_en_ext_d_0),
		.qe(),
		.q(reg2hw[85]),
		.qs(timeout_ctrl_en_qs)
	);
	// Trace: design.sv:86924:3
	localparam signed [31:0] sv2v_uu_u_target_id_address0_DW = 7;
	// removed localparam type sv2v_uu_u_target_id_address0_d
	localparam [6:0] sv2v_uu_u_target_id_address0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(7),
		.SWACCESS("RW"),
		.RESVAL(7'h00)
	) u_target_id_address0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(target_id_address0_we),
		.wd(target_id_address0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_target_id_address0_ext_d_0),
		.qe(),
		.q(reg2hw[84-:7]),
		.qs(target_id_address0_qs)
	);
	// Trace: design.sv:86950:3
	localparam signed [31:0] sv2v_uu_u_target_id_mask0_DW = 7;
	// removed localparam type sv2v_uu_u_target_id_mask0_d
	localparam [6:0] sv2v_uu_u_target_id_mask0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(7),
		.SWACCESS("RW"),
		.RESVAL(7'h00)
	) u_target_id_mask0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(target_id_mask0_we),
		.wd(target_id_mask0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_target_id_mask0_ext_d_0),
		.qe(),
		.q(reg2hw[77-:7]),
		.qs(target_id_mask0_qs)
	);
	// Trace: design.sv:86976:3
	localparam signed [31:0] sv2v_uu_u_target_id_address1_DW = 7;
	// removed localparam type sv2v_uu_u_target_id_address1_d
	localparam [6:0] sv2v_uu_u_target_id_address1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(7),
		.SWACCESS("RW"),
		.RESVAL(7'h00)
	) u_target_id_address1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(target_id_address1_we),
		.wd(target_id_address1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_target_id_address1_ext_d_0),
		.qe(),
		.q(reg2hw[70-:7]),
		.qs(target_id_address1_qs)
	);
	// Trace: design.sv:87002:3
	localparam signed [31:0] sv2v_uu_u_target_id_mask1_DW = 7;
	// removed localparam type sv2v_uu_u_target_id_mask1_d
	localparam [6:0] sv2v_uu_u_target_id_mask1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(7),
		.SWACCESS("RW"),
		.RESVAL(7'h00)
	) u_target_id_mask1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(target_id_mask1_we),
		.wd(target_id_mask1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_target_id_mask1_ext_d_0),
		.qe(),
		.q(reg2hw[63-:7]),
		.qs(target_id_mask1_qs)
	);
	// Trace: design.sv:87030:3
	localparam [31:0] sv2v_uu_u_acqdata_abyte_DW = 8;
	// removed localparam type sv2v_uu_u_acqdata_abyte_wd
	localparam [7:0] sv2v_uu_u_acqdata_abyte_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(8)) u_acqdata_abyte(
		.re(acqdata_abyte_re),
		.we(1'b0),
		.wd(sv2v_uu_u_acqdata_abyte_ext_wd_0),
		.d(hw2reg[9-:8]),
		.qre(reg2hw[48]),
		.qe(),
		.q(reg2hw[56-:8]),
		.qs(acqdata_abyte_qs)
	);
	// Trace: design.sv:87045:3
	localparam [31:0] sv2v_uu_u_acqdata_signal_DW = 2;
	// removed localparam type sv2v_uu_u_acqdata_signal_wd
	localparam [1:0] sv2v_uu_u_acqdata_signal_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(2)) u_acqdata_signal(
		.re(acqdata_signal_re),
		.we(1'b0),
		.wd(sv2v_uu_u_acqdata_signal_ext_wd_0),
		.d(hw2reg[1-:2]),
		.qre(reg2hw[45]),
		.qe(),
		.q(reg2hw[47-:2]),
		.qs(acqdata_signal_qs)
	);
	// Trace: design.sv:87061:3
	localparam signed [31:0] sv2v_uu_u_txdata_DW = 8;
	// removed localparam type sv2v_uu_u_txdata_d
	localparam [7:0] sv2v_uu_u_txdata_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("WO"),
		.RESVAL(8'h00)
	) u_txdata(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(txdata_we),
		.wd(txdata_wd),
		.de(1'b0),
		.d(sv2v_uu_u_txdata_ext_d_0),
		.qe(reg2hw[36]),
		.q(reg2hw[44-:8]),
		.qs()
	);
	// Trace: design.sv:87088:3
	localparam signed [31:0] sv2v_uu_u_stretch_ctrl_enableaddr_DW = 1;
	// removed localparam type sv2v_uu_u_stretch_ctrl_enableaddr_d
	localparam [0:0] sv2v_uu_u_stretch_ctrl_enableaddr_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_stretch_ctrl_enableaddr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(stretch_ctrl_enableaddr_we),
		.wd(stretch_ctrl_enableaddr_wd),
		.de(1'b0),
		.d(sv2v_uu_u_stretch_ctrl_enableaddr_ext_d_0),
		.qe(),
		.q(reg2hw[35]),
		.qs(stretch_ctrl_enableaddr_qs)
	);
	// Trace: design.sv:87114:3
	localparam signed [31:0] sv2v_uu_u_stretch_ctrl_enabletx_DW = 1;
	// removed localparam type sv2v_uu_u_stretch_ctrl_enabletx_d
	localparam [0:0] sv2v_uu_u_stretch_ctrl_enabletx_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_stretch_ctrl_enabletx(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(stretch_ctrl_enabletx_we),
		.wd(stretch_ctrl_enabletx_wd),
		.de(1'b0),
		.d(sv2v_uu_u_stretch_ctrl_enabletx_ext_d_0),
		.qe(),
		.q(reg2hw[34]),
		.qs(stretch_ctrl_enabletx_qs)
	);
	// Trace: design.sv:87140:3
	localparam signed [31:0] sv2v_uu_u_stretch_ctrl_enableacq_DW = 1;
	// removed localparam type sv2v_uu_u_stretch_ctrl_enableacq_d
	localparam [0:0] sv2v_uu_u_stretch_ctrl_enableacq_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_stretch_ctrl_enableacq(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(stretch_ctrl_enableacq_we),
		.wd(stretch_ctrl_enableacq_wd),
		.de(1'b0),
		.d(sv2v_uu_u_stretch_ctrl_enableacq_ext_d_0),
		.qe(),
		.q(reg2hw[33]),
		.qs(stretch_ctrl_enableacq_qs)
	);
	// Trace: design.sv:87166:3
	localparam signed [31:0] sv2v_uu_u_stretch_ctrl_stop_DW = 1;
	// removed localparam type sv2v_uu_u_stretch_ctrl_stop_d
	localparam [0:0] sv2v_uu_u_stretch_ctrl_stop_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_stretch_ctrl_stop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(stretch_ctrl_stop_we),
		.wd(stretch_ctrl_stop_wd),
		.de(1'b0),
		.d(sv2v_uu_u_stretch_ctrl_stop_ext_d_0),
		.qe(),
		.q(reg2hw[32]),
		.qs(stretch_ctrl_stop_qs)
	);
	// Trace: design.sv:87193:3
	localparam signed [31:0] sv2v_uu_u_host_timeout_ctrl_DW = 32;
	// removed localparam type sv2v_uu_u_host_timeout_ctrl_d
	localparam [31:0] sv2v_uu_u_host_timeout_ctrl_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_host_timeout_ctrl(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(host_timeout_ctrl_we),
		.wd(host_timeout_ctrl_wd),
		.de(1'b0),
		.d(sv2v_uu_u_host_timeout_ctrl_ext_d_0),
		.qe(),
		.q(reg2hw[31-:32]),
		.qs(host_timeout_ctrl_qs)
	);
	// Trace: design.sv:87220:3
	reg [21:0] addr_hit;
	// Trace: design.sv:87221:3
	localparam signed [31:0] i2c_reg_pkg_BlockAw = 7;
	localparam [6:0] i2c_reg_pkg_I2C_ACQDATA_OFFSET = 7'h48;
	localparam [6:0] i2c_reg_pkg_I2C_CTRL_OFFSET = 7'h0c;
	localparam [6:0] i2c_reg_pkg_I2C_FDATA_OFFSET = 7'h18;
	localparam [6:0] i2c_reg_pkg_I2C_FIFO_CTRL_OFFSET = 7'h1c;
	localparam [6:0] i2c_reg_pkg_I2C_FIFO_STATUS_OFFSET = 7'h20;
	localparam [6:0] i2c_reg_pkg_I2C_HOST_TIMEOUT_CTRL_OFFSET = 7'h54;
	localparam [6:0] i2c_reg_pkg_I2C_INTR_ENABLE_OFFSET = 7'h04;
	localparam [6:0] i2c_reg_pkg_I2C_INTR_STATE_OFFSET = 7'h00;
	localparam [6:0] i2c_reg_pkg_I2C_INTR_TEST_OFFSET = 7'h08;
	localparam [6:0] i2c_reg_pkg_I2C_OVRD_OFFSET = 7'h24;
	localparam [6:0] i2c_reg_pkg_I2C_RDATA_OFFSET = 7'h14;
	localparam [6:0] i2c_reg_pkg_I2C_STATUS_OFFSET = 7'h10;
	localparam [6:0] i2c_reg_pkg_I2C_STRETCH_CTRL_OFFSET = 7'h50;
	localparam [6:0] i2c_reg_pkg_I2C_TARGET_ID_OFFSET = 7'h44;
	localparam [6:0] i2c_reg_pkg_I2C_TIMEOUT_CTRL_OFFSET = 7'h40;
	localparam [6:0] i2c_reg_pkg_I2C_TIMING0_OFFSET = 7'h2c;
	localparam [6:0] i2c_reg_pkg_I2C_TIMING1_OFFSET = 7'h30;
	localparam [6:0] i2c_reg_pkg_I2C_TIMING2_OFFSET = 7'h34;
	localparam [6:0] i2c_reg_pkg_I2C_TIMING3_OFFSET = 7'h38;
	localparam [6:0] i2c_reg_pkg_I2C_TIMING4_OFFSET = 7'h3c;
	localparam [6:0] i2c_reg_pkg_I2C_TXDATA_OFFSET = 7'h4c;
	localparam [6:0] i2c_reg_pkg_I2C_VAL_OFFSET = 7'h28;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:87222:5
		addr_hit = 1'sb0;
		// Trace: design.sv:87223:5
		addr_hit[0] = reg_addr == i2c_reg_pkg_I2C_INTR_STATE_OFFSET;
		// Trace: design.sv:87224:5
		addr_hit[1] = reg_addr == i2c_reg_pkg_I2C_INTR_ENABLE_OFFSET;
		// Trace: design.sv:87225:5
		addr_hit[2] = reg_addr == i2c_reg_pkg_I2C_INTR_TEST_OFFSET;
		// Trace: design.sv:87226:5
		addr_hit[3] = reg_addr == i2c_reg_pkg_I2C_CTRL_OFFSET;
		// Trace: design.sv:87227:5
		addr_hit[4] = reg_addr == i2c_reg_pkg_I2C_STATUS_OFFSET;
		// Trace: design.sv:87228:5
		addr_hit[5] = reg_addr == i2c_reg_pkg_I2C_RDATA_OFFSET;
		// Trace: design.sv:87229:5
		addr_hit[6] = reg_addr == i2c_reg_pkg_I2C_FDATA_OFFSET;
		// Trace: design.sv:87230:5
		addr_hit[7] = reg_addr == i2c_reg_pkg_I2C_FIFO_CTRL_OFFSET;
		// Trace: design.sv:87231:5
		addr_hit[8] = reg_addr == i2c_reg_pkg_I2C_FIFO_STATUS_OFFSET;
		// Trace: design.sv:87232:5
		addr_hit[9] = reg_addr == i2c_reg_pkg_I2C_OVRD_OFFSET;
		// Trace: design.sv:87233:5
		addr_hit[10] = reg_addr == i2c_reg_pkg_I2C_VAL_OFFSET;
		// Trace: design.sv:87234:5
		addr_hit[11] = reg_addr == i2c_reg_pkg_I2C_TIMING0_OFFSET;
		// Trace: design.sv:87235:5
		addr_hit[12] = reg_addr == i2c_reg_pkg_I2C_TIMING1_OFFSET;
		// Trace: design.sv:87236:5
		addr_hit[13] = reg_addr == i2c_reg_pkg_I2C_TIMING2_OFFSET;
		// Trace: design.sv:87237:5
		addr_hit[14] = reg_addr == i2c_reg_pkg_I2C_TIMING3_OFFSET;
		// Trace: design.sv:87238:5
		addr_hit[15] = reg_addr == i2c_reg_pkg_I2C_TIMING4_OFFSET;
		// Trace: design.sv:87239:5
		addr_hit[16] = reg_addr == i2c_reg_pkg_I2C_TIMEOUT_CTRL_OFFSET;
		// Trace: design.sv:87240:5
		addr_hit[17] = reg_addr == i2c_reg_pkg_I2C_TARGET_ID_OFFSET;
		// Trace: design.sv:87241:5
		addr_hit[18] = reg_addr == i2c_reg_pkg_I2C_ACQDATA_OFFSET;
		// Trace: design.sv:87242:5
		addr_hit[19] = reg_addr == i2c_reg_pkg_I2C_TXDATA_OFFSET;
		// Trace: design.sv:87243:5
		addr_hit[20] = reg_addr == i2c_reg_pkg_I2C_STRETCH_CTRL_OFFSET;
		// Trace: design.sv:87244:5
		addr_hit[21] = reg_addr == i2c_reg_pkg_I2C_HOST_TIMEOUT_CTRL_OFFSET;
	end
	// Trace: design.sv:87247:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:87250:3
	localparam [87:0] i2c_reg_pkg_I2C_PERMIT = 88'b0011001100110001001100010011001111110001111111111111111111111111111111110011000100011111;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:87251:5
		wr_err = reg_we & ((((((((((((((((((((((addr_hit[0] & |(i2c_reg_pkg_I2C_PERMIT[84+:4] & ~reg_be)) | (addr_hit[1] & |(i2c_reg_pkg_I2C_PERMIT[80+:4] & ~reg_be))) | (addr_hit[2] & |(i2c_reg_pkg_I2C_PERMIT[76+:4] & ~reg_be))) | (addr_hit[3] & |(i2c_reg_pkg_I2C_PERMIT[72+:4] & ~reg_be))) | (addr_hit[4] & |(i2c_reg_pkg_I2C_PERMIT[68+:4] & ~reg_be))) | (addr_hit[5] & |(i2c_reg_pkg_I2C_PERMIT[64+:4] & ~reg_be))) | (addr_hit[6] & |(i2c_reg_pkg_I2C_PERMIT[60+:4] & ~reg_be))) | (addr_hit[7] & |(i2c_reg_pkg_I2C_PERMIT[56+:4] & ~reg_be))) | (addr_hit[8] & |(i2c_reg_pkg_I2C_PERMIT[52+:4] & ~reg_be))) | (addr_hit[9] & |(i2c_reg_pkg_I2C_PERMIT[48+:4] & ~reg_be))) | (addr_hit[10] & |(i2c_reg_pkg_I2C_PERMIT[44+:4] & ~reg_be))) | (addr_hit[11] & |(i2c_reg_pkg_I2C_PERMIT[40+:4] & ~reg_be))) | (addr_hit[12] & |(i2c_reg_pkg_I2C_PERMIT[36+:4] & ~reg_be))) | (addr_hit[13] & |(i2c_reg_pkg_I2C_PERMIT[32+:4] & ~reg_be))) | (addr_hit[14] & |(i2c_reg_pkg_I2C_PERMIT[28+:4] & ~reg_be))) | (addr_hit[15] & |(i2c_reg_pkg_I2C_PERMIT[24+:4] & ~reg_be))) | (addr_hit[16] & |(i2c_reg_pkg_I2C_PERMIT[20+:4] & ~reg_be))) | (addr_hit[17] & |(i2c_reg_pkg_I2C_PERMIT[16+:4] & ~reg_be))) | (addr_hit[18] & |(i2c_reg_pkg_I2C_PERMIT[12+:4] & ~reg_be))) | (addr_hit[19] & |(i2c_reg_pkg_I2C_PERMIT[8+:4] & ~reg_be))) | (addr_hit[20] & |(i2c_reg_pkg_I2C_PERMIT[4+:4] & ~reg_be))) | (addr_hit[21] & |(i2c_reg_pkg_I2C_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:87276:3
	assign intr_state_fmt_watermark_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87277:3
	assign intr_state_fmt_watermark_wd = reg_wdata[0];
	// Trace: design.sv:87279:3
	assign intr_state_rx_watermark_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87280:3
	assign intr_state_rx_watermark_wd = reg_wdata[1];
	// Trace: design.sv:87282:3
	assign intr_state_fmt_overflow_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87283:3
	assign intr_state_fmt_overflow_wd = reg_wdata[2];
	// Trace: design.sv:87285:3
	assign intr_state_rx_overflow_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87286:3
	assign intr_state_rx_overflow_wd = reg_wdata[3];
	// Trace: design.sv:87288:3
	assign intr_state_nak_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87289:3
	assign intr_state_nak_wd = reg_wdata[4];
	// Trace: design.sv:87291:3
	assign intr_state_scl_interference_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87292:3
	assign intr_state_scl_interference_wd = reg_wdata[5];
	// Trace: design.sv:87294:3
	assign intr_state_sda_interference_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87295:3
	assign intr_state_sda_interference_wd = reg_wdata[6];
	// Trace: design.sv:87297:3
	assign intr_state_stretch_timeout_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87298:3
	assign intr_state_stretch_timeout_wd = reg_wdata[7];
	// Trace: design.sv:87300:3
	assign intr_state_sda_unstable_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87301:3
	assign intr_state_sda_unstable_wd = reg_wdata[8];
	// Trace: design.sv:87303:3
	assign intr_state_trans_complete_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87304:3
	assign intr_state_trans_complete_wd = reg_wdata[9];
	// Trace: design.sv:87306:3
	assign intr_state_tx_empty_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87307:3
	assign intr_state_tx_empty_wd = reg_wdata[10];
	// Trace: design.sv:87309:3
	assign intr_state_tx_nonempty_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87310:3
	assign intr_state_tx_nonempty_wd = reg_wdata[11];
	// Trace: design.sv:87312:3
	assign intr_state_tx_overflow_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87313:3
	assign intr_state_tx_overflow_wd = reg_wdata[12];
	// Trace: design.sv:87315:3
	assign intr_state_acq_overflow_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87316:3
	assign intr_state_acq_overflow_wd = reg_wdata[13];
	// Trace: design.sv:87318:3
	assign intr_state_ack_stop_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87319:3
	assign intr_state_ack_stop_wd = reg_wdata[14];
	// Trace: design.sv:87321:3
	assign intr_state_host_timeout_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:87322:3
	assign intr_state_host_timeout_wd = reg_wdata[15];
	// Trace: design.sv:87324:3
	assign intr_enable_fmt_watermark_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87325:3
	assign intr_enable_fmt_watermark_wd = reg_wdata[0];
	// Trace: design.sv:87327:3
	assign intr_enable_rx_watermark_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87328:3
	assign intr_enable_rx_watermark_wd = reg_wdata[1];
	// Trace: design.sv:87330:3
	assign intr_enable_fmt_overflow_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87331:3
	assign intr_enable_fmt_overflow_wd = reg_wdata[2];
	// Trace: design.sv:87333:3
	assign intr_enable_rx_overflow_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87334:3
	assign intr_enable_rx_overflow_wd = reg_wdata[3];
	// Trace: design.sv:87336:3
	assign intr_enable_nak_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87337:3
	assign intr_enable_nak_wd = reg_wdata[4];
	// Trace: design.sv:87339:3
	assign intr_enable_scl_interference_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87340:3
	assign intr_enable_scl_interference_wd = reg_wdata[5];
	// Trace: design.sv:87342:3
	assign intr_enable_sda_interference_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87343:3
	assign intr_enable_sda_interference_wd = reg_wdata[6];
	// Trace: design.sv:87345:3
	assign intr_enable_stretch_timeout_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87346:3
	assign intr_enable_stretch_timeout_wd = reg_wdata[7];
	// Trace: design.sv:87348:3
	assign intr_enable_sda_unstable_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87349:3
	assign intr_enable_sda_unstable_wd = reg_wdata[8];
	// Trace: design.sv:87351:3
	assign intr_enable_trans_complete_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87352:3
	assign intr_enable_trans_complete_wd = reg_wdata[9];
	// Trace: design.sv:87354:3
	assign intr_enable_tx_empty_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87355:3
	assign intr_enable_tx_empty_wd = reg_wdata[10];
	// Trace: design.sv:87357:3
	assign intr_enable_tx_nonempty_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87358:3
	assign intr_enable_tx_nonempty_wd = reg_wdata[11];
	// Trace: design.sv:87360:3
	assign intr_enable_tx_overflow_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87361:3
	assign intr_enable_tx_overflow_wd = reg_wdata[12];
	// Trace: design.sv:87363:3
	assign intr_enable_acq_overflow_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87364:3
	assign intr_enable_acq_overflow_wd = reg_wdata[13];
	// Trace: design.sv:87366:3
	assign intr_enable_ack_stop_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87367:3
	assign intr_enable_ack_stop_wd = reg_wdata[14];
	// Trace: design.sv:87369:3
	assign intr_enable_host_timeout_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:87370:3
	assign intr_enable_host_timeout_wd = reg_wdata[15];
	// Trace: design.sv:87372:3
	assign intr_test_fmt_watermark_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87373:3
	assign intr_test_fmt_watermark_wd = reg_wdata[0];
	// Trace: design.sv:87375:3
	assign intr_test_rx_watermark_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87376:3
	assign intr_test_rx_watermark_wd = reg_wdata[1];
	// Trace: design.sv:87378:3
	assign intr_test_fmt_overflow_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87379:3
	assign intr_test_fmt_overflow_wd = reg_wdata[2];
	// Trace: design.sv:87381:3
	assign intr_test_rx_overflow_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87382:3
	assign intr_test_rx_overflow_wd = reg_wdata[3];
	// Trace: design.sv:87384:3
	assign intr_test_nak_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87385:3
	assign intr_test_nak_wd = reg_wdata[4];
	// Trace: design.sv:87387:3
	assign intr_test_scl_interference_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87388:3
	assign intr_test_scl_interference_wd = reg_wdata[5];
	// Trace: design.sv:87390:3
	assign intr_test_sda_interference_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87391:3
	assign intr_test_sda_interference_wd = reg_wdata[6];
	// Trace: design.sv:87393:3
	assign intr_test_stretch_timeout_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87394:3
	assign intr_test_stretch_timeout_wd = reg_wdata[7];
	// Trace: design.sv:87396:3
	assign intr_test_sda_unstable_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87397:3
	assign intr_test_sda_unstable_wd = reg_wdata[8];
	// Trace: design.sv:87399:3
	assign intr_test_trans_complete_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87400:3
	assign intr_test_trans_complete_wd = reg_wdata[9];
	// Trace: design.sv:87402:3
	assign intr_test_tx_empty_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87403:3
	assign intr_test_tx_empty_wd = reg_wdata[10];
	// Trace: design.sv:87405:3
	assign intr_test_tx_nonempty_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87406:3
	assign intr_test_tx_nonempty_wd = reg_wdata[11];
	// Trace: design.sv:87408:3
	assign intr_test_tx_overflow_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87409:3
	assign intr_test_tx_overflow_wd = reg_wdata[12];
	// Trace: design.sv:87411:3
	assign intr_test_acq_overflow_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87412:3
	assign intr_test_acq_overflow_wd = reg_wdata[13];
	// Trace: design.sv:87414:3
	assign intr_test_ack_stop_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87415:3
	assign intr_test_ack_stop_wd = reg_wdata[14];
	// Trace: design.sv:87417:3
	assign intr_test_host_timeout_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:87418:3
	assign intr_test_host_timeout_wd = reg_wdata[15];
	// Trace: design.sv:87420:3
	assign ctrl_enablehost_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:87421:3
	assign ctrl_enablehost_wd = reg_wdata[0];
	// Trace: design.sv:87423:3
	assign ctrl_enabletarget_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:87424:3
	assign ctrl_enabletarget_wd = reg_wdata[1];
	// Trace: design.sv:87426:3
	assign status_fmtfull_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87428:3
	assign status_rxfull_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87430:3
	assign status_fmtempty_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87432:3
	assign status_hostidle_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87434:3
	assign status_targetidle_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87436:3
	assign status_rxempty_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87438:3
	assign status_txfull_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87440:3
	assign status_acqfull_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87442:3
	assign status_txempty_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87444:3
	assign status_acqempty_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:87446:3
	assign rdata_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:87448:3
	assign fdata_fbyte_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:87449:3
	assign fdata_fbyte_wd = reg_wdata[7:0];
	// Trace: design.sv:87451:3
	assign fdata_start_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:87452:3
	assign fdata_start_wd = reg_wdata[8];
	// Trace: design.sv:87454:3
	assign fdata_stop_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:87455:3
	assign fdata_stop_wd = reg_wdata[9];
	// Trace: design.sv:87457:3
	assign fdata_read_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:87458:3
	assign fdata_read_wd = reg_wdata[10];
	// Trace: design.sv:87460:3
	assign fdata_rcont_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:87461:3
	assign fdata_rcont_wd = reg_wdata[11];
	// Trace: design.sv:87463:3
	assign fdata_nakok_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:87464:3
	assign fdata_nakok_wd = reg_wdata[12];
	// Trace: design.sv:87466:3
	assign fifo_ctrl_rxrst_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:87467:3
	assign fifo_ctrl_rxrst_wd = reg_wdata[0];
	// Trace: design.sv:87469:3
	assign fifo_ctrl_fmtrst_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:87470:3
	assign fifo_ctrl_fmtrst_wd = reg_wdata[1];
	// Trace: design.sv:87472:3
	assign fifo_ctrl_rxilvl_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:87473:3
	assign fifo_ctrl_rxilvl_wd = reg_wdata[4:2];
	// Trace: design.sv:87475:3
	assign fifo_ctrl_fmtilvl_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:87476:3
	assign fifo_ctrl_fmtilvl_wd = reg_wdata[6:5];
	// Trace: design.sv:87478:3
	assign fifo_ctrl_acqrst_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:87479:3
	assign fifo_ctrl_acqrst_wd = reg_wdata[7];
	// Trace: design.sv:87481:3
	assign fifo_ctrl_txrst_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:87482:3
	assign fifo_ctrl_txrst_wd = reg_wdata[8];
	// Trace: design.sv:87484:3
	assign fifo_status_fmtlvl_re = (addr_hit[8] & reg_re) & !reg_error;
	// Trace: design.sv:87486:3
	assign fifo_status_txlvl_re = (addr_hit[8] & reg_re) & !reg_error;
	// Trace: design.sv:87488:3
	assign fifo_status_rxlvl_re = (addr_hit[8] & reg_re) & !reg_error;
	// Trace: design.sv:87490:3
	assign fifo_status_acqlvl_re = (addr_hit[8] & reg_re) & !reg_error;
	// Trace: design.sv:87492:3
	assign ovrd_txovrden_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:87493:3
	assign ovrd_txovrden_wd = reg_wdata[0];
	// Trace: design.sv:87495:3
	assign ovrd_sclval_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:87496:3
	assign ovrd_sclval_wd = reg_wdata[1];
	// Trace: design.sv:87498:3
	assign ovrd_sdaval_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:87499:3
	assign ovrd_sdaval_wd = reg_wdata[2];
	// Trace: design.sv:87501:3
	assign val_scl_rx_re = (addr_hit[10] & reg_re) & !reg_error;
	// Trace: design.sv:87503:3
	assign val_sda_rx_re = (addr_hit[10] & reg_re) & !reg_error;
	// Trace: design.sv:87505:3
	assign timing0_thigh_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:87506:3
	assign timing0_thigh_wd = reg_wdata[15:0];
	// Trace: design.sv:87508:3
	assign timing0_tlow_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:87509:3
	assign timing0_tlow_wd = reg_wdata[31:16];
	// Trace: design.sv:87511:3
	assign timing1_t_r_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:87512:3
	assign timing1_t_r_wd = reg_wdata[15:0];
	// Trace: design.sv:87514:3
	assign timing1_t_f_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:87515:3
	assign timing1_t_f_wd = reg_wdata[31:16];
	// Trace: design.sv:87517:3
	assign timing2_tsu_sta_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:87518:3
	assign timing2_tsu_sta_wd = reg_wdata[15:0];
	// Trace: design.sv:87520:3
	assign timing2_thd_sta_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:87521:3
	assign timing2_thd_sta_wd = reg_wdata[31:16];
	// Trace: design.sv:87523:3
	assign timing3_tsu_dat_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:87524:3
	assign timing3_tsu_dat_wd = reg_wdata[15:0];
	// Trace: design.sv:87526:3
	assign timing3_thd_dat_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:87527:3
	assign timing3_thd_dat_wd = reg_wdata[31:16];
	// Trace: design.sv:87529:3
	assign timing4_tsu_sto_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:87530:3
	assign timing4_tsu_sto_wd = reg_wdata[15:0];
	// Trace: design.sv:87532:3
	assign timing4_t_buf_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:87533:3
	assign timing4_t_buf_wd = reg_wdata[31:16];
	// Trace: design.sv:87535:3
	assign timeout_ctrl_val_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:87536:3
	assign timeout_ctrl_val_wd = reg_wdata[30:0];
	// Trace: design.sv:87538:3
	assign timeout_ctrl_en_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:87539:3
	assign timeout_ctrl_en_wd = reg_wdata[31];
	// Trace: design.sv:87541:3
	assign target_id_address0_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:87542:3
	assign target_id_address0_wd = reg_wdata[6:0];
	// Trace: design.sv:87544:3
	assign target_id_mask0_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:87545:3
	assign target_id_mask0_wd = reg_wdata[13:7];
	// Trace: design.sv:87547:3
	assign target_id_address1_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:87548:3
	assign target_id_address1_wd = reg_wdata[20:14];
	// Trace: design.sv:87550:3
	assign target_id_mask1_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:87551:3
	assign target_id_mask1_wd = reg_wdata[27:21];
	// Trace: design.sv:87553:3
	assign acqdata_abyte_re = (addr_hit[18] & reg_re) & !reg_error;
	// Trace: design.sv:87555:3
	assign acqdata_signal_re = (addr_hit[18] & reg_re) & !reg_error;
	// Trace: design.sv:87557:3
	assign txdata_we = (addr_hit[19] & reg_we) & !reg_error;
	// Trace: design.sv:87558:3
	assign txdata_wd = reg_wdata[7:0];
	// Trace: design.sv:87560:3
	assign stretch_ctrl_enableaddr_we = (addr_hit[20] & reg_we) & !reg_error;
	// Trace: design.sv:87561:3
	assign stretch_ctrl_enableaddr_wd = reg_wdata[0];
	// Trace: design.sv:87563:3
	assign stretch_ctrl_enabletx_we = (addr_hit[20] & reg_we) & !reg_error;
	// Trace: design.sv:87564:3
	assign stretch_ctrl_enabletx_wd = reg_wdata[1];
	// Trace: design.sv:87566:3
	assign stretch_ctrl_enableacq_we = (addr_hit[20] & reg_we) & !reg_error;
	// Trace: design.sv:87567:3
	assign stretch_ctrl_enableacq_wd = reg_wdata[2];
	// Trace: design.sv:87569:3
	assign stretch_ctrl_stop_we = (addr_hit[20] & reg_we) & !reg_error;
	// Trace: design.sv:87570:3
	assign stretch_ctrl_stop_wd = reg_wdata[3];
	// Trace: design.sv:87572:3
	assign host_timeout_ctrl_we = (addr_hit[21] & reg_we) & !reg_error;
	// Trace: design.sv:87573:3
	assign host_timeout_ctrl_wd = reg_wdata[31:0];
	// Trace: design.sv:87576:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:87577:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:87578:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]: begin
				// Trace: design.sv:87580:9
				reg_rdata_next[0] = intr_state_fmt_watermark_qs;
				// Trace: design.sv:87581:9
				reg_rdata_next[1] = intr_state_rx_watermark_qs;
				// Trace: design.sv:87582:9
				reg_rdata_next[2] = intr_state_fmt_overflow_qs;
				// Trace: design.sv:87583:9
				reg_rdata_next[3] = intr_state_rx_overflow_qs;
				// Trace: design.sv:87584:9
				reg_rdata_next[4] = intr_state_nak_qs;
				// Trace: design.sv:87585:9
				reg_rdata_next[5] = intr_state_scl_interference_qs;
				// Trace: design.sv:87586:9
				reg_rdata_next[6] = intr_state_sda_interference_qs;
				// Trace: design.sv:87587:9
				reg_rdata_next[7] = intr_state_stretch_timeout_qs;
				// Trace: design.sv:87588:9
				reg_rdata_next[8] = intr_state_sda_unstable_qs;
				// Trace: design.sv:87589:9
				reg_rdata_next[9] = intr_state_trans_complete_qs;
				// Trace: design.sv:87590:9
				reg_rdata_next[10] = intr_state_tx_empty_qs;
				// Trace: design.sv:87591:9
				reg_rdata_next[11] = intr_state_tx_nonempty_qs;
				// Trace: design.sv:87592:9
				reg_rdata_next[12] = intr_state_tx_overflow_qs;
				// Trace: design.sv:87593:9
				reg_rdata_next[13] = intr_state_acq_overflow_qs;
				// Trace: design.sv:87594:9
				reg_rdata_next[14] = intr_state_ack_stop_qs;
				// Trace: design.sv:87595:9
				reg_rdata_next[15] = intr_state_host_timeout_qs;
			end
			addr_hit[1]: begin
				// Trace: design.sv:87599:9
				reg_rdata_next[0] = intr_enable_fmt_watermark_qs;
				// Trace: design.sv:87600:9
				reg_rdata_next[1] = intr_enable_rx_watermark_qs;
				// Trace: design.sv:87601:9
				reg_rdata_next[2] = intr_enable_fmt_overflow_qs;
				// Trace: design.sv:87602:9
				reg_rdata_next[3] = intr_enable_rx_overflow_qs;
				// Trace: design.sv:87603:9
				reg_rdata_next[4] = intr_enable_nak_qs;
				// Trace: design.sv:87604:9
				reg_rdata_next[5] = intr_enable_scl_interference_qs;
				// Trace: design.sv:87605:9
				reg_rdata_next[6] = intr_enable_sda_interference_qs;
				// Trace: design.sv:87606:9
				reg_rdata_next[7] = intr_enable_stretch_timeout_qs;
				// Trace: design.sv:87607:9
				reg_rdata_next[8] = intr_enable_sda_unstable_qs;
				// Trace: design.sv:87608:9
				reg_rdata_next[9] = intr_enable_trans_complete_qs;
				// Trace: design.sv:87609:9
				reg_rdata_next[10] = intr_enable_tx_empty_qs;
				// Trace: design.sv:87610:9
				reg_rdata_next[11] = intr_enable_tx_nonempty_qs;
				// Trace: design.sv:87611:9
				reg_rdata_next[12] = intr_enable_tx_overflow_qs;
				// Trace: design.sv:87612:9
				reg_rdata_next[13] = intr_enable_acq_overflow_qs;
				// Trace: design.sv:87613:9
				reg_rdata_next[14] = intr_enable_ack_stop_qs;
				// Trace: design.sv:87614:9
				reg_rdata_next[15] = intr_enable_host_timeout_qs;
			end
			addr_hit[2]: begin
				// Trace: design.sv:87618:9
				reg_rdata_next[0] = 1'sb0;
				// Trace: design.sv:87619:9
				reg_rdata_next[1] = 1'sb0;
				// Trace: design.sv:87620:9
				reg_rdata_next[2] = 1'sb0;
				// Trace: design.sv:87621:9
				reg_rdata_next[3] = 1'sb0;
				// Trace: design.sv:87622:9
				reg_rdata_next[4] = 1'sb0;
				// Trace: design.sv:87623:9
				reg_rdata_next[5] = 1'sb0;
				// Trace: design.sv:87624:9
				reg_rdata_next[6] = 1'sb0;
				// Trace: design.sv:87625:9
				reg_rdata_next[7] = 1'sb0;
				// Trace: design.sv:87626:9
				reg_rdata_next[8] = 1'sb0;
				// Trace: design.sv:87627:9
				reg_rdata_next[9] = 1'sb0;
				// Trace: design.sv:87628:9
				reg_rdata_next[10] = 1'sb0;
				// Trace: design.sv:87629:9
				reg_rdata_next[11] = 1'sb0;
				// Trace: design.sv:87630:9
				reg_rdata_next[12] = 1'sb0;
				// Trace: design.sv:87631:9
				reg_rdata_next[13] = 1'sb0;
				// Trace: design.sv:87632:9
				reg_rdata_next[14] = 1'sb0;
				// Trace: design.sv:87633:9
				reg_rdata_next[15] = 1'sb0;
			end
			addr_hit[3]: begin
				// Trace: design.sv:87637:9
				reg_rdata_next[0] = ctrl_enablehost_qs;
				// Trace: design.sv:87638:9
				reg_rdata_next[1] = ctrl_enabletarget_qs;
			end
			addr_hit[4]: begin
				// Trace: design.sv:87642:9
				reg_rdata_next[0] = status_fmtfull_qs;
				// Trace: design.sv:87643:9
				reg_rdata_next[1] = status_rxfull_qs;
				// Trace: design.sv:87644:9
				reg_rdata_next[2] = status_fmtempty_qs;
				// Trace: design.sv:87645:9
				reg_rdata_next[3] = status_hostidle_qs;
				// Trace: design.sv:87646:9
				reg_rdata_next[4] = status_targetidle_qs;
				// Trace: design.sv:87647:9
				reg_rdata_next[5] = status_rxempty_qs;
				// Trace: design.sv:87648:9
				reg_rdata_next[6] = status_txfull_qs;
				// Trace: design.sv:87649:9
				reg_rdata_next[7] = status_acqfull_qs;
				// Trace: design.sv:87650:9
				reg_rdata_next[8] = status_txempty_qs;
				// Trace: design.sv:87651:9
				reg_rdata_next[9] = status_acqempty_qs;
			end
			addr_hit[5]:
				// Trace: design.sv:87655:9
				reg_rdata_next[7:0] = rdata_qs;
			addr_hit[6]: begin
				// Trace: design.sv:87659:9
				reg_rdata_next[7:0] = 1'sb0;
				// Trace: design.sv:87660:9
				reg_rdata_next[8] = 1'sb0;
				// Trace: design.sv:87661:9
				reg_rdata_next[9] = 1'sb0;
				// Trace: design.sv:87662:9
				reg_rdata_next[10] = 1'sb0;
				// Trace: design.sv:87663:9
				reg_rdata_next[11] = 1'sb0;
				// Trace: design.sv:87664:9
				reg_rdata_next[12] = 1'sb0;
			end
			addr_hit[7]: begin
				// Trace: design.sv:87668:9
				reg_rdata_next[0] = 1'sb0;
				// Trace: design.sv:87669:9
				reg_rdata_next[1] = 1'sb0;
				// Trace: design.sv:87670:9
				reg_rdata_next[4:2] = fifo_ctrl_rxilvl_qs;
				// Trace: design.sv:87671:9
				reg_rdata_next[6:5] = fifo_ctrl_fmtilvl_qs;
				// Trace: design.sv:87672:9
				reg_rdata_next[7] = 1'sb0;
				// Trace: design.sv:87673:9
				reg_rdata_next[8] = 1'sb0;
			end
			addr_hit[8]: begin
				// Trace: design.sv:87677:9
				reg_rdata_next[5:0] = fifo_status_fmtlvl_qs;
				// Trace: design.sv:87678:9
				reg_rdata_next[13:8] = fifo_status_txlvl_qs;
				// Trace: design.sv:87679:9
				reg_rdata_next[21:16] = fifo_status_rxlvl_qs;
				// Trace: design.sv:87680:9
				reg_rdata_next[29:24] = fifo_status_acqlvl_qs;
			end
			addr_hit[9]: begin
				// Trace: design.sv:87684:9
				reg_rdata_next[0] = ovrd_txovrden_qs;
				// Trace: design.sv:87685:9
				reg_rdata_next[1] = ovrd_sclval_qs;
				// Trace: design.sv:87686:9
				reg_rdata_next[2] = ovrd_sdaval_qs;
			end
			addr_hit[10]: begin
				// Trace: design.sv:87690:9
				reg_rdata_next[15:0] = val_scl_rx_qs;
				// Trace: design.sv:87691:9
				reg_rdata_next[31:16] = val_sda_rx_qs;
			end
			addr_hit[11]: begin
				// Trace: design.sv:87695:9
				reg_rdata_next[15:0] = timing0_thigh_qs;
				// Trace: design.sv:87696:9
				reg_rdata_next[31:16] = timing0_tlow_qs;
			end
			addr_hit[12]: begin
				// Trace: design.sv:87700:9
				reg_rdata_next[15:0] = timing1_t_r_qs;
				// Trace: design.sv:87701:9
				reg_rdata_next[31:16] = timing1_t_f_qs;
			end
			addr_hit[13]: begin
				// Trace: design.sv:87705:9
				reg_rdata_next[15:0] = timing2_tsu_sta_qs;
				// Trace: design.sv:87706:9
				reg_rdata_next[31:16] = timing2_thd_sta_qs;
			end
			addr_hit[14]: begin
				// Trace: design.sv:87710:9
				reg_rdata_next[15:0] = timing3_tsu_dat_qs;
				// Trace: design.sv:87711:9
				reg_rdata_next[31:16] = timing3_thd_dat_qs;
			end
			addr_hit[15]: begin
				// Trace: design.sv:87715:9
				reg_rdata_next[15:0] = timing4_tsu_sto_qs;
				// Trace: design.sv:87716:9
				reg_rdata_next[31:16] = timing4_t_buf_qs;
			end
			addr_hit[16]: begin
				// Trace: design.sv:87720:9
				reg_rdata_next[30:0] = timeout_ctrl_val_qs;
				// Trace: design.sv:87721:9
				reg_rdata_next[31] = timeout_ctrl_en_qs;
			end
			addr_hit[17]: begin
				// Trace: design.sv:87725:9
				reg_rdata_next[6:0] = target_id_address0_qs;
				// Trace: design.sv:87726:9
				reg_rdata_next[13:7] = target_id_mask0_qs;
				// Trace: design.sv:87727:9
				reg_rdata_next[20:14] = target_id_address1_qs;
				// Trace: design.sv:87728:9
				reg_rdata_next[27:21] = target_id_mask1_qs;
			end
			addr_hit[18]: begin
				// Trace: design.sv:87732:9
				reg_rdata_next[7:0] = acqdata_abyte_qs;
				// Trace: design.sv:87733:9
				reg_rdata_next[9:8] = acqdata_signal_qs;
			end
			addr_hit[19]:
				// Trace: design.sv:87737:9
				reg_rdata_next[7:0] = 1'sb0;
			addr_hit[20]: begin
				// Trace: design.sv:87741:9
				reg_rdata_next[0] = stretch_ctrl_enableaddr_qs;
				// Trace: design.sv:87742:9
				reg_rdata_next[1] = stretch_ctrl_enabletx_qs;
				// Trace: design.sv:87743:9
				reg_rdata_next[2] = stretch_ctrl_enableacq_qs;
				// Trace: design.sv:87744:9
				reg_rdata_next[3] = stretch_ctrl_stop_qs;
			end
			addr_hit[21]:
				// Trace: design.sv:87748:9
				reg_rdata_next[31:0] = host_timeout_ctrl_qs;
			default:
				// Trace: design.sv:87752:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:87761:3
	wire unused_wdata;
	// Trace: design.sv:87762:3
	wire unused_be;
	// Trace: design.sv:87763:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:87764:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module i2c_core (
	clk_i,
	rst_ni,
	reg2hw,
	hw2reg,
	scl_i,
	scl_o,
	sda_i,
	sda_o,
	intr_fmt_watermark_o,
	intr_rx_watermark_o,
	intr_fmt_overflow_o,
	intr_rx_overflow_o,
	intr_nak_o,
	intr_scl_interference_o,
	intr_sda_interference_o,
	intr_stretch_timeout_o,
	intr_sda_unstable_o,
	intr_trans_complete_o,
	intr_tx_empty_o,
	intr_tx_nonempty_o,
	intr_tx_overflow_o,
	intr_acq_overflow_o,
	intr_ack_stop_o,
	intr_host_timeout_o
);
	reg _sv2v_0;
	// Trace: design.sv:87786:3
	input clk_i;
	// Trace: design.sv:87787:3
	input rst_ni;
	// Trace: design.sv:87789:3
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_acqdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_fdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_fifo_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_host_timeout_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_enable_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_state_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_test_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_ovrd_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_rdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_stretch_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_target_id_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timeout_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing0_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing1_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing2_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing3_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing4_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_txdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_t
	input wire [388:0] reg2hw;
	// Trace: design.sv:87790:3
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_acqdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_fifo_status_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_intr_state_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_rdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_status_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_val_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_t
	output wire [115:0] hw2reg;
	// Trace: design.sv:87792:3
	input scl_i;
	// Trace: design.sv:87793:3
	output wire scl_o;
	// Trace: design.sv:87794:3
	input sda_i;
	// Trace: design.sv:87795:3
	output wire sda_o;
	// Trace: design.sv:87797:3
	output wire intr_fmt_watermark_o;
	// Trace: design.sv:87798:3
	output wire intr_rx_watermark_o;
	// Trace: design.sv:87799:3
	output wire intr_fmt_overflow_o;
	// Trace: design.sv:87800:3
	output wire intr_rx_overflow_o;
	// Trace: design.sv:87801:3
	output wire intr_nak_o;
	// Trace: design.sv:87802:3
	output wire intr_scl_interference_o;
	// Trace: design.sv:87803:3
	output wire intr_sda_interference_o;
	// Trace: design.sv:87804:3
	output wire intr_stretch_timeout_o;
	// Trace: design.sv:87805:3
	output wire intr_sda_unstable_o;
	// Trace: design.sv:87806:3
	output wire intr_trans_complete_o;
	// Trace: design.sv:87807:3
	output wire intr_tx_empty_o;
	// Trace: design.sv:87808:3
	output wire intr_tx_nonempty_o;
	// Trace: design.sv:87809:3
	output wire intr_tx_overflow_o;
	// Trace: design.sv:87810:3
	output wire intr_acq_overflow_o;
	// Trace: design.sv:87811:3
	output wire intr_ack_stop_o;
	// Trace: design.sv:87812:3
	output wire intr_host_timeout_o;
	// Trace: design.sv:87815:3
	wire [15:0] thigh;
	// Trace: design.sv:87816:3
	wire [15:0] tlow;
	// Trace: design.sv:87817:3
	wire [15:0] t_r;
	// Trace: design.sv:87818:3
	wire [15:0] t_f;
	// Trace: design.sv:87819:3
	wire [15:0] thd_sta;
	// Trace: design.sv:87820:3
	wire [15:0] tsu_sta;
	// Trace: design.sv:87821:3
	wire [15:0] tsu_sto;
	// Trace: design.sv:87822:3
	wire [15:0] tsu_dat;
	// Trace: design.sv:87823:3
	wire [15:0] thd_dat;
	// Trace: design.sv:87824:3
	wire [15:0] t_buf;
	// Trace: design.sv:87825:3
	wire [30:0] stretch_timeout;
	// Trace: design.sv:87826:3
	wire timeout_enable;
	// Trace: design.sv:87827:3
	wire stretch_en_addr;
	// Trace: design.sv:87828:3
	wire stretch_en_tx;
	// Trace: design.sv:87829:3
	wire stretch_en_acq;
	// Trace: design.sv:87830:3
	wire stretch_stop;
	// Trace: design.sv:87831:3
	wire [31:0] host_timeout;
	// Trace: design.sv:87833:3
	wire scl_out_fsm;
	// Trace: design.sv:87834:3
	wire sda_out_fsm;
	// Trace: design.sv:87836:3
	wire event_fmt_watermark;
	// Trace: design.sv:87837:3
	wire event_rx_watermark;
	// Trace: design.sv:87838:3
	wire event_fmt_overflow;
	// Trace: design.sv:87839:3
	wire event_rx_overflow;
	// Trace: design.sv:87840:3
	wire event_nak;
	// Trace: design.sv:87841:3
	wire event_scl_interference;
	// Trace: design.sv:87842:3
	wire event_sda_interference;
	// Trace: design.sv:87843:3
	wire event_stretch_timeout;
	// Trace: design.sv:87844:3
	wire event_sda_unstable;
	// Trace: design.sv:87845:3
	wire event_trans_complete;
	// Trace: design.sv:87846:3
	wire event_tx_empty;
	// Trace: design.sv:87847:3
	wire event_tx_nonempty;
	// Trace: design.sv:87848:3
	wire event_tx_overflow;
	// Trace: design.sv:87849:3
	wire event_acq_overflow;
	// Trace: design.sv:87850:3
	wire event_ack_stop;
	// Trace: design.sv:87851:3
	wire event_host_timeout;
	// Trace: design.sv:87853:3
	reg [15:0] scl_rx_val;
	// Trace: design.sv:87854:3
	reg [15:0] sda_rx_val;
	// Trace: design.sv:87856:3
	wire override;
	// Trace: design.sv:87858:3
	wire fmt_fifo_wvalid;
	// Trace: design.sv:87859:3
	wire fmt_fifo_wready;
	// Trace: design.sv:87860:3
	wire [12:0] fmt_fifo_wdata;
	// Trace: design.sv:87861:3
	wire [5:0] fmt_fifo_depth;
	// Trace: design.sv:87862:3
	wire fmt_fifo_rvalid;
	// Trace: design.sv:87863:3
	wire fmt_fifo_rready;
	// Trace: design.sv:87864:3
	wire [12:0] fmt_fifo_rdata;
	// Trace: design.sv:87865:3
	wire [7:0] fmt_byte;
	// Trace: design.sv:87866:3
	wire fmt_flag_start_before;
	// Trace: design.sv:87867:3
	wire fmt_flag_stop_after;
	// Trace: design.sv:87868:3
	wire fmt_flag_read_bytes;
	// Trace: design.sv:87869:3
	wire fmt_flag_read_continue;
	// Trace: design.sv:87870:3
	wire fmt_flag_nak_ok;
	// Trace: design.sv:87872:3
	wire i2c_fifo_rxrst;
	// Trace: design.sv:87873:3
	wire i2c_fifo_fmtrst;
	// Trace: design.sv:87874:3
	wire [2:0] i2c_fifo_rxilvl;
	// Trace: design.sv:87875:3
	wire [1:0] i2c_fifo_fmtilvl;
	// Trace: design.sv:87877:3
	wire rx_fifo_wvalid;
	// Trace: design.sv:87878:3
	wire rx_fifo_wready;
	// Trace: design.sv:87879:3
	wire [7:0] rx_fifo_wdata;
	// Trace: design.sv:87880:3
	wire [5:0] rx_fifo_depth;
	// Trace: design.sv:87881:3
	wire rx_fifo_rvalid;
	// Trace: design.sv:87882:3
	wire rx_fifo_rready;
	// Trace: design.sv:87883:3
	wire [7:0] rx_fifo_rdata;
	// Trace: design.sv:87885:3
	reg fmt_watermark_d;
	// Trace: design.sv:87886:3
	reg fmt_watermark_q;
	// Trace: design.sv:87887:3
	reg rx_watermark_d;
	// Trace: design.sv:87888:3
	reg rx_watermark_q;
	// Trace: design.sv:87890:3
	wire tx_fifo_wvalid;
	// Trace: design.sv:87891:3
	wire tx_fifo_wready;
	// Trace: design.sv:87892:3
	wire [7:0] tx_fifo_wdata;
	// Trace: design.sv:87893:3
	wire [5:0] tx_fifo_depth;
	// Trace: design.sv:87894:3
	wire tx_fifo_rvalid;
	// Trace: design.sv:87895:3
	wire tx_fifo_rready;
	// Trace: design.sv:87896:3
	wire [7:0] tx_fifo_rdata;
	// Trace: design.sv:87898:3
	wire acq_fifo_wvalid;
	// Trace: design.sv:87899:3
	wire acq_fifo_wready;
	// Trace: design.sv:87900:3
	wire [9:0] acq_fifo_wdata;
	// Trace: design.sv:87901:3
	wire [5:0] acq_fifo_depth;
	// Trace: design.sv:87902:3
	wire acq_fifo_rvalid;
	// Trace: design.sv:87903:3
	wire acq_fifo_rready;
	// Trace: design.sv:87904:3
	wire [9:0] acq_fifo_rdata;
	// Trace: design.sv:87906:3
	wire i2c_fifo_txrst;
	// Trace: design.sv:87907:3
	wire i2c_fifo_acqrst;
	// Trace: design.sv:87909:3
	wire host_idle;
	// Trace: design.sv:87910:3
	wire target_idle;
	// Trace: design.sv:87912:3
	wire host_enable;
	// Trace: design.sv:87913:3
	wire target_enable;
	// Trace: design.sv:87915:3
	wire [6:0] target_address0;
	// Trace: design.sv:87916:3
	wire [6:0] target_mask0;
	// Trace: design.sv:87917:3
	wire [6:0] target_address1;
	// Trace: design.sv:87918:3
	wire [6:0] target_mask1;
	// Trace: design.sv:87921:3
	wire unused_fifo_ctrl_rxilvl_qe;
	// Trace: design.sv:87922:3
	wire unused_fifo_ctrl_fmtilvl_qe;
	// Trace: design.sv:87923:3
	wire [7:0] unused_rx_fifo_rdata_q;
	// Trace: design.sv:87924:3
	wire [7:0] unused_acq_fifo_adata_q;
	// Trace: design.sv:87925:3
	wire [1:0] unused_acq_fifo_signal_q;
	// Trace: design.sv:87927:3
	assign hw2reg[83] = ~fmt_fifo_wready;
	// Trace: design.sv:87928:3
	assign hw2reg[82] = ~rx_fifo_wready;
	// Trace: design.sv:87929:3
	assign hw2reg[81] = ~fmt_fifo_rvalid;
	// Trace: design.sv:87930:3
	assign hw2reg[80] = host_idle;
	// Trace: design.sv:87931:3
	assign hw2reg[79] = target_idle;
	// Trace: design.sv:87932:3
	assign hw2reg[78] = ~rx_fifo_rvalid;
	// Trace: design.sv:87933:3
	assign hw2reg[73-:8] = rx_fifo_rdata;
	// Trace: design.sv:87934:3
	assign hw2reg[65-:6] = fmt_fifo_depth;
	// Trace: design.sv:87935:3
	assign hw2reg[53-:6] = rx_fifo_depth;
	// Trace: design.sv:87936:3
	assign hw2reg[41-:16] = scl_rx_val;
	// Trace: design.sv:87937:3
	assign hw2reg[25-:16] = sda_rx_val;
	// Trace: design.sv:87939:3
	assign hw2reg[77] = ~tx_fifo_wready;
	// Trace: design.sv:87940:3
	assign hw2reg[76] = ~acq_fifo_wready;
	// Trace: design.sv:87941:3
	assign hw2reg[75] = ~tx_fifo_rvalid;
	// Trace: design.sv:87942:3
	assign hw2reg[74] = ~acq_fifo_rvalid;
	// Trace: design.sv:87943:3
	assign hw2reg[59-:6] = tx_fifo_depth;
	// Trace: design.sv:87944:3
	assign hw2reg[47-:6] = acq_fifo_depth;
	// Trace: design.sv:87945:3
	assign hw2reg[9-:8] = acq_fifo_rdata[7:0];
	// Trace: design.sv:87946:3
	assign hw2reg[1-:2] = acq_fifo_rdata[9:8];
	// Trace: design.sv:87948:3
	assign override = reg2hw[279];
	// Trace: design.sv:87950:3
	assign scl_o = (override ? reg2hw[278] : scl_out_fsm);
	// Trace: design.sv:87951:3
	assign sda_o = (override ? reg2hw[277] : sda_out_fsm);
	// Trace: design.sv:87953:3
	assign host_enable = reg2hw[324];
	// Trace: design.sv:87954:3
	assign target_enable = reg2hw[323];
	// Trace: design.sv:87956:3
	assign target_address0 = reg2hw[84-:7];
	// Trace: design.sv:87957:3
	assign target_mask0 = reg2hw[77-:7];
	// Trace: design.sv:87958:3
	assign target_address1 = reg2hw[70-:7];
	// Trace: design.sv:87959:3
	assign target_mask1 = reg2hw[63-:7];
	// Trace: design.sv:87962:3
	always @(posedge clk_i or negedge rst_ni) begin : rx_oversampling
		// Trace: design.sv:87963:5
		if (!rst_ni) begin
			// Trace: design.sv:87964:8
			scl_rx_val <= 16'h0000;
			// Trace: design.sv:87965:8
			sda_rx_val <= 16'h0000;
		end
		else begin
			// Trace: design.sv:87967:8
			scl_rx_val <= {scl_rx_val[14:0], scl_i};
			// Trace: design.sv:87968:8
			sda_rx_val <= {sda_rx_val[14:0], sda_i};
		end
	end
	// Trace: design.sv:87972:3
	assign thigh = reg2hw[276-:16];
	// Trace: design.sv:87973:3
	assign tlow = reg2hw[260-:16];
	// Trace: design.sv:87974:3
	assign t_r = reg2hw[244-:16];
	// Trace: design.sv:87975:3
	assign t_f = reg2hw[228-:16];
	// Trace: design.sv:87976:3
	assign tsu_sta = reg2hw[212-:16];
	// Trace: design.sv:87977:3
	assign thd_sta = reg2hw[196-:16];
	// Trace: design.sv:87978:3
	assign tsu_dat = reg2hw[180-:16];
	// Trace: design.sv:87979:3
	assign thd_dat = reg2hw[164-:16];
	// Trace: design.sv:87980:3
	assign tsu_sto = reg2hw[148-:16];
	// Trace: design.sv:87981:3
	assign t_buf = reg2hw[132-:16];
	// Trace: design.sv:87982:3
	assign stretch_timeout = reg2hw[116-:31];
	// Trace: design.sv:87983:3
	assign timeout_enable = reg2hw[85];
	// Trace: design.sv:87984:3
	assign stretch_en_addr = reg2hw[35];
	// Trace: design.sv:87985:3
	assign stretch_en_tx = reg2hw[34];
	// Trace: design.sv:87986:3
	assign stretch_en_acq = reg2hw[33];
	// Trace: design.sv:87987:3
	assign stretch_stop = reg2hw[32];
	// Trace: design.sv:87988:3
	assign host_timeout = reg2hw[31-:32];
	// Trace: design.sv:87990:3
	assign i2c_fifo_rxrst = reg2hw[294] & reg2hw[293];
	// Trace: design.sv:87991:3
	assign i2c_fifo_fmtrst = reg2hw[292] & reg2hw[291];
	// Trace: design.sv:87992:3
	assign i2c_fifo_rxilvl = reg2hw[290-:3];
	// Trace: design.sv:87993:3
	assign i2c_fifo_fmtilvl = reg2hw[286-:2];
	// Trace: design.sv:87995:3
	assign i2c_fifo_txrst = reg2hw[281] & reg2hw[280];
	// Trace: design.sv:87996:3
	assign i2c_fifo_acqrst = reg2hw[283] & reg2hw[282];
	// Trace: design.sv:87998:3
	always @(posedge clk_i or negedge rst_ni) begin : watermark_transition
		// Trace: design.sv:87999:5
		if (!rst_ni) begin
			// Trace: design.sv:88000:7
			fmt_watermark_q <= 1'b1;
			// Trace: design.sv:88001:7
			rx_watermark_q <= 1'b0;
		end
		else begin
			// Trace: design.sv:88003:7
			fmt_watermark_q <= fmt_watermark_d;
			// Trace: design.sv:88004:7
			rx_watermark_q <= rx_watermark_d;
		end
	end
	// Trace: design.sv:88008:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:88009:5
		(* full_case, parallel_case *)
		case (i2c_fifo_fmtilvl)
			2'h0:
				// Trace: design.sv:88010:16
				fmt_watermark_d = fmt_fifo_depth <= 6'd1;
			2'h1:
				// Trace: design.sv:88011:16
				fmt_watermark_d = fmt_fifo_depth <= 6'd4;
			2'h2:
				// Trace: design.sv:88012:16
				fmt_watermark_d = fmt_fifo_depth <= 6'd8;
			default:
				// Trace: design.sv:88013:16
				fmt_watermark_d = fmt_fifo_depth <= 6'd16;
		endcase
	end
	// Trace: design.sv:88017:3
	assign event_fmt_watermark = fmt_watermark_d & ~fmt_watermark_q;
	// Trace: design.sv:88019:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:88020:5
		(* full_case, parallel_case *)
		case (i2c_fifo_rxilvl)
			3'h0:
				// Trace: design.sv:88021:16
				rx_watermark_d = rx_fifo_depth >= 6'd1;
			3'h1:
				// Trace: design.sv:88022:16
				rx_watermark_d = rx_fifo_depth >= 6'd4;
			3'h2:
				// Trace: design.sv:88023:16
				rx_watermark_d = rx_fifo_depth >= 6'd8;
			3'h3:
				// Trace: design.sv:88024:16
				rx_watermark_d = rx_fifo_depth >= 6'd16;
			3'h4:
				// Trace: design.sv:88025:16
				rx_watermark_d = rx_fifo_depth >= 6'd30;
			default:
				// Trace: design.sv:88026:16
				rx_watermark_d = 1'b0;
		endcase
	end
	// Trace: design.sv:88030:3
	assign event_rx_watermark = rx_watermark_d & ~rx_watermark_q;
	// Trace: design.sv:88032:3
	assign event_fmt_overflow = fmt_fifo_wvalid & ~fmt_fifo_wready;
	// Trace: design.sv:88033:3
	assign event_rx_overflow = rx_fifo_wvalid & ~rx_fifo_wready;
	// Trace: design.sv:88038:3
	assign fmt_fifo_wvalid = ((((reg2hw[305] & reg2hw[303]) & reg2hw[301]) & reg2hw[299]) & reg2hw[297]) & reg2hw[295];
	// Trace: design.sv:88044:3
	assign fmt_fifo_wdata[7:0] = reg2hw[313-:8];
	// Trace: design.sv:88045:3
	assign fmt_fifo_wdata[8] = reg2hw[304];
	// Trace: design.sv:88046:3
	assign fmt_fifo_wdata[9] = reg2hw[302];
	// Trace: design.sv:88047:3
	assign fmt_fifo_wdata[10] = reg2hw[300];
	// Trace: design.sv:88048:3
	assign fmt_fifo_wdata[11] = reg2hw[298];
	// Trace: design.sv:88049:3
	assign fmt_fifo_wdata[12] = reg2hw[296];
	// Trace: design.sv:88051:3
	assign fmt_byte = (fmt_fifo_rvalid ? fmt_fifo_rdata[7:0] : {8 {1'sb0}});
	// Trace: design.sv:88052:3
	assign fmt_flag_start_before = (fmt_fifo_rvalid ? fmt_fifo_rdata[8] : 1'b0);
	// Trace: design.sv:88053:3
	assign fmt_flag_stop_after = (fmt_fifo_rvalid ? fmt_fifo_rdata[9] : 1'b0);
	// Trace: design.sv:88054:3
	assign fmt_flag_read_bytes = (fmt_fifo_rvalid ? fmt_fifo_rdata[10] : 1'b0);
	// Trace: design.sv:88055:3
	assign fmt_flag_read_continue = (fmt_fifo_rvalid ? fmt_fifo_rdata[11] : 1'b0);
	// Trace: design.sv:88056:3
	assign fmt_flag_nak_ok = (fmt_fifo_rvalid ? fmt_fifo_rdata[12] : 1'b0);
	// Trace: design.sv:88059:3
	assign unused_fifo_ctrl_rxilvl_qe = reg2hw[287];
	// Trace: design.sv:88060:3
	assign unused_fifo_ctrl_fmtilvl_qe = reg2hw[284];
	// Trace: design.sv:88061:3
	assign unused_rx_fifo_rdata_q = reg2hw[322-:8];
	// Trace: design.sv:88062:3
	assign unused_acq_fifo_adata_q = reg2hw[56-:8];
	// Trace: design.sv:88063:3
	assign unused_acq_fifo_signal_q = reg2hw[47-:2];
	// Trace: design.sv:88065:3
	prim_fifo_sync #(
		.Width(13),
		.Pass(1'b1),
		.Depth(32)
	) u_i2c_fmtfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(i2c_fifo_fmtrst),
		.wvalid_i(fmt_fifo_wvalid),
		.wready_o(fmt_fifo_wready),
		.wdata_i(fmt_fifo_wdata),
		.depth_o(fmt_fifo_depth),
		.rvalid_o(fmt_fifo_rvalid),
		.rready_i(fmt_fifo_rready),
		.rdata_o(fmt_fifo_rdata),
		.full_o()
	);
	// Trace: design.sv:88083:3
	assign rx_fifo_rready = reg2hw[314];
	// Trace: design.sv:88085:3
	prim_fifo_sync #(
		.Width(8),
		.Pass(1'b0),
		.Depth(32)
	) u_i2c_rxfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(i2c_fifo_rxrst),
		.wvalid_i(rx_fifo_wvalid),
		.wready_o(rx_fifo_wready),
		.wdata_i(rx_fifo_wdata),
		.depth_o(rx_fifo_depth),
		.rvalid_o(rx_fifo_rvalid),
		.rready_i(rx_fifo_rready),
		.rdata_o(rx_fifo_rdata),
		.full_o()
	);
	// Trace: design.sv:88104:3
	assign event_tx_overflow = tx_fifo_wvalid & ~tx_fifo_wready;
	// Trace: design.sv:88105:3
	assign event_acq_overflow = acq_fifo_wvalid & ~acq_fifo_wready;
	// Trace: design.sv:88107:3
	assign tx_fifo_wvalid = reg2hw[36];
	// Trace: design.sv:88108:3
	assign tx_fifo_wdata = reg2hw[44-:8];
	// Trace: design.sv:88110:3
	prim_fifo_sync #(
		.Width(8),
		.Pass(1'b1),
		.Depth(32)
	) u_i2c_txfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(i2c_fifo_txrst),
		.wvalid_i(tx_fifo_wvalid),
		.wready_o(tx_fifo_wready),
		.wdata_i(tx_fifo_wdata),
		.depth_o(tx_fifo_depth),
		.rvalid_o(tx_fifo_rvalid),
		.rready_i(tx_fifo_rready),
		.rdata_o(tx_fifo_rdata),
		.full_o()
	);
	// Trace: design.sv:88128:3
	assign acq_fifo_rready = reg2hw[48] & reg2hw[45];
	// Trace: design.sv:88130:3
	prim_fifo_sync #(
		.Width(10),
		.Pass(1'b0),
		.Depth(32)
	) u_i2c_acqfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(i2c_fifo_acqrst),
		.wvalid_i(acq_fifo_wvalid),
		.wready_o(acq_fifo_wready),
		.wdata_i(acq_fifo_wdata),
		.depth_o(acq_fifo_depth),
		.rvalid_o(acq_fifo_rvalid),
		.rready_i(acq_fifo_rready),
		.rdata_o(acq_fifo_rdata),
		.full_o()
	);
	// Trace: design.sv:88148:3
	i2c_fsm u_i2c_fsm(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.scl_i(scl_i),
		.scl_o(scl_out_fsm),
		.sda_i(sda_i),
		.sda_o(sda_out_fsm),
		.host_enable_i(host_enable),
		.target_enable_i(target_enable),
		.fmt_fifo_rvalid_i(fmt_fifo_rvalid),
		.fmt_fifo_wvalid_i(fmt_fifo_wvalid),
		.fmt_fifo_depth_i(fmt_fifo_depth),
		.fmt_fifo_rready_o(fmt_fifo_rready),
		.fmt_byte_i(fmt_byte),
		.fmt_flag_start_before_i(fmt_flag_start_before),
		.fmt_flag_stop_after_i(fmt_flag_stop_after),
		.fmt_flag_read_bytes_i(fmt_flag_read_bytes),
		.fmt_flag_read_continue_i(fmt_flag_read_continue),
		.fmt_flag_nak_ok_i(fmt_flag_nak_ok),
		.rx_fifo_wvalid_o(rx_fifo_wvalid),
		.rx_fifo_wdata_o(rx_fifo_wdata),
		.tx_fifo_rvalid_i(tx_fifo_rvalid),
		.tx_fifo_wvalid_i(tx_fifo_wvalid),
		.tx_fifo_depth_i(tx_fifo_depth),
		.tx_fifo_rready_o(tx_fifo_rready),
		.tx_fifo_rdata_i(tx_fifo_rdata),
		.acq_fifo_wready_i(acq_fifo_wready),
		.acq_fifo_wvalid_o(acq_fifo_wvalid),
		.acq_fifo_wdata_o(acq_fifo_wdata),
		.host_idle_o(host_idle),
		.target_idle_o(target_idle),
		.thigh_i(thigh),
		.tlow_i(tlow),
		.t_r_i(t_r),
		.t_f_i(t_f),
		.thd_sta_i(thd_sta),
		.tsu_sta_i(tsu_sta),
		.tsu_sto_i(tsu_sto),
		.tsu_dat_i(tsu_dat),
		.thd_dat_i(thd_dat),
		.t_buf_i(t_buf),
		.stretch_timeout_i(stretch_timeout),
		.timeout_enable_i(timeout_enable),
		.stretch_en_addr_i(stretch_en_addr),
		.stretch_en_tx_i(stretch_en_tx),
		.stretch_en_acq_i(stretch_en_acq),
		.stretch_stop_i(stretch_stop),
		.host_timeout_i(host_timeout),
		.target_address0_i(target_address0),
		.target_mask0_i(target_mask0),
		.target_address1_i(target_address1),
		.target_mask1_i(target_mask1),
		.event_nak_o(event_nak),
		.event_scl_interference_o(event_scl_interference),
		.event_sda_interference_o(event_sda_interference),
		.event_stretch_timeout_o(event_stretch_timeout),
		.event_sda_unstable_o(event_sda_unstable),
		.event_trans_complete_o(event_trans_complete),
		.event_tx_empty_o(event_tx_empty),
		.event_tx_nonempty_o(event_tx_nonempty),
		.event_ack_stop_o(event_ack_stop),
		.event_host_timeout_o(event_host_timeout)
	);
	// Trace: design.sv:88223:3
	prim_intr_hw #(.Width(1)) intr_hw_fmt_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_fmt_watermark),
		.reg2hw_intr_enable_q_i(reg2hw[372]),
		.reg2hw_intr_test_q_i(reg2hw[356]),
		.reg2hw_intr_test_qe_i(reg2hw[355]),
		.reg2hw_intr_state_q_i(reg2hw[388]),
		.hw2reg_intr_state_de_o(hw2reg[114]),
		.hw2reg_intr_state_d_o(hw2reg[115]),
		.intr_o(intr_fmt_watermark_o)
	);
	// Trace: design.sv:88236:3
	prim_intr_hw #(.Width(1)) intr_hw_rx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_rx_watermark),
		.reg2hw_intr_enable_q_i(reg2hw[371]),
		.reg2hw_intr_test_q_i(reg2hw[354]),
		.reg2hw_intr_test_qe_i(reg2hw[353]),
		.reg2hw_intr_state_q_i(reg2hw[387]),
		.hw2reg_intr_state_de_o(hw2reg[112]),
		.hw2reg_intr_state_d_o(hw2reg[113]),
		.intr_o(intr_rx_watermark_o)
	);
	// Trace: design.sv:88249:3
	prim_intr_hw #(.Width(1)) intr_hw_fmt_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_fmt_overflow),
		.reg2hw_intr_enable_q_i(reg2hw[370]),
		.reg2hw_intr_test_q_i(reg2hw[352]),
		.reg2hw_intr_test_qe_i(reg2hw[351]),
		.reg2hw_intr_state_q_i(reg2hw[386]),
		.hw2reg_intr_state_de_o(hw2reg[110]),
		.hw2reg_intr_state_d_o(hw2reg[111]),
		.intr_o(intr_fmt_overflow_o)
	);
	// Trace: design.sv:88262:3
	prim_intr_hw #(.Width(1)) intr_hw_rx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_rx_overflow),
		.reg2hw_intr_enable_q_i(reg2hw[369]),
		.reg2hw_intr_test_q_i(reg2hw[350]),
		.reg2hw_intr_test_qe_i(reg2hw[349]),
		.reg2hw_intr_state_q_i(reg2hw[385]),
		.hw2reg_intr_state_de_o(hw2reg[108]),
		.hw2reg_intr_state_d_o(hw2reg[109]),
		.intr_o(intr_rx_overflow_o)
	);
	// Trace: design.sv:88275:3
	prim_intr_hw #(.Width(1)) intr_hw_nak(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_nak),
		.reg2hw_intr_enable_q_i(reg2hw[368]),
		.reg2hw_intr_test_q_i(reg2hw[348]),
		.reg2hw_intr_test_qe_i(reg2hw[347]),
		.reg2hw_intr_state_q_i(reg2hw[384]),
		.hw2reg_intr_state_de_o(hw2reg[106]),
		.hw2reg_intr_state_d_o(hw2reg[107]),
		.intr_o(intr_nak_o)
	);
	// Trace: design.sv:88288:3
	prim_intr_hw #(.Width(1)) intr_hw_scl_interference(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_scl_interference),
		.reg2hw_intr_enable_q_i(reg2hw[367]),
		.reg2hw_intr_test_q_i(reg2hw[346]),
		.reg2hw_intr_test_qe_i(reg2hw[345]),
		.reg2hw_intr_state_q_i(reg2hw[383]),
		.hw2reg_intr_state_de_o(hw2reg[104]),
		.hw2reg_intr_state_d_o(hw2reg[105]),
		.intr_o(intr_scl_interference_o)
	);
	// Trace: design.sv:88301:3
	prim_intr_hw #(.Width(1)) intr_hw_sda_interference(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_sda_interference),
		.reg2hw_intr_enable_q_i(reg2hw[366]),
		.reg2hw_intr_test_q_i(reg2hw[344]),
		.reg2hw_intr_test_qe_i(reg2hw[343]),
		.reg2hw_intr_state_q_i(reg2hw[382]),
		.hw2reg_intr_state_de_o(hw2reg[102]),
		.hw2reg_intr_state_d_o(hw2reg[103]),
		.intr_o(intr_sda_interference_o)
	);
	// Trace: design.sv:88314:3
	prim_intr_hw #(.Width(1)) intr_hw_stretch_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_stretch_timeout),
		.reg2hw_intr_enable_q_i(reg2hw[365]),
		.reg2hw_intr_test_q_i(reg2hw[342]),
		.reg2hw_intr_test_qe_i(reg2hw[341]),
		.reg2hw_intr_state_q_i(reg2hw[381]),
		.hw2reg_intr_state_de_o(hw2reg[100]),
		.hw2reg_intr_state_d_o(hw2reg[101]),
		.intr_o(intr_stretch_timeout_o)
	);
	// Trace: design.sv:88327:3
	prim_intr_hw #(.Width(1)) intr_hw_sda_unstable(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_sda_unstable),
		.reg2hw_intr_enable_q_i(reg2hw[364]),
		.reg2hw_intr_test_q_i(reg2hw[340]),
		.reg2hw_intr_test_qe_i(reg2hw[339]),
		.reg2hw_intr_state_q_i(reg2hw[380]),
		.hw2reg_intr_state_de_o(hw2reg[98]),
		.hw2reg_intr_state_d_o(hw2reg[99]),
		.intr_o(intr_sda_unstable_o)
	);
	// Trace: design.sv:88340:3
	prim_intr_hw #(.Width(1)) intr_hw_trans_complete(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_trans_complete),
		.reg2hw_intr_enable_q_i(reg2hw[363]),
		.reg2hw_intr_test_q_i(reg2hw[338]),
		.reg2hw_intr_test_qe_i(reg2hw[337]),
		.reg2hw_intr_state_q_i(reg2hw[379]),
		.hw2reg_intr_state_de_o(hw2reg[96]),
		.hw2reg_intr_state_d_o(hw2reg[97]),
		.intr_o(intr_trans_complete_o)
	);
	// Trace: design.sv:88353:3
	prim_intr_hw #(.Width(1)) intr_hw_tx_empty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_tx_empty),
		.reg2hw_intr_enable_q_i(reg2hw[362]),
		.reg2hw_intr_test_q_i(reg2hw[336]),
		.reg2hw_intr_test_qe_i(reg2hw[335]),
		.reg2hw_intr_state_q_i(reg2hw[378]),
		.hw2reg_intr_state_de_o(hw2reg[94]),
		.hw2reg_intr_state_d_o(hw2reg[95]),
		.intr_o(intr_tx_empty_o)
	);
	// Trace: design.sv:88366:3
	prim_intr_hw #(.Width(1)) intr_hw_tx_nonempty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_tx_nonempty),
		.reg2hw_intr_enable_q_i(reg2hw[361]),
		.reg2hw_intr_test_q_i(reg2hw[334]),
		.reg2hw_intr_test_qe_i(reg2hw[333]),
		.reg2hw_intr_state_q_i(reg2hw[377]),
		.hw2reg_intr_state_de_o(hw2reg[92]),
		.hw2reg_intr_state_d_o(hw2reg[93]),
		.intr_o(intr_tx_nonempty_o)
	);
	// Trace: design.sv:88379:3
	prim_intr_hw #(.Width(1)) intr_hw_tx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_tx_overflow),
		.reg2hw_intr_enable_q_i(reg2hw[360]),
		.reg2hw_intr_test_q_i(reg2hw[332]),
		.reg2hw_intr_test_qe_i(reg2hw[331]),
		.reg2hw_intr_state_q_i(reg2hw[376]),
		.hw2reg_intr_state_de_o(hw2reg[90]),
		.hw2reg_intr_state_d_o(hw2reg[91]),
		.intr_o(intr_tx_overflow_o)
	);
	// Trace: design.sv:88392:3
	prim_intr_hw #(.Width(1)) intr_hw_acq_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_acq_overflow),
		.reg2hw_intr_enable_q_i(reg2hw[359]),
		.reg2hw_intr_test_q_i(reg2hw[330]),
		.reg2hw_intr_test_qe_i(reg2hw[329]),
		.reg2hw_intr_state_q_i(reg2hw[375]),
		.hw2reg_intr_state_de_o(hw2reg[88]),
		.hw2reg_intr_state_d_o(hw2reg[89]),
		.intr_o(intr_acq_overflow_o)
	);
	// Trace: design.sv:88405:3
	prim_intr_hw #(.Width(1)) intr_hw_ack_stop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_ack_stop),
		.reg2hw_intr_enable_q_i(reg2hw[358]),
		.reg2hw_intr_test_q_i(reg2hw[328]),
		.reg2hw_intr_test_qe_i(reg2hw[327]),
		.reg2hw_intr_state_q_i(reg2hw[374]),
		.hw2reg_intr_state_de_o(hw2reg[86]),
		.hw2reg_intr_state_d_o(hw2reg[87]),
		.intr_o(intr_ack_stop_o)
	);
	// Trace: design.sv:88418:3
	prim_intr_hw #(.Width(1)) intr_hw_host_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_host_timeout),
		.reg2hw_intr_enable_q_i(reg2hw[357]),
		.reg2hw_intr_test_q_i(reg2hw[326]),
		.reg2hw_intr_test_qe_i(reg2hw[325]),
		.reg2hw_intr_state_q_i(reg2hw[373]),
		.hw2reg_intr_state_de_o(hw2reg[84]),
		.hw2reg_intr_state_d_o(hw2reg[85]),
		.intr_o(intr_host_timeout_o)
	);
	initial _sv2v_0 = 0;
endmodule
module i2c_fsm (
	clk_i,
	rst_ni,
	scl_i,
	scl_o,
	sda_i,
	sda_o,
	host_enable_i,
	target_enable_i,
	fmt_fifo_rvalid_i,
	fmt_fifo_wvalid_i,
	fmt_fifo_depth_i,
	fmt_fifo_rready_o,
	fmt_byte_i,
	fmt_flag_start_before_i,
	fmt_flag_stop_after_i,
	fmt_flag_read_bytes_i,
	fmt_flag_read_continue_i,
	fmt_flag_nak_ok_i,
	rx_fifo_wvalid_o,
	rx_fifo_wdata_o,
	tx_fifo_rvalid_i,
	tx_fifo_wvalid_i,
	tx_fifo_depth_i,
	tx_fifo_rready_o,
	tx_fifo_rdata_i,
	acq_fifo_wready_i,
	acq_fifo_wvalid_o,
	acq_fifo_wdata_o,
	host_idle_o,
	target_idle_o,
	thigh_i,
	tlow_i,
	t_r_i,
	t_f_i,
	thd_sta_i,
	tsu_sta_i,
	tsu_sto_i,
	tsu_dat_i,
	thd_dat_i,
	t_buf_i,
	stretch_timeout_i,
	timeout_enable_i,
	stretch_en_addr_i,
	stretch_en_tx_i,
	stretch_en_acq_i,
	stretch_stop_i,
	host_timeout_i,
	target_address0_i,
	target_mask0_i,
	target_address1_i,
	target_mask1_i,
	event_nak_o,
	event_scl_interference_o,
	event_sda_interference_o,
	event_stretch_timeout_o,
	event_sda_unstable_o,
	event_trans_complete_o,
	event_tx_empty_o,
	event_tx_nonempty_o,
	event_ack_stop_o,
	event_host_timeout_o
);
	reg _sv2v_0;
	// Trace: design.sv:88441:3
	input clk_i;
	// Trace: design.sv:88442:3
	input rst_ni;
	// Trace: design.sv:88444:3
	input scl_i;
	// Trace: design.sv:88445:3
	output wire scl_o;
	// Trace: design.sv:88446:3
	input sda_i;
	// Trace: design.sv:88447:3
	output wire sda_o;
	// Trace: design.sv:88449:3
	input host_enable_i;
	// Trace: design.sv:88450:3
	input target_enable_i;
	// Trace: design.sv:88452:3
	input fmt_fifo_rvalid_i;
	// Trace: design.sv:88453:3
	input fmt_fifo_wvalid_i;
	// Trace: design.sv:88454:3
	input [5:0] fmt_fifo_depth_i;
	// Trace: design.sv:88455:3
	output reg fmt_fifo_rready_o;
	// Trace: design.sv:88456:3
	input [7:0] fmt_byte_i;
	// Trace: design.sv:88457:3
	input fmt_flag_start_before_i;
	// Trace: design.sv:88458:3
	input fmt_flag_stop_after_i;
	// Trace: design.sv:88459:3
	input fmt_flag_read_bytes_i;
	// Trace: design.sv:88460:3
	input fmt_flag_read_continue_i;
	// Trace: design.sv:88461:3
	input fmt_flag_nak_ok_i;
	// Trace: design.sv:88463:3
	output reg rx_fifo_wvalid_o;
	// Trace: design.sv:88464:3
	output reg [7:0] rx_fifo_wdata_o;
	// Trace: design.sv:88466:3
	input tx_fifo_rvalid_i;
	// Trace: design.sv:88467:3
	input tx_fifo_wvalid_i;
	// Trace: design.sv:88468:3
	input [5:0] tx_fifo_depth_i;
	// Trace: design.sv:88469:3
	output reg tx_fifo_rready_o;
	// Trace: design.sv:88470:3
	input [7:0] tx_fifo_rdata_i;
	// Trace: design.sv:88472:3
	input wire acq_fifo_wready_i;
	// Trace: design.sv:88473:3
	output reg acq_fifo_wvalid_o;
	// Trace: design.sv:88474:3
	output reg [9:0] acq_fifo_wdata_o;
	// Trace: design.sv:88476:3
	output reg host_idle_o;
	// Trace: design.sv:88477:3
	output reg target_idle_o;
	// Trace: design.sv:88479:3
	input [15:0] thigh_i;
	// Trace: design.sv:88480:3
	input [15:0] tlow_i;
	// Trace: design.sv:88481:3
	input [15:0] t_r_i;
	// Trace: design.sv:88482:3
	input [15:0] t_f_i;
	// Trace: design.sv:88483:3
	input [15:0] thd_sta_i;
	// Trace: design.sv:88484:3
	input [15:0] tsu_sta_i;
	// Trace: design.sv:88485:3
	input [15:0] tsu_sto_i;
	// Trace: design.sv:88486:3
	input [15:0] tsu_dat_i;
	// Trace: design.sv:88487:3
	input [15:0] thd_dat_i;
	// Trace: design.sv:88488:3
	input [15:0] t_buf_i;
	// Trace: design.sv:88489:3
	input [30:0] stretch_timeout_i;
	// Trace: design.sv:88490:3
	input timeout_enable_i;
	// Trace: design.sv:88491:3
	input stretch_en_addr_i;
	// Trace: design.sv:88492:3
	input stretch_en_tx_i;
	// Trace: design.sv:88493:3
	input stretch_en_acq_i;
	// Trace: design.sv:88494:3
	input stretch_stop_i;
	// Trace: design.sv:88495:3
	input [31:0] host_timeout_i;
	// Trace: design.sv:88497:3
	input wire [6:0] target_address0_i;
	// Trace: design.sv:88498:3
	input wire [6:0] target_mask0_i;
	// Trace: design.sv:88499:3
	input wire [6:0] target_address1_i;
	// Trace: design.sv:88500:3
	input wire [6:0] target_mask1_i;
	// Trace: design.sv:88502:3
	output reg event_nak_o;
	// Trace: design.sv:88503:3
	output reg event_scl_interference_o;
	// Trace: design.sv:88504:3
	output reg event_sda_interference_o;
	// Trace: design.sv:88505:3
	output reg event_stretch_timeout_o;
	// Trace: design.sv:88506:3
	output reg event_sda_unstable_o;
	// Trace: design.sv:88507:3
	output reg event_trans_complete_o;
	// Trace: design.sv:88508:3
	output reg event_tx_empty_o;
	// Trace: design.sv:88509:3
	output reg event_tx_nonempty_o;
	// Trace: design.sv:88510:3
	output reg event_ack_stop_o;
	// Trace: design.sv:88511:3
	output wire event_host_timeout_o;
	// Trace: design.sv:88515:3
	reg [19:0] tcount_q;
	// Trace: design.sv:88516:3
	reg [19:0] tcount_d;
	// Trace: design.sv:88517:3
	reg load_tcount;
	// Trace: design.sv:88518:3
	reg [30:0] stretch;
	// Trace: design.sv:88521:3
	reg [2:0] bit_index;
	// Trace: design.sv:88522:3
	reg bit_decr;
	// Trace: design.sv:88523:3
	reg bit_clr;
	// Trace: design.sv:88524:3
	reg [8:0] byte_num;
	// Trace: design.sv:88525:3
	reg [8:0] byte_index;
	// Trace: design.sv:88526:3
	reg byte_decr;
	// Trace: design.sv:88527:3
	reg byte_clr;
	// Trace: design.sv:88530:3
	reg scl_temp;
	// Trace: design.sv:88531:3
	reg sda_temp;
	// Trace: design.sv:88532:3
	reg scl_i_q;
	// Trace: design.sv:88533:3
	reg sda_i_q;
	// Trace: design.sv:88534:3
	reg [7:0] read_byte;
	// Trace: design.sv:88535:3
	reg read_byte_clr;
	// Trace: design.sv:88536:3
	reg shift_data_en;
	// Trace: design.sv:88537:3
	reg no_stop;
	// Trace: design.sv:88538:3
	reg log_start;
	// Trace: design.sv:88539:3
	reg log_stop;
	// Trace: design.sv:88540:3
	reg restart;
	// Trace: design.sv:88543:3
	reg start_det;
	// Trace: design.sv:88544:3
	reg stop_det;
	// Trace: design.sv:88545:3
	wire address0_match;
	// Trace: design.sv:88546:3
	wire address1_match;
	// Trace: design.sv:88547:3
	wire address_match;
	// Trace: design.sv:88548:3
	reg [7:0] input_byte;
	// Trace: design.sv:88549:3
	reg input_byte_clr;
	// Trace: design.sv:88550:3
	reg [31:0] scl_high_cnt;
	// Trace: design.sv:88553:3
	reg [3:0] bit_idx;
	// Trace: design.sv:88554:3
	wire bit_ack;
	// Trace: design.sv:88555:3
	wire rw_bit;
	// Trace: design.sv:88556:3
	reg host_ack;
	// Trace: design.sv:88559:3
	// removed localparam type tcount_sel_e
	// Trace: design.sv:88564:3
	reg [3:0] tcount_sel;
	// Trace: design.sv:88566:3
	function automatic [19:0] sv2v_cast_20;
		input reg [19:0] inp;
		sv2v_cast_20 = inp;
	endfunction
	always @(*) begin : counter_functions
		if (_sv2v_0)
			;
		// Trace: design.sv:88567:5
		tcount_d = tcount_q;
		// Trace: design.sv:88568:5
		if (load_tcount)
			// Trace: design.sv:88569:7
			(* full_case, parallel_case *)
			case (tcount_sel)
				4'd0:
					// Trace: design.sv:88570:23
					tcount_d = sv2v_cast_20(t_r_i) + sv2v_cast_20(tsu_sta_i);
				4'd1:
					// Trace: design.sv:88571:23
					tcount_d = sv2v_cast_20(t_f_i) + sv2v_cast_20(thd_sta_i);
				4'd6:
					// Trace: design.sv:88572:23
					tcount_d = sv2v_cast_20(thd_dat_i);
				4'd2:
					// Trace: design.sv:88573:23
					tcount_d = ((sv2v_cast_20(tlow_i) - sv2v_cast_20(t_r_i)) - sv2v_cast_20(tsu_dat_i)) - sv2v_cast_20(thd_dat_i);
				4'd3:
					// Trace: design.sv:88574:23
					tcount_d = sv2v_cast_20(t_r_i) + sv2v_cast_20(tsu_dat_i);
				4'd4:
					// Trace: design.sv:88575:23
					tcount_d = (sv2v_cast_20(t_r_i) + sv2v_cast_20(thigh_i)) + sv2v_cast_20(t_f_i);
				4'd5:
					// Trace: design.sv:88576:23
					tcount_d = sv2v_cast_20(t_f_i) + sv2v_cast_20(thd_dat_i);
				4'd7:
					// Trace: design.sv:88577:23
					tcount_d = (sv2v_cast_20(t_f_i) + sv2v_cast_20(tlow_i)) - sv2v_cast_20(thd_dat_i);
				4'd8:
					// Trace: design.sv:88578:23
					tcount_d = sv2v_cast_20(t_r_i) + sv2v_cast_20(tsu_sto_i);
				4'd9:
					// Trace: design.sv:88579:23
					tcount_d = (sv2v_cast_20(t_r_i) + sv2v_cast_20(t_buf_i)) - sv2v_cast_20(tsu_sta_i);
				4'd10:
					// Trace: design.sv:88580:23
					tcount_d = 20'h00001;
				default:
					// Trace: design.sv:88581:23
					tcount_d = 20'h00001;
			endcase
		else if (stretch == {31 {1'sb0}})
			// Trace: design.sv:88584:7
			tcount_d = tcount_q - 1'b1;
		else
			// Trace: design.sv:88586:7
			tcount_d = tcount_q;
	end
	// Trace: design.sv:88590:3
	always @(posedge clk_i or negedge rst_ni) begin : clk_counter
		// Trace: design.sv:88591:5
		if (!rst_ni)
			// Trace: design.sv:88592:7
			tcount_q <= 1'sb1;
		else
			// Trace: design.sv:88594:7
			tcount_q <= tcount_d;
	end
	// Trace: design.sv:88599:3
	always @(posedge clk_i or negedge rst_ni) begin : clk_stretch
		// Trace: design.sv:88600:5
		if (!rst_ni)
			// Trace: design.sv:88601:7
			stretch <= 1'sb0;
		else if (scl_temp && !scl_i)
			// Trace: design.sv:88603:7
			stretch <= stretch + 1'b1;
		else
			// Trace: design.sv:88605:7
			stretch <= 1'sb0;
	end
	// Trace: design.sv:88610:3
	always @(posedge clk_i or negedge rst_ni) begin : bit_counter
		// Trace: design.sv:88611:5
		if (!rst_ni)
			// Trace: design.sv:88612:7
			bit_index <= 3'd7;
		else if (bit_clr)
			// Trace: design.sv:88614:7
			bit_index <= 3'd7;
		else if (bit_decr)
			// Trace: design.sv:88616:7
			bit_index <= bit_index - 1'b1;
		else
			// Trace: design.sv:88618:7
			bit_index <= bit_index;
	end
	// Trace: design.sv:88623:3
	always @(posedge clk_i or negedge rst_ni) begin : read_register
		// Trace: design.sv:88624:5
		if (!rst_ni)
			// Trace: design.sv:88625:7
			read_byte <= 8'h00;
		else if (read_byte_clr)
			// Trace: design.sv:88627:7
			read_byte <= 8'h00;
		else if (shift_data_en)
			// Trace: design.sv:88629:7
			read_byte[7:0] <= {read_byte[6:0], sda_i};
	end
	// Trace: design.sv:88634:3
	function automatic [8:0] sv2v_cast_9;
		input reg [8:0] inp;
		sv2v_cast_9 = inp;
	endfunction
	always @(*) begin : byte_number
		if (_sv2v_0)
			;
		// Trace: design.sv:88635:5
		if (!fmt_flag_read_bytes_i)
			// Trace: design.sv:88635:33
			byte_num = 9'd0;
		else if (fmt_byte_i == {8 {1'sb0}})
			// Trace: design.sv:88636:32
			byte_num = 9'd256;
		else
			// Trace: design.sv:88637:10
			byte_num = sv2v_cast_9(fmt_byte_i);
	end
	// Trace: design.sv:88641:3
	always @(posedge clk_i or negedge rst_ni) begin : byte_counter
		// Trace: design.sv:88642:5
		if (!rst_ni)
			// Trace: design.sv:88643:7
			byte_index <= 1'sb0;
		else if (byte_clr)
			// Trace: design.sv:88645:7
			byte_index <= byte_num;
		else if (byte_decr)
			// Trace: design.sv:88647:7
			byte_index <= byte_index - 1'b1;
		else
			// Trace: design.sv:88649:7
			byte_index <= byte_index;
	end
	// Trace: design.sv:88654:3
	always @(posedge clk_i or negedge rst_ni) begin : bus_prev
		// Trace: design.sv:88655:5
		if (!rst_ni) begin
			// Trace: design.sv:88656:7
			scl_i_q <= 1'b1;
			// Trace: design.sv:88657:7
			sda_i_q <= 1'b1;
		end
		else begin
			// Trace: design.sv:88659:7
			scl_i_q <= scl_i;
			// Trace: design.sv:88660:7
			sda_i_q <= sda_i;
		end
	end
	// Trace: design.sv:88665:3
	always @(posedge clk_i or negedge rst_ni) begin : stop_state
		// Trace: design.sv:88666:5
		if (!rst_ni)
			// Trace: design.sv:88667:7
			no_stop <= 1'b0;
		else if (log_stop)
			// Trace: design.sv:88669:7
			no_stop <= 1'b0;
		else if (log_start)
			// Trace: design.sv:88671:7
			no_stop <= 1'b1;
		else
			// Trace: design.sv:88673:7
			no_stop <= no_stop;
	end
	// Trace: design.sv:88678:3
	always @(posedge clk_i or negedge rst_ni) begin : s_detect
		// Trace: design.sv:88679:5
		if (!rst_ni)
			// Trace: design.sv:88680:7
			start_det <= 1'b0;
		else if (scl_i_q && scl_i) begin
			begin
				// Trace: design.sv:88682:7
				if (sda_i_q && !sda_i)
					// Trace: design.sv:88682:30
					start_det <= 1'b1;
				else
					// Trace: design.sv:88683:12
					start_det <= 1'b0;
			end
		end
		else
			// Trace: design.sv:88685:7
			start_det <= 1'b0;
	end
	// Trace: design.sv:88690:3
	always @(posedge clk_i or negedge rst_ni) begin : p_detect
		// Trace: design.sv:88691:5
		if (!rst_ni)
			// Trace: design.sv:88692:7
			stop_det <= 1'b0;
		else if (scl_i_q && scl_i) begin
			begin
				// Trace: design.sv:88694:7
				if (!sda_i_q && sda_i)
					// Trace: design.sv:88694:30
					stop_det <= 1'b1;
				else
					// Trace: design.sv:88695:12
					stop_det <= 1'b0;
			end
		end
		else
			// Trace: design.sv:88697:7
			stop_det <= 1'b0;
	end
	// Trace: design.sv:88702:3
	assign bit_ack = (bit_idx == 4'd8) && !start_det;
	// Trace: design.sv:88705:3
	always @(posedge clk_i or negedge rst_ni) begin : tgt_bit_counter
		// Trace: design.sv:88706:5
		if (!rst_ni)
			// Trace: design.sv:88707:7
			bit_idx <= 4'd0;
		else if (start_det || bit_ack)
			// Trace: design.sv:88709:7
			bit_idx <= 4'd0;
		else if (scl_i_q && !scl_i)
			// Trace: design.sv:88711:7
			bit_idx <= bit_idx + 1'b1;
		else
			// Trace: design.sv:88713:7
			bit_idx <= bit_idx;
	end
	// Trace: design.sv:88718:3
	always @(posedge clk_i or negedge rst_ni) begin : scl_high_counter
		// Trace: design.sv:88719:5
		if (!rst_ni)
			// Trace: design.sv:88720:7
			scl_high_cnt <= 32'd0;
		else if (scl_i)
			// Trace: design.sv:88722:7
			scl_high_cnt <= scl_high_cnt + 1'b1;
		else
			// Trace: design.sv:88724:7
			scl_high_cnt <= 32'd0;
	end
	// Trace: design.sv:88729:3
	assign address0_match = (input_byte[7:1] & target_mask0_i) == target_address0_i;
	// Trace: design.sv:88730:3
	assign address1_match = (input_byte[7:1] & target_mask1_i) == target_address1_i;
	// Trace: design.sv:88731:3
	assign address_match = address0_match || address1_match;
	// Trace: design.sv:88732:3
	assign rw_bit = input_byte[0];
	// Trace: design.sv:88735:3
	always @(posedge clk_i or negedge rst_ni) begin : tgt_input_register
		// Trace: design.sv:88736:5
		if (!rst_ni)
			// Trace: design.sv:88737:7
			input_byte <= 8'h00;
		else if (input_byte_clr)
			// Trace: design.sv:88739:7
			input_byte <= 8'h00;
		else if (!scl_i_q && scl_i) begin
			begin
				// Trace: design.sv:88741:7
				if (!bit_ack)
					// Trace: design.sv:88741:21
					input_byte[7:0] <= {input_byte[6:0], sda_i};
			end
		end
	end
	// Trace: design.sv:88746:3
	always @(posedge clk_i or negedge rst_ni) begin : host_ack_register
		// Trace: design.sv:88747:5
		if (!rst_ni)
			// Trace: design.sv:88748:7
			host_ack <= 1'b0;
		else if (!scl_i_q && scl_i) begin
			begin
				// Trace: design.sv:88750:7
				if (bit_ack)
					// Trace: design.sv:88750:20
					host_ack <= ~sda_i;
			end
		end
	end
	// Trace: design.sv:88755:3
	// removed localparam type state_e
	// Trace: design.sv:88769:3
	reg [5:0] state_q;
	reg [5:0] state_d;
	// Trace: design.sv:88772:3
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	always @(*) begin : state_outputs
		if (_sv2v_0)
			;
		// Trace: design.sv:88773:5
		host_idle_o = 1'b1;
		// Trace: design.sv:88774:5
		target_idle_o = 1'b1;
		// Trace: design.sv:88775:5
		sda_temp = 1'b1;
		// Trace: design.sv:88776:5
		scl_temp = 1'b1;
		// Trace: design.sv:88777:5
		fmt_fifo_rready_o = 1'b0;
		// Trace: design.sv:88778:5
		rx_fifo_wvalid_o = 1'b0;
		// Trace: design.sv:88779:5
		rx_fifo_wdata_o = 8'h00;
		// Trace: design.sv:88780:5
		tx_fifo_rready_o = 1'b0;
		// Trace: design.sv:88781:5
		acq_fifo_wvalid_o = 1'b0;
		// Trace: design.sv:88782:5
		acq_fifo_wdata_o = 10'b0000000000;
		// Trace: design.sv:88783:5
		event_nak_o = 1'b0;
		// Trace: design.sv:88784:5
		event_scl_interference_o = 1'b0;
		// Trace: design.sv:88785:5
		event_sda_interference_o = 1'b0;
		// Trace: design.sv:88786:5
		event_sda_unstable_o = 1'b0;
		// Trace: design.sv:88787:5
		event_stretch_timeout_o = 1'b0;
		// Trace: design.sv:88788:5
		event_trans_complete_o = 1'b0;
		// Trace: design.sv:88789:5
		event_tx_empty_o = 1'b0;
		// Trace: design.sv:88790:5
		event_tx_nonempty_o = 1'b0;
		// Trace: design.sv:88791:5
		event_ack_stop_o = 1'b0;
		// Trace: design.sv:88792:5
		(* full_case, parallel_case *)
		case (state_q)
			6'd0: begin
				// Trace: design.sv:88795:9
				host_idle_o = 1'b1;
				// Trace: design.sv:88796:9
				sda_temp = 1'b1;
				// Trace: design.sv:88797:9
				scl_temp = 1'b1;
				// Trace: design.sv:88798:9
				if (host_enable_i && !sda_i)
					// Trace: design.sv:88798:38
					event_sda_interference_o = 1'b1;
			end
			6'd2: begin
				// Trace: design.sv:88802:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88803:9
				sda_temp = 1'b1;
				// Trace: design.sv:88804:9
				scl_temp = 1'b1;
				// Trace: design.sv:88805:9
				if (!sda_i)
					// Trace: design.sv:88805:21
					event_sda_interference_o = 1'b1;
				if (restart)
					// Trace: design.sv:88806:22
					event_trans_complete_o = 1'b1;
			end
			6'd3: begin
				// Trace: design.sv:88810:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88811:9
				sda_temp = 1'b0;
				// Trace: design.sv:88812:9
				scl_temp = 1'b1;
			end
			6'd23: begin
				// Trace: design.sv:88816:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88817:9
				sda_temp = 1'b0;
				// Trace: design.sv:88818:9
				scl_temp = 1'b0;
			end
			6'd6: begin
				// Trace: design.sv:88822:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88823:9
				sda_temp = 1'b0;
				// Trace: design.sv:88824:9
				scl_temp = 1'b0;
			end
			6'd7: begin
				// Trace: design.sv:88828:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88829:9
				sda_temp = fmt_byte_i[bit_index];
				// Trace: design.sv:88830:9
				scl_temp = 1'b0;
				// Trace: design.sv:88831:9
				if (sda_temp && !sda_i)
					// Trace: design.sv:88831:33
					event_sda_interference_o = 1'b1;
			end
			6'd8: begin
				// Trace: design.sv:88835:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88836:9
				sda_temp = fmt_byte_i[bit_index];
				// Trace: design.sv:88837:9
				scl_temp = 1'b1;
				// Trace: design.sv:88838:9
				if ((stretch > stretch_timeout_i) && timeout_enable_i)
					// Trace: design.sv:88839:11
					event_stretch_timeout_o = 1'b1;
				if (scl_i_q && !scl_i)
					// Trace: design.sv:88841:33
					event_scl_interference_o = 1'b1;
				if (sda_temp && !sda_i)
					// Trace: design.sv:88842:33
					event_sda_interference_o = 1'b1;
				if (sda_i_q != sda_i)
					// Trace: design.sv:88843:33
					event_sda_unstable_o = 1'b1;
			end
			6'd9: begin
				// Trace: design.sv:88847:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88848:9
				sda_temp = fmt_byte_i[bit_index];
				// Trace: design.sv:88849:9
				scl_temp = 1'b0;
				// Trace: design.sv:88850:9
				if (sda_temp && !sda_i)
					// Trace: design.sv:88850:33
					event_sda_interference_o = 1'b1;
			end
			6'd10: begin
				// Trace: design.sv:88854:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88855:9
				sda_temp = 1'b0;
				// Trace: design.sv:88856:9
				scl_temp = 1'b0;
			end
			6'd11: begin
				// Trace: design.sv:88860:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88861:9
				sda_temp = 1'b1;
				// Trace: design.sv:88862:9
				scl_temp = 1'b0;
			end
			6'd12: begin
				// Trace: design.sv:88866:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88867:9
				sda_temp = 1'b1;
				// Trace: design.sv:88868:9
				scl_temp = 1'b1;
				// Trace: design.sv:88869:9
				if (!sda_i && !fmt_flag_nak_ok_i)
					// Trace: design.sv:88869:43
					event_nak_o = 1'b1;
				if ((stretch > stretch_timeout_i) && timeout_enable_i)
					// Trace: design.sv:88871:11
					event_stretch_timeout_o = 1'b1;
				if (scl_i_q && !scl_i)
					// Trace: design.sv:88873:33
					event_scl_interference_o = 1'b1;
				if (sda_i_q != sda_i)
					// Trace: design.sv:88874:33
					event_sda_unstable_o = 1'b1;
			end
			6'd13: begin
				// Trace: design.sv:88878:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88879:9
				sda_temp = 1'b1;
				// Trace: design.sv:88880:9
				scl_temp = 1'b0;
			end
			6'd14: begin
				// Trace: design.sv:88884:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88885:9
				sda_temp = 1'b1;
				// Trace: design.sv:88886:9
				scl_temp = 1'b0;
			end
			6'd15: begin
				// Trace: design.sv:88890:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88891:9
				scl_temp = 1'b0;
			end
			6'd16: begin
				// Trace: design.sv:88895:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88896:9
				scl_temp = 1'b1;
				// Trace: design.sv:88897:9
				if ((stretch > stretch_timeout_i) && timeout_enable_i)
					// Trace: design.sv:88898:11
					event_stretch_timeout_o = 1'b1;
				if (scl_i_q && !scl_i)
					// Trace: design.sv:88900:33
					event_scl_interference_o = 1'b1;
				if (sda_i_q != sda_i)
					// Trace: design.sv:88901:33
					event_sda_unstable_o = 1'b1;
			end
			6'd17: begin
				// Trace: design.sv:88905:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88906:9
				scl_temp = 1'b0;
				// Trace: design.sv:88907:9
				if ((bit_index == {3 {1'sb0}}) && (tcount_q == 20'd1)) begin
					// Trace: design.sv:88908:11
					rx_fifo_wdata_o = read_byte;
					// Trace: design.sv:88909:11
					rx_fifo_wvalid_o = 1'b1;
				end
			end
			6'd18: begin
				// Trace: design.sv:88914:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88915:9
				sda_temp = 1'b0;
				// Trace: design.sv:88916:9
				scl_temp = 1'b0;
			end
			6'd19: begin
				// Trace: design.sv:88920:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88921:9
				if (fmt_flag_read_continue_i)
					// Trace: design.sv:88921:39
					sda_temp = 1'b0;
				else if (byte_index == 9'd1)
					// Trace: design.sv:88922:38
					sda_temp = 1'b1;
				else
					// Trace: design.sv:88923:14
					sda_temp = 1'b0;
				// Trace: design.sv:88924:9
				scl_temp = 1'b0;
				if (sda_temp && !sda_i)
					// Trace: design.sv:88925:33
					event_sda_interference_o = 1'b1;
			end
			6'd20: begin
				// Trace: design.sv:88929:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88930:9
				if (fmt_flag_read_continue_i)
					// Trace: design.sv:88930:39
					sda_temp = 1'b0;
				else if (byte_index == 9'd1)
					// Trace: design.sv:88931:38
					sda_temp = 1'b1;
				else
					// Trace: design.sv:88932:14
					sda_temp = 1'b0;
				// Trace: design.sv:88933:9
				scl_temp = 1'b1;
				if ((stretch > stretch_timeout_i) && timeout_enable_i)
					// Trace: design.sv:88935:11
					event_stretch_timeout_o = 1'b1;
				if (scl_i_q && !scl_i)
					// Trace: design.sv:88937:33
					event_scl_interference_o = 1'b1;
				if (sda_temp && !sda_i)
					// Trace: design.sv:88938:33
					event_sda_interference_o = 1'b1;
				if (sda_i_q != sda_i)
					// Trace: design.sv:88939:33
					event_sda_unstable_o = 1'b1;
			end
			6'd21: begin
				// Trace: design.sv:88943:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88944:9
				if (fmt_flag_read_continue_i)
					// Trace: design.sv:88944:39
					sda_temp = 1'b0;
				else if (byte_index == 9'd1)
					// Trace: design.sv:88945:38
					sda_temp = 1'b1;
				else
					// Trace: design.sv:88946:14
					sda_temp = 1'b0;
				// Trace: design.sv:88947:9
				scl_temp = 1'b0;
				if (sda_temp && !sda_i)
					// Trace: design.sv:88948:33
					event_sda_interference_o = 1'b1;
			end
			6'd24: begin
				// Trace: design.sv:88952:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88953:9
				sda_temp = 1'b0;
				// Trace: design.sv:88954:9
				scl_temp = 1'b0;
			end
			6'd4: begin
				// Trace: design.sv:88958:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88959:9
				sda_temp = 1'b0;
				// Trace: design.sv:88960:9
				scl_temp = 1'b1;
			end
			6'd5: begin
				// Trace: design.sv:88964:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88965:9
				sda_temp = 1'b1;
				// Trace: design.sv:88966:9
				scl_temp = 1'b1;
				// Trace: design.sv:88967:9
				if (!sda_i)
					// Trace: design.sv:88967:21
					event_sda_interference_o = 1'b1;
				// Trace: design.sv:88968:9
				event_trans_complete_o = 1'b1;
			end
			6'd22: begin
				// Trace: design.sv:88972:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88973:9
				scl_temp = 1'b0;
			end
			6'd1: begin
				// Trace: design.sv:88977:9
				host_idle_o = 1'b0;
				// Trace: design.sv:88978:9
				if (fmt_flag_stop_after_i)
					// Trace: design.sv:88978:36
					scl_temp = 1'b1;
				else
					// Trace: design.sv:88979:14
					scl_temp = 1'b0;
				// Trace: design.sv:88980:9
				fmt_fifo_rready_o = 1'b1;
			end
			6'd25: begin
				// Trace: design.sv:88984:9
				target_idle_o = 1'b0;
				// Trace: design.sv:88985:9
				if (bit_ack && address_match) begin
					// Trace: design.sv:88986:11
					acq_fifo_wdata_o = {2'b01, input_byte};
					// Trace: design.sv:88987:11
					acq_fifo_wvalid_o = 1'b1;
					// Trace: design.sv:88988:11
					if ((tx_fifo_depth_i == {6 {1'sb0}}) && rw_bit)
						// Trace: design.sv:88988:48
						event_tx_empty_o = 1'b1;
				end
			end
			6'd26:
				// Trace: design.sv:88993:9
				target_idle_o = 1'b0;
			6'd27: begin
				// Trace: design.sv:88997:9
				target_idle_o = 1'b0;
				// Trace: design.sv:88998:9
				sda_temp = 1'b0;
			end
			6'd28: begin
				// Trace: design.sv:89002:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89003:9
				sda_temp = 1'b0;
			end
			6'd29: begin
				// Trace: design.sv:89007:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89008:9
				sda_temp = 1'b0;
			end
			6'd30:
				// Trace: design.sv:89012:9
				target_idle_o = 1'b0;
			6'd31: begin
				// Trace: design.sv:89016:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89017:9
				sda_temp = tx_fifo_rdata_i[sv2v_cast_3(bit_idx)];
			end
			6'd32: begin
				// Trace: design.sv:89021:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89022:9
				sda_temp = tx_fifo_rdata_i[sv2v_cast_3(bit_idx)];
			end
			6'd33: begin
				// Trace: design.sv:89026:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89027:9
				sda_temp = tx_fifo_rdata_i[sv2v_cast_3(bit_idx)];
			end
			6'd34: begin
				// Trace: design.sv:89031:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89032:9
				if (((tx_fifo_depth_i == 6'd1) && !tx_fifo_wvalid_i) && host_ack)
					// Trace: design.sv:89032:71
					event_tx_empty_o = 1'b1;
				if (host_ack && (start_det || stop_det))
					// Trace: design.sv:89033:50
					event_ack_stop_o = 1'b1;
			end
			6'd40: begin
				// Trace: design.sv:89037:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89038:9
				tx_fifo_rready_o = 1'b1;
			end
			6'd35: begin
				// Trace: design.sv:89042:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89043:9
				if (bit_ack) begin
					// Trace: design.sv:89044:11
					acq_fifo_wdata_o = {2'b00, input_byte};
					// Trace: design.sv:89045:11
					acq_fifo_wvalid_o = 1'b1;
				end
			end
			6'd36:
				// Trace: design.sv:89050:9
				target_idle_o = 1'b0;
			6'd37: begin
				// Trace: design.sv:89054:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89055:9
				sda_temp = 1'b0;
			end
			6'd38: begin
				// Trace: design.sv:89059:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89060:9
				sda_temp = 1'b0;
			end
			6'd39: begin
				// Trace: design.sv:89064:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89065:9
				sda_temp = 1'b0;
			end
			6'd41: begin
				// Trace: design.sv:89069:9
				if (start_det)
					// Trace: design.sv:89069:24
					acq_fifo_wdata_o = {2'b11, input_byte};
				else
					// Trace: design.sv:89070:14
					acq_fifo_wdata_o = {2'b10, input_byte};
				// Trace: design.sv:89071:9
				acq_fifo_wvalid_o = 1'b1;
				if (tx_fifo_depth_i != {6 {1'sb0}})
					// Trace: design.sv:89072:36
					event_tx_nonempty_o = 1'b1;
			end
			6'd44: begin
				// Trace: design.sv:89076:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89077:9
				scl_temp = 1'b0;
			end
			6'd45: begin
				// Trace: design.sv:89081:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89082:9
				scl_temp = 1'b0;
			end
			6'd46: begin
				// Trace: design.sv:89086:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89087:9
				scl_temp = 1'b0;
			end
			6'd42: begin
				// Trace: design.sv:89091:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89092:9
				tx_fifo_rready_o = 1'b1;
				// Trace: design.sv:89093:9
				scl_temp = 1'b0;
				// Trace: design.sv:89094:9
				if (tx_fifo_depth_i == {6 {1'sb0}})
					// Trace: design.sv:89094:36
					event_tx_empty_o = 1'b1;
			end
			6'd43: begin
				// Trace: design.sv:89098:9
				target_idle_o = 1'b0;
				// Trace: design.sv:89099:9
				scl_temp = 1'b0;
			end
			default: begin
				// Trace: design.sv:89103:9
				host_idle_o = 1'b1;
				// Trace: design.sv:89104:9
				target_idle_o = 1'b1;
				// Trace: design.sv:89105:9
				sda_temp = 1'b1;
				// Trace: design.sv:89106:9
				scl_temp = 1'b1;
				// Trace: design.sv:89107:9
				fmt_fifo_rready_o = 1'b0;
				// Trace: design.sv:89108:9
				rx_fifo_wvalid_o = 1'b0;
				// Trace: design.sv:89109:9
				rx_fifo_wdata_o = 8'h00;
				// Trace: design.sv:89110:9
				tx_fifo_rready_o = 1'b0;
				// Trace: design.sv:89111:9
				acq_fifo_wvalid_o = 1'b0;
				// Trace: design.sv:89112:9
				acq_fifo_wdata_o = 10'b0000000000;
				// Trace: design.sv:89113:9
				event_nak_o = 1'b0;
				// Trace: design.sv:89114:9
				event_scl_interference_o = 1'b0;
				// Trace: design.sv:89115:9
				event_sda_interference_o = 1'b0;
				// Trace: design.sv:89116:9
				event_sda_unstable_o = 1'b0;
				// Trace: design.sv:89117:9
				event_stretch_timeout_o = 1'b0;
				// Trace: design.sv:89118:9
				event_trans_complete_o = 1'b0;
				// Trace: design.sv:89119:9
				event_tx_empty_o = 1'b0;
				// Trace: design.sv:89120:9
				event_tx_nonempty_o = 1'b0;
				// Trace: design.sv:89121:9
				event_ack_stop_o = 1'b0;
			end
		endcase
	end
	// Trace: design.sv:89127:3
	always @(*) begin : state_functions
		if (_sv2v_0)
			;
		// Trace: design.sv:89128:5
		state_d = state_q;
		// Trace: design.sv:89129:5
		load_tcount = 1'b0;
		// Trace: design.sv:89130:5
		tcount_sel = 4'd10;
		// Trace: design.sv:89131:5
		bit_decr = 1'b0;
		// Trace: design.sv:89132:5
		bit_clr = 1'b0;
		// Trace: design.sv:89133:5
		byte_decr = 1'b0;
		// Trace: design.sv:89134:5
		byte_clr = 1'b0;
		// Trace: design.sv:89135:5
		read_byte_clr = 1'b0;
		// Trace: design.sv:89136:5
		shift_data_en = 1'b0;
		// Trace: design.sv:89137:5
		log_start = 1'b0;
		// Trace: design.sv:89138:5
		log_stop = 1'b0;
		// Trace: design.sv:89139:5
		restart = 1'b0;
		// Trace: design.sv:89140:5
		input_byte_clr = 1'b0;
		// Trace: design.sv:89142:5
		(* full_case, parallel_case *)
		case (state_q)
			6'd0:
				// Trace: design.sv:89145:9
				if (!host_enable_i && !target_enable_i)
					// Trace: design.sv:89145:49
					state_d = 6'd0;
				else if (host_enable_i) begin
					begin
						// Trace: design.sv:89147:11
						if (!fmt_fifo_rvalid_i)
							// Trace: design.sv:89147:35
							state_d = 6'd0;
						else
							// Trace: design.sv:89148:16
							state_d = 6'd22;
					end
				end
				else if (target_enable_i) begin
					begin
						// Trace: design.sv:89150:11
						if (!start_det)
							// Trace: design.sv:89150:27
							state_d = 6'd0;
						else begin
							// Trace: design.sv:89152:13
							state_d = 6'd25;
							// Trace: design.sv:89153:13
							input_byte_clr = 1'b1;
						end
					end
				end
			6'd2: begin
				// Trace: design.sv:89160:9
				if (no_stop)
					// Trace: design.sv:89160:22
					restart = 1'b1;
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89162:11
					state_d = 6'd3;
					// Trace: design.sv:89163:11
					load_tcount = 1'b1;
					// Trace: design.sv:89164:11
					tcount_sel = 4'd1;
					// Trace: design.sv:89165:11
					log_start = 1'b1;
				end
			end
			6'd3:
				// Trace: design.sv:89170:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89171:11
					state_d = 6'd23;
					// Trace: design.sv:89172:11
					load_tcount = 1'b1;
					// Trace: design.sv:89173:11
					tcount_sel = 4'd6;
				end
			6'd23:
				// Trace: design.sv:89178:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89179:11
					state_d = 6'd6;
					// Trace: design.sv:89180:11
					load_tcount = 1'b1;
					// Trace: design.sv:89181:11
					tcount_sel = 4'd2;
				end
			6'd6:
				// Trace: design.sv:89187:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89188:11
					state_d = 6'd7;
					// Trace: design.sv:89189:11
					load_tcount = 1'b1;
					// Trace: design.sv:89190:11
					tcount_sel = 4'd3;
				end
			6'd7:
				// Trace: design.sv:89195:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89196:11
					state_d = 6'd8;
					// Trace: design.sv:89197:11
					load_tcount = 1'b1;
					// Trace: design.sv:89198:11
					tcount_sel = 4'd4;
				end
			6'd8:
				// Trace: design.sv:89203:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89204:11
					state_d = 6'd9;
					// Trace: design.sv:89205:11
					load_tcount = 1'b1;
					// Trace: design.sv:89206:11
					tcount_sel = 4'd5;
				end
			6'd9:
				// Trace: design.sv:89211:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89212:11
					load_tcount = 1'b1;
					// Trace: design.sv:89213:11
					tcount_sel = 4'd2;
					// Trace: design.sv:89214:11
					if (bit_index == {3 {1'sb0}}) begin
						// Trace: design.sv:89215:13
						state_d = 6'd10;
						// Trace: design.sv:89216:13
						bit_clr = 1'b1;
					end
					else begin
						// Trace: design.sv:89218:13
						state_d = 6'd6;
						// Trace: design.sv:89219:13
						bit_decr = 1'b1;
					end
				end
			6'd10:
				// Trace: design.sv:89226:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89227:11
					state_d = 6'd11;
					// Trace: design.sv:89228:11
					load_tcount = 1'b1;
					// Trace: design.sv:89229:11
					tcount_sel = 4'd3;
				end
			6'd11:
				// Trace: design.sv:89234:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89235:11
					state_d = 6'd12;
					// Trace: design.sv:89236:11
					load_tcount = 1'b1;
					// Trace: design.sv:89237:11
					tcount_sel = 4'd4;
				end
			6'd12:
				// Trace: design.sv:89242:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89243:11
					state_d = 6'd13;
					// Trace: design.sv:89244:11
					load_tcount = 1'b1;
					// Trace: design.sv:89245:11
					tcount_sel = 4'd5;
				end
			6'd13:
				// Trace: design.sv:89250:9
				if (tcount_q == 20'd1) begin
					begin
						// Trace: design.sv:89251:11
						if (fmt_flag_stop_after_i) begin
							// Trace: design.sv:89252:13
							state_d = 6'd24;
							// Trace: design.sv:89253:13
							load_tcount = 1'b1;
							// Trace: design.sv:89254:13
							tcount_sel = 4'd7;
						end
						else begin
							// Trace: design.sv:89256:13
							state_d = 6'd1;
							// Trace: design.sv:89257:13
							load_tcount = 1'b1;
							// Trace: design.sv:89258:13
							tcount_sel = 4'd10;
						end
					end
				end
			6'd14:
				// Trace: design.sv:89265:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89266:11
					state_d = 6'd15;
					// Trace: design.sv:89267:11
					load_tcount = 1'b1;
					// Trace: design.sv:89268:11
					tcount_sel = 4'd3;
				end
			6'd15:
				// Trace: design.sv:89273:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89274:11
					state_d = 6'd16;
					// Trace: design.sv:89275:11
					load_tcount = 1'b1;
					// Trace: design.sv:89276:11
					tcount_sel = 4'd4;
				end
			6'd16:
				// Trace: design.sv:89281:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89282:11
					state_d = 6'd17;
					// Trace: design.sv:89283:11
					load_tcount = 1'b1;
					// Trace: design.sv:89284:11
					tcount_sel = 4'd5;
					// Trace: design.sv:89285:11
					shift_data_en = 1'b1;
				end
			6'd17:
				// Trace: design.sv:89290:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89291:11
					load_tcount = 1'b1;
					// Trace: design.sv:89292:11
					tcount_sel = 4'd2;
					// Trace: design.sv:89293:11
					if (bit_index == {3 {1'sb0}}) begin
						// Trace: design.sv:89294:13
						state_d = 6'd18;
						// Trace: design.sv:89295:13
						bit_clr = 1'b1;
						// Trace: design.sv:89296:13
						read_byte_clr = 1'b1;
					end
					else begin
						// Trace: design.sv:89298:13
						state_d = 6'd14;
						// Trace: design.sv:89299:13
						bit_decr = 1'b1;
					end
				end
			6'd18:
				// Trace: design.sv:89306:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89307:11
					state_d = 6'd19;
					// Trace: design.sv:89308:11
					load_tcount = 1'b1;
					// Trace: design.sv:89309:11
					tcount_sel = 4'd3;
				end
			6'd19:
				// Trace: design.sv:89314:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89315:11
					state_d = 6'd20;
					// Trace: design.sv:89316:11
					load_tcount = 1'b1;
					// Trace: design.sv:89317:11
					tcount_sel = 4'd4;
				end
			6'd20:
				// Trace: design.sv:89322:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89323:11
					state_d = 6'd21;
					// Trace: design.sv:89324:11
					load_tcount = 1'b1;
					// Trace: design.sv:89325:11
					tcount_sel = 4'd5;
				end
			6'd21:
				// Trace: design.sv:89330:9
				if (tcount_q == 20'd1) begin
					begin
						// Trace: design.sv:89331:11
						if (byte_index == 9'd1) begin
							begin
								// Trace: design.sv:89332:13
								if (fmt_flag_stop_after_i) begin
									// Trace: design.sv:89333:15
									state_d = 6'd24;
									// Trace: design.sv:89334:15
									load_tcount = 1'b1;
									// Trace: design.sv:89335:15
									tcount_sel = 4'd7;
								end
								else begin
									// Trace: design.sv:89337:15
									state_d = 6'd1;
									// Trace: design.sv:89338:15
									load_tcount = 1'b1;
									// Trace: design.sv:89339:15
									tcount_sel = 4'd10;
								end
							end
						end
						else begin
							// Trace: design.sv:89342:13
							state_d = 6'd14;
							// Trace: design.sv:89343:13
							load_tcount = 1'b1;
							// Trace: design.sv:89344:13
							tcount_sel = 4'd2;
							// Trace: design.sv:89345:13
							byte_decr = 1'b1;
						end
					end
				end
			6'd24:
				// Trace: design.sv:89352:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89353:11
					state_d = 6'd4;
					// Trace: design.sv:89354:11
					load_tcount = 1'b1;
					// Trace: design.sv:89355:11
					tcount_sel = 4'd8;
				end
			6'd4:
				// Trace: design.sv:89360:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89361:11
					state_d = 6'd5;
					// Trace: design.sv:89362:11
					load_tcount = 1'b1;
					// Trace: design.sv:89363:11
					tcount_sel = 4'd9;
					// Trace: design.sv:89364:11
					log_stop = 1'b1;
				end
			6'd5:
				// Trace: design.sv:89369:9
				if (tcount_q == 20'd1) begin
					begin
						// Trace: design.sv:89370:11
						if (!host_enable_i) begin
							// Trace: design.sv:89371:13
							state_d = 6'd0;
							// Trace: design.sv:89372:13
							load_tcount = 1'b1;
							// Trace: design.sv:89373:13
							tcount_sel = 4'd10;
						end
						else begin
							// Trace: design.sv:89375:13
							state_d = 6'd1;
							// Trace: design.sv:89376:13
							load_tcount = 1'b1;
							// Trace: design.sv:89377:13
							tcount_sel = 4'd10;
						end
					end
				end
			6'd22:
				// Trace: design.sv:89384:9
				if (fmt_flag_read_bytes_i) begin
					// Trace: design.sv:89385:11
					byte_clr = 1'b1;
					// Trace: design.sv:89386:11
					state_d = 6'd14;
					// Trace: design.sv:89387:11
					load_tcount = 1'b1;
					// Trace: design.sv:89388:11
					tcount_sel = 4'd2;
				end
				else if (fmt_flag_start_before_i) begin
					// Trace: design.sv:89390:11
					state_d = 6'd2;
					// Trace: design.sv:89391:11
					load_tcount = 1'b1;
					// Trace: design.sv:89392:11
					tcount_sel = 4'd0;
				end
				else begin
					// Trace: design.sv:89394:11
					state_d = 6'd6;
					// Trace: design.sv:89395:11
					load_tcount = 1'b1;
					// Trace: design.sv:89396:11
					tcount_sel = 4'd2;
				end
			6'd1:
				// Trace: design.sv:89402:9
				if (!host_enable_i) begin
					// Trace: design.sv:89403:11
					state_d = 6'd24;
					// Trace: design.sv:89404:11
					load_tcount = 1'b1;
					// Trace: design.sv:89405:11
					tcount_sel = 4'd7;
				end
				else if ((fmt_fifo_depth_i == 6'd1) && !fmt_fifo_wvalid_i) begin
					// Trace: design.sv:89407:11
					state_d = 6'd0;
					// Trace: design.sv:89408:11
					load_tcount = 1'b1;
					// Trace: design.sv:89409:11
					tcount_sel = 4'd10;
				end
				else begin
					// Trace: design.sv:89411:11
					state_d = 6'd22;
					// Trace: design.sv:89412:11
					load_tcount = 1'b1;
					// Trace: design.sv:89413:11
					tcount_sel = 4'd10;
				end
			6'd25:
				// Trace: design.sv:89419:9
				if (bit_ack) begin
					begin
						// Trace: design.sv:89420:11
						if (address_match) begin
							// Trace: design.sv:89421:13
							state_d = 6'd26;
							// Trace: design.sv:89422:13
							load_tcount = 1'b1;
							// Trace: design.sv:89423:13
							tcount_sel = 4'd6;
						end
						else
							// Trace: design.sv:89424:20
							state_d = 6'd0;
					end
				end
			6'd26:
				// Trace: design.sv:89430:9
				if (tcount_q == 20'd1) begin
					begin
						// Trace: design.sv:89431:11
						if (stretch_en_addr_i)
							// Trace: design.sv:89431:34
							state_d = 6'd44;
						else
							// Trace: design.sv:89432:16
							state_d = 6'd27;
					end
				end
			6'd27:
				// Trace: design.sv:89437:9
				if (scl_i)
					// Trace: design.sv:89437:20
					state_d = 6'd28;
			6'd28:
				// Trace: design.sv:89441:9
				if (!scl_i) begin
					// Trace: design.sv:89442:11
					state_d = 6'd29;
					// Trace: design.sv:89443:11
					load_tcount = 1'b1;
					// Trace: design.sv:89444:11
					tcount_sel = 4'd6;
				end
			6'd29:
				// Trace: design.sv:89449:9
				if (tcount_q == 20'd1) begin
					begin
						// Trace: design.sv:89450:11
						if (rw_bit) begin
							begin
								// Trace: design.sv:89451:13
								if (tx_fifo_rvalid_i) begin
									// Trace: design.sv:89452:15
									state_d = 6'd30;
									// Trace: design.sv:89453:15
									load_tcount = 1'b1;
									// Trace: design.sv:89454:15
									tcount_sel = 4'd2;
								end
								else
									// Trace: design.sv:89455:22
									state_d = 6'd42;
							end
						end
						else
							// Trace: design.sv:89457:13
							if (acq_fifo_wready_i)
								// Trace: design.sv:89457:36
								state_d = 6'd35;
							else
								// Trace: design.sv:89458:18
								state_d = 6'd43;
					end
				end
			6'd30:
				// Trace: design.sv:89465:9
				if (tcount_q == 20'd1)
					// Trace: design.sv:89466:11
					state_d = 6'd31;
			6'd31:
				// Trace: design.sv:89471:9
				if (scl_i)
					// Trace: design.sv:89471:20
					state_d = 6'd32;
			6'd32:
				// Trace: design.sv:89475:9
				if (!scl_i) begin
					// Trace: design.sv:89476:11
					state_d = 6'd33;
					// Trace: design.sv:89477:11
					load_tcount = 1'b1;
					// Trace: design.sv:89478:11
					tcount_sel = 4'd6;
				end
			6'd33:
				// Trace: design.sv:89483:9
				if (tcount_q == 20'd1) begin
					// Trace: design.sv:89484:11
					load_tcount = 1'b1;
					// Trace: design.sv:89485:11
					tcount_sel = 4'd2;
					// Trace: design.sv:89486:11
					if (bit_ack)
						// Trace: design.sv:89487:13
						state_d = 6'd34;
					else
						// Trace: design.sv:89489:13
						state_d = 6'd30;
				end
			6'd34:
				// Trace: design.sv:89495:9
				if (scl_i) begin
					begin
						// Trace: design.sv:89496:11
						if (host_ack) begin
							begin
								// Trace: design.sv:89497:13
								if (stretch_en_tx_i)
									// Trace: design.sv:89497:34
									state_d = 6'd46;
								else
									// Trace: design.sv:89498:18
									state_d = 6'd40;
							end
						end
						else
							// Trace: design.sv:89500:13
							if (start_det || stop_det)
								// Trace: design.sv:89500:40
								state_d = 6'd41;
					end
				end
			6'd40:
				// Trace: design.sv:89507:9
				if (!target_enable_i)
					// Trace: design.sv:89508:11
					state_d = 6'd0;
				else if ((tx_fifo_depth_i == 6'd1) && !tx_fifo_wvalid_i)
					// Trace: design.sv:89510:11
					state_d = 6'd42;
				else begin
					// Trace: design.sv:89512:11
					state_d = 6'd30;
					// Trace: design.sv:89513:11
					load_tcount = 1'b1;
					// Trace: design.sv:89514:11
					tcount_sel = 4'd2;
				end
			6'd35:
				// Trace: design.sv:89520:9
				if (bit_ack) begin
					// Trace: design.sv:89521:11
					state_d = 6'd36;
					// Trace: design.sv:89522:11
					load_tcount = 1'b1;
					// Trace: design.sv:89523:11
					tcount_sel = 4'd6;
				end
			6'd36:
				// Trace: design.sv:89529:9
				if (tcount_q == 20'd1) begin
					begin
						// Trace: design.sv:89530:11
						if (stretch_en_acq_i)
							// Trace: design.sv:89530:33
							state_d = 6'd45;
						else
							// Trace: design.sv:89531:16
							state_d = 6'd37;
					end
				end
			6'd37:
				// Trace: design.sv:89536:9
				if (scl_i)
					// Trace: design.sv:89536:20
					state_d = 6'd38;
			6'd38:
				// Trace: design.sv:89540:9
				if (!scl_i) begin
					// Trace: design.sv:89541:11
					state_d = 6'd39;
					// Trace: design.sv:89542:11
					load_tcount = 1'b1;
					// Trace: design.sv:89543:11
					tcount_sel = 4'd6;
				end
			6'd39:
				// Trace: design.sv:89548:9
				if (tcount_q == 20'd1) begin
					begin
						// Trace: design.sv:89549:11
						if (bit_ack) begin
							begin
								// Trace: design.sv:89550:13
								if (start_det || stop_det)
									// Trace: design.sv:89550:40
									state_d = 6'd41;
								else
									// Trace: design.sv:89551:18
									state_d = 6'd35;
							end
						end
					end
				end
			6'd41:
				// Trace: design.sv:89558:9
				state_d = 6'd0;
			6'd44:
				// Trace: design.sv:89563:9
				if (!stretch_stop_i)
					// Trace: design.sv:89563:30
					state_d = 6'd44;
				else
					// Trace: design.sv:89564:14
					state_d = 6'd27;
			6'd45:
				// Trace: design.sv:89569:9
				if (!stretch_stop_i)
					// Trace: design.sv:89569:30
					state_d = 6'd45;
				else
					// Trace: design.sv:89570:14
					state_d = 6'd37;
			6'd46:
				// Trace: design.sv:89575:9
				if (!stretch_stop_i)
					// Trace: design.sv:89575:30
					state_d = 6'd46;
				else
					// Trace: design.sv:89576:14
					state_d = 6'd40;
			6'd42:
				// Trace: design.sv:89581:9
				if (tx_fifo_depth_i == {6 {1'sb0}})
					// Trace: design.sv:89582:11
					state_d = 6'd42;
				else begin
					// Trace: design.sv:89584:11
					state_d = 6'd30;
					// Trace: design.sv:89585:11
					load_tcount = 1'b1;
					// Trace: design.sv:89586:11
					tcount_sel = 4'd2;
				end
			6'd43:
				// Trace: design.sv:89592:9
				if (acq_fifo_wready_i)
					// Trace: design.sv:89592:32
					state_d = 6'd35;
				else
					// Trace: design.sv:89593:14
					state_d = 6'd43;
			default: begin
				// Trace: design.sv:89598:9
				state_d = 6'd0;
				// Trace: design.sv:89599:9
				load_tcount = 1'b0;
				// Trace: design.sv:89600:9
				tcount_sel = 4'd10;
				// Trace: design.sv:89601:9
				bit_decr = 1'b0;
				// Trace: design.sv:89602:9
				bit_clr = 1'b0;
				// Trace: design.sv:89603:9
				byte_decr = 1'b0;
				// Trace: design.sv:89604:9
				byte_clr = 1'b0;
				// Trace: design.sv:89605:9
				read_byte_clr = 1'b0;
				// Trace: design.sv:89606:9
				shift_data_en = 1'b0;
				// Trace: design.sv:89607:9
				log_start = 1'b0;
				// Trace: design.sv:89608:9
				log_stop = 1'b0;
				// Trace: design.sv:89609:9
				restart = 1'b0;
				// Trace: design.sv:89610:9
				input_byte_clr = 1'b0;
			end
		endcase
	end
	// Trace: design.sv:89616:3
	always @(posedge clk_i or negedge rst_ni) begin : state_transition
		// Trace: design.sv:89617:5
		if (!rst_ni)
			// Trace: design.sv:89618:7
			state_q <= 6'd0;
		else
			// Trace: design.sv:89620:7
			state_q <= state_d;
	end
	// Trace: design.sv:89625:3
	assign scl_o = scl_temp;
	// Trace: design.sv:89626:3
	assign sda_o = sda_temp;
	// Trace: design.sv:89629:3
	assign event_host_timeout_o = (!target_idle_o & (scl_high_cnt > host_timeout_i) ? 1'b1 : 1'b0);
	initial _sv2v_0 = 0;
endmodule
module i2c (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	cio_scl_i,
	cio_scl_o,
	cio_scl_en_o,
	cio_sda_i,
	cio_sda_o,
	cio_sda_en_o,
	intr_fmt_watermark_o,
	intr_rx_watermark_o,
	intr_fmt_overflow_o,
	intr_rx_overflow_o,
	intr_nak_o,
	intr_scl_interference_o,
	intr_sda_interference_o,
	intr_stretch_timeout_o,
	intr_sda_unstable_o,
	intr_trans_complete_o,
	intr_tx_empty_o,
	intr_tx_nonempty_o,
	intr_tx_overflow_o,
	intr_acq_overflow_o,
	intr_ack_stop_o,
	intr_host_timeout_o
);
	// Trace: design.sv:89641:3
	input clk_i;
	// Trace: design.sv:89642:3
	input rst_ni;
	// Trace: design.sv:89645:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:89646:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:89649:3
	input cio_scl_i;
	// Trace: design.sv:89650:3
	output wire cio_scl_o;
	// Trace: design.sv:89651:3
	output wire cio_scl_en_o;
	// Trace: design.sv:89652:3
	input cio_sda_i;
	// Trace: design.sv:89653:3
	output wire cio_sda_o;
	// Trace: design.sv:89654:3
	output wire cio_sda_en_o;
	// Trace: design.sv:89657:3
	output wire intr_fmt_watermark_o;
	// Trace: design.sv:89658:3
	output wire intr_rx_watermark_o;
	// Trace: design.sv:89659:3
	output wire intr_fmt_overflow_o;
	// Trace: design.sv:89660:3
	output wire intr_rx_overflow_o;
	// Trace: design.sv:89661:3
	output wire intr_nak_o;
	// Trace: design.sv:89662:3
	output wire intr_scl_interference_o;
	// Trace: design.sv:89663:3
	output wire intr_sda_interference_o;
	// Trace: design.sv:89664:3
	output wire intr_stretch_timeout_o;
	// Trace: design.sv:89665:3
	output wire intr_sda_unstable_o;
	// Trace: design.sv:89666:3
	output wire intr_trans_complete_o;
	// Trace: design.sv:89667:3
	output wire intr_tx_empty_o;
	// Trace: design.sv:89668:3
	output wire intr_tx_nonempty_o;
	// Trace: design.sv:89669:3
	output wire intr_tx_overflow_o;
	// Trace: design.sv:89670:3
	output wire intr_acq_overflow_o;
	// Trace: design.sv:89671:3
	output wire intr_ack_stop_o;
	// Trace: design.sv:89672:3
	output wire intr_host_timeout_o;
	// Trace: design.sv:89675:3
	// removed import i2c_reg_pkg::*;
	// Trace: design.sv:89677:3
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_acqdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_fdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_fifo_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_host_timeout_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_enable_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_state_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_intr_test_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_ovrd_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_rdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_stretch_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_target_id_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timeout_ctrl_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing0_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing1_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing2_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing3_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_timing4_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_txdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_reg2hw_t
	wire [388:0] reg2hw;
	// Trace: design.sv:89678:3
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_acqdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_fifo_status_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_intr_state_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_rdata_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_status_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_val_reg_t
	// removed localparam type i2c_reg_pkg_i2c_hw2reg_t
	wire [115:0] hw2reg;
	// Trace: design.sv:89680:3
	i2c_reg_top u_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.tl_o(tl_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.intg_err_o(),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:89691:3
	wire scl_int;
	// Trace: design.sv:89692:3
	wire sda_int;
	// Trace: design.sv:89694:3
	i2c_core i2c_core(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.scl_i(cio_scl_i),
		.scl_o(scl_int),
		.sda_i(cio_sda_i),
		.sda_o(sda_int),
		.intr_fmt_watermark_o(intr_fmt_watermark_o),
		.intr_rx_watermark_o(intr_rx_watermark_o),
		.intr_fmt_overflow_o(intr_fmt_overflow_o),
		.intr_rx_overflow_o(intr_rx_overflow_o),
		.intr_nak_o(intr_nak_o),
		.intr_scl_interference_o(intr_scl_interference_o),
		.intr_sda_interference_o(intr_sda_interference_o),
		.intr_stretch_timeout_o(intr_stretch_timeout_o),
		.intr_sda_unstable_o(intr_sda_unstable_o),
		.intr_trans_complete_o(intr_trans_complete_o),
		.intr_tx_empty_o(intr_tx_empty_o),
		.intr_tx_nonempty_o(intr_tx_nonempty_o),
		.intr_tx_overflow_o(intr_tx_overflow_o),
		.intr_acq_overflow_o(intr_acq_overflow_o),
		.intr_ack_stop_o(intr_ack_stop_o),
		.intr_host_timeout_o(intr_host_timeout_o)
	);
	// Trace: design.sv:89727:3
	assign cio_scl_o = 1'b0;
	// Trace: design.sv:89728:3
	assign cio_sda_o = 1'b0;
	// Trace: design.sv:89730:3
	assign cio_scl_en_o = ~scl_int;
	// Trace: design.sv:89731:3
	assign cio_sda_en_o = ~sda_int;
endmodule
// removed package "rv_plic_reg_pkg"
module rv_plic_reg_top (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	reg2hw,
	hw2reg,
	intg_err_o,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:90387:15
	parameter signed [31:0] AW = 10;
	// Trace: design.sv:90389:3
	input clk_i;
	// Trace: design.sv:90390:3
	input rst_ni;
	// Trace: design.sv:90391:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:90392:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:90394:3
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_cc0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_ie0_mreg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_le_mreg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_msip0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio10_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio11_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio12_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio13_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio14_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio15_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio16_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio17_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio18_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio19_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio1_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio20_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio21_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio22_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio23_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio24_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio25_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio26_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio27_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio28_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio29_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio2_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio30_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio31_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio32_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio33_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio34_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio35_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio36_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio37_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio38_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio39_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio3_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio40_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio41_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio42_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio43_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio44_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio45_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio46_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio47_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio48_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio49_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio4_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio50_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio51_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio52_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio53_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio54_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio55_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio56_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio57_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio58_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio59_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio5_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio60_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio61_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio62_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio63_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio6_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio7_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio8_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio9_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_threshold0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_t
	output wire [331:0] reg2hw;
	// Trace: design.sv:90395:3
	// removed localparam type rv_plic_reg_pkg_rv_plic_hw2reg_cc0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_hw2reg_ip_mreg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_hw2reg_t
	input wire [133:0] hw2reg;
	// Trace: design.sv:90398:3
	output wire intg_err_o;
	// Trace: design.sv:90401:3
	input devmode_i;
	// Trace: design.sv:90404:3
	// removed import rv_plic_reg_pkg::*;
	// Trace: design.sv:90406:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:90407:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:90410:3
	wire reg_we;
	// Trace: design.sv:90411:3
	wire reg_re;
	// Trace: design.sv:90412:3
	wire [AW - 1:0] reg_addr;
	// Trace: design.sv:90413:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:90414:3
	wire [3:0] reg_be;
	// Trace: design.sv:90415:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:90416:3
	wire reg_error;
	// Trace: design.sv:90418:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:90420:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:90422:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_reg_h2d;
	// Trace: design.sv:90423:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_reg_d2h;
	// Trace: design.sv:90427:3
	assign intg_err_o = 1'b0;
	// Trace: design.sv:90429:3
	assign tl_reg_h2d = tl_i;
	// Trace: design.sv:90430:3
	assign tl_o = tl_reg_d2h;
	// Trace: design.sv:90433:3
	tlul_adapter_reg #(
		.RegAw(AW),
		.RegDw(DW),
		.EnableDataIntgGen(0)
	) u_reg_if(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_reg_h2d),
		.tl_o(tl_reg_d2h),
		.we_o(reg_we),
		.re_o(reg_re),
		.addr_o(reg_addr),
		.wdata_o(reg_wdata),
		.be_o(reg_be),
		.rdata_i(reg_rdata),
		.error_i(reg_error)
	);
	// Trace: design.sv:90453:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:90454:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:90460:3
	wire ip_0_p_0_qs;
	// Trace: design.sv:90461:3
	wire ip_0_p_1_qs;
	// Trace: design.sv:90462:3
	wire ip_0_p_2_qs;
	// Trace: design.sv:90463:3
	wire ip_0_p_3_qs;
	// Trace: design.sv:90464:3
	wire ip_0_p_4_qs;
	// Trace: design.sv:90465:3
	wire ip_0_p_5_qs;
	// Trace: design.sv:90466:3
	wire ip_0_p_6_qs;
	// Trace: design.sv:90467:3
	wire ip_0_p_7_qs;
	// Trace: design.sv:90468:3
	wire ip_0_p_8_qs;
	// Trace: design.sv:90469:3
	wire ip_0_p_9_qs;
	// Trace: design.sv:90470:3
	wire ip_0_p_10_qs;
	// Trace: design.sv:90471:3
	wire ip_0_p_11_qs;
	// Trace: design.sv:90472:3
	wire ip_0_p_12_qs;
	// Trace: design.sv:90473:3
	wire ip_0_p_13_qs;
	// Trace: design.sv:90474:3
	wire ip_0_p_14_qs;
	// Trace: design.sv:90475:3
	wire ip_0_p_15_qs;
	// Trace: design.sv:90476:3
	wire ip_0_p_16_qs;
	// Trace: design.sv:90477:3
	wire ip_0_p_17_qs;
	// Trace: design.sv:90478:3
	wire ip_0_p_18_qs;
	// Trace: design.sv:90479:3
	wire ip_0_p_19_qs;
	// Trace: design.sv:90480:3
	wire ip_0_p_20_qs;
	// Trace: design.sv:90481:3
	wire ip_0_p_21_qs;
	// Trace: design.sv:90482:3
	wire ip_0_p_22_qs;
	// Trace: design.sv:90483:3
	wire ip_0_p_23_qs;
	// Trace: design.sv:90484:3
	wire ip_0_p_24_qs;
	// Trace: design.sv:90485:3
	wire ip_0_p_25_qs;
	// Trace: design.sv:90486:3
	wire ip_0_p_26_qs;
	// Trace: design.sv:90487:3
	wire ip_0_p_27_qs;
	// Trace: design.sv:90488:3
	wire ip_0_p_28_qs;
	// Trace: design.sv:90489:3
	wire ip_0_p_29_qs;
	// Trace: design.sv:90490:3
	wire ip_0_p_30_qs;
	// Trace: design.sv:90491:3
	wire ip_0_p_31_qs;
	// Trace: design.sv:90492:3
	wire ip_1_p_32_qs;
	// Trace: design.sv:90493:3
	wire ip_1_p_33_qs;
	// Trace: design.sv:90494:3
	wire ip_1_p_34_qs;
	// Trace: design.sv:90495:3
	wire ip_1_p_35_qs;
	// Trace: design.sv:90496:3
	wire ip_1_p_36_qs;
	// Trace: design.sv:90497:3
	wire ip_1_p_37_qs;
	// Trace: design.sv:90498:3
	wire ip_1_p_38_qs;
	// Trace: design.sv:90499:3
	wire ip_1_p_39_qs;
	// Trace: design.sv:90500:3
	wire ip_1_p_40_qs;
	// Trace: design.sv:90501:3
	wire ip_1_p_41_qs;
	// Trace: design.sv:90502:3
	wire ip_1_p_42_qs;
	// Trace: design.sv:90503:3
	wire ip_1_p_43_qs;
	// Trace: design.sv:90504:3
	wire ip_1_p_44_qs;
	// Trace: design.sv:90505:3
	wire ip_1_p_45_qs;
	// Trace: design.sv:90506:3
	wire ip_1_p_46_qs;
	// Trace: design.sv:90507:3
	wire ip_1_p_47_qs;
	// Trace: design.sv:90508:3
	wire ip_1_p_48_qs;
	// Trace: design.sv:90509:3
	wire ip_1_p_49_qs;
	// Trace: design.sv:90510:3
	wire ip_1_p_50_qs;
	// Trace: design.sv:90511:3
	wire ip_1_p_51_qs;
	// Trace: design.sv:90512:3
	wire ip_1_p_52_qs;
	// Trace: design.sv:90513:3
	wire ip_1_p_53_qs;
	// Trace: design.sv:90514:3
	wire ip_1_p_54_qs;
	// Trace: design.sv:90515:3
	wire ip_1_p_55_qs;
	// Trace: design.sv:90516:3
	wire ip_1_p_56_qs;
	// Trace: design.sv:90517:3
	wire ip_1_p_57_qs;
	// Trace: design.sv:90518:3
	wire ip_1_p_58_qs;
	// Trace: design.sv:90519:3
	wire ip_1_p_59_qs;
	// Trace: design.sv:90520:3
	wire ip_1_p_60_qs;
	// Trace: design.sv:90521:3
	wire ip_1_p_61_qs;
	// Trace: design.sv:90522:3
	wire ip_1_p_62_qs;
	// Trace: design.sv:90523:3
	wire ip_1_p_63_qs;
	// Trace: design.sv:90524:3
	wire le_0_le_0_qs;
	// Trace: design.sv:90525:3
	wire le_0_le_0_wd;
	// Trace: design.sv:90526:3
	wire le_0_le_0_we;
	// Trace: design.sv:90527:3
	wire le_0_le_1_qs;
	// Trace: design.sv:90528:3
	wire le_0_le_1_wd;
	// Trace: design.sv:90529:3
	wire le_0_le_1_we;
	// Trace: design.sv:90530:3
	wire le_0_le_2_qs;
	// Trace: design.sv:90531:3
	wire le_0_le_2_wd;
	// Trace: design.sv:90532:3
	wire le_0_le_2_we;
	// Trace: design.sv:90533:3
	wire le_0_le_3_qs;
	// Trace: design.sv:90534:3
	wire le_0_le_3_wd;
	// Trace: design.sv:90535:3
	wire le_0_le_3_we;
	// Trace: design.sv:90536:3
	wire le_0_le_4_qs;
	// Trace: design.sv:90537:3
	wire le_0_le_4_wd;
	// Trace: design.sv:90538:3
	wire le_0_le_4_we;
	// Trace: design.sv:90539:3
	wire le_0_le_5_qs;
	// Trace: design.sv:90540:3
	wire le_0_le_5_wd;
	// Trace: design.sv:90541:3
	wire le_0_le_5_we;
	// Trace: design.sv:90542:3
	wire le_0_le_6_qs;
	// Trace: design.sv:90543:3
	wire le_0_le_6_wd;
	// Trace: design.sv:90544:3
	wire le_0_le_6_we;
	// Trace: design.sv:90545:3
	wire le_0_le_7_qs;
	// Trace: design.sv:90546:3
	wire le_0_le_7_wd;
	// Trace: design.sv:90547:3
	wire le_0_le_7_we;
	// Trace: design.sv:90548:3
	wire le_0_le_8_qs;
	// Trace: design.sv:90549:3
	wire le_0_le_8_wd;
	// Trace: design.sv:90550:3
	wire le_0_le_8_we;
	// Trace: design.sv:90551:3
	wire le_0_le_9_qs;
	// Trace: design.sv:90552:3
	wire le_0_le_9_wd;
	// Trace: design.sv:90553:3
	wire le_0_le_9_we;
	// Trace: design.sv:90554:3
	wire le_0_le_10_qs;
	// Trace: design.sv:90555:3
	wire le_0_le_10_wd;
	// Trace: design.sv:90556:3
	wire le_0_le_10_we;
	// Trace: design.sv:90557:3
	wire le_0_le_11_qs;
	// Trace: design.sv:90558:3
	wire le_0_le_11_wd;
	// Trace: design.sv:90559:3
	wire le_0_le_11_we;
	// Trace: design.sv:90560:3
	wire le_0_le_12_qs;
	// Trace: design.sv:90561:3
	wire le_0_le_12_wd;
	// Trace: design.sv:90562:3
	wire le_0_le_12_we;
	// Trace: design.sv:90563:3
	wire le_0_le_13_qs;
	// Trace: design.sv:90564:3
	wire le_0_le_13_wd;
	// Trace: design.sv:90565:3
	wire le_0_le_13_we;
	// Trace: design.sv:90566:3
	wire le_0_le_14_qs;
	// Trace: design.sv:90567:3
	wire le_0_le_14_wd;
	// Trace: design.sv:90568:3
	wire le_0_le_14_we;
	// Trace: design.sv:90569:3
	wire le_0_le_15_qs;
	// Trace: design.sv:90570:3
	wire le_0_le_15_wd;
	// Trace: design.sv:90571:3
	wire le_0_le_15_we;
	// Trace: design.sv:90572:3
	wire le_0_le_16_qs;
	// Trace: design.sv:90573:3
	wire le_0_le_16_wd;
	// Trace: design.sv:90574:3
	wire le_0_le_16_we;
	// Trace: design.sv:90575:3
	wire le_0_le_17_qs;
	// Trace: design.sv:90576:3
	wire le_0_le_17_wd;
	// Trace: design.sv:90577:3
	wire le_0_le_17_we;
	// Trace: design.sv:90578:3
	wire le_0_le_18_qs;
	// Trace: design.sv:90579:3
	wire le_0_le_18_wd;
	// Trace: design.sv:90580:3
	wire le_0_le_18_we;
	// Trace: design.sv:90581:3
	wire le_0_le_19_qs;
	// Trace: design.sv:90582:3
	wire le_0_le_19_wd;
	// Trace: design.sv:90583:3
	wire le_0_le_19_we;
	// Trace: design.sv:90584:3
	wire le_0_le_20_qs;
	// Trace: design.sv:90585:3
	wire le_0_le_20_wd;
	// Trace: design.sv:90586:3
	wire le_0_le_20_we;
	// Trace: design.sv:90587:3
	wire le_0_le_21_qs;
	// Trace: design.sv:90588:3
	wire le_0_le_21_wd;
	// Trace: design.sv:90589:3
	wire le_0_le_21_we;
	// Trace: design.sv:90590:3
	wire le_0_le_22_qs;
	// Trace: design.sv:90591:3
	wire le_0_le_22_wd;
	// Trace: design.sv:90592:3
	wire le_0_le_22_we;
	// Trace: design.sv:90593:3
	wire le_0_le_23_qs;
	// Trace: design.sv:90594:3
	wire le_0_le_23_wd;
	// Trace: design.sv:90595:3
	wire le_0_le_23_we;
	// Trace: design.sv:90596:3
	wire le_0_le_24_qs;
	// Trace: design.sv:90597:3
	wire le_0_le_24_wd;
	// Trace: design.sv:90598:3
	wire le_0_le_24_we;
	// Trace: design.sv:90599:3
	wire le_0_le_25_qs;
	// Trace: design.sv:90600:3
	wire le_0_le_25_wd;
	// Trace: design.sv:90601:3
	wire le_0_le_25_we;
	// Trace: design.sv:90602:3
	wire le_0_le_26_qs;
	// Trace: design.sv:90603:3
	wire le_0_le_26_wd;
	// Trace: design.sv:90604:3
	wire le_0_le_26_we;
	// Trace: design.sv:90605:3
	wire le_0_le_27_qs;
	// Trace: design.sv:90606:3
	wire le_0_le_27_wd;
	// Trace: design.sv:90607:3
	wire le_0_le_27_we;
	// Trace: design.sv:90608:3
	wire le_0_le_28_qs;
	// Trace: design.sv:90609:3
	wire le_0_le_28_wd;
	// Trace: design.sv:90610:3
	wire le_0_le_28_we;
	// Trace: design.sv:90611:3
	wire le_0_le_29_qs;
	// Trace: design.sv:90612:3
	wire le_0_le_29_wd;
	// Trace: design.sv:90613:3
	wire le_0_le_29_we;
	// Trace: design.sv:90614:3
	wire le_0_le_30_qs;
	// Trace: design.sv:90615:3
	wire le_0_le_30_wd;
	// Trace: design.sv:90616:3
	wire le_0_le_30_we;
	// Trace: design.sv:90617:3
	wire le_0_le_31_qs;
	// Trace: design.sv:90618:3
	wire le_0_le_31_wd;
	// Trace: design.sv:90619:3
	wire le_0_le_31_we;
	// Trace: design.sv:90620:3
	wire le_1_le_32_qs;
	// Trace: design.sv:90621:3
	wire le_1_le_32_wd;
	// Trace: design.sv:90622:3
	wire le_1_le_32_we;
	// Trace: design.sv:90623:3
	wire le_1_le_33_qs;
	// Trace: design.sv:90624:3
	wire le_1_le_33_wd;
	// Trace: design.sv:90625:3
	wire le_1_le_33_we;
	// Trace: design.sv:90626:3
	wire le_1_le_34_qs;
	// Trace: design.sv:90627:3
	wire le_1_le_34_wd;
	// Trace: design.sv:90628:3
	wire le_1_le_34_we;
	// Trace: design.sv:90629:3
	wire le_1_le_35_qs;
	// Trace: design.sv:90630:3
	wire le_1_le_35_wd;
	// Trace: design.sv:90631:3
	wire le_1_le_35_we;
	// Trace: design.sv:90632:3
	wire le_1_le_36_qs;
	// Trace: design.sv:90633:3
	wire le_1_le_36_wd;
	// Trace: design.sv:90634:3
	wire le_1_le_36_we;
	// Trace: design.sv:90635:3
	wire le_1_le_37_qs;
	// Trace: design.sv:90636:3
	wire le_1_le_37_wd;
	// Trace: design.sv:90637:3
	wire le_1_le_37_we;
	// Trace: design.sv:90638:3
	wire le_1_le_38_qs;
	// Trace: design.sv:90639:3
	wire le_1_le_38_wd;
	// Trace: design.sv:90640:3
	wire le_1_le_38_we;
	// Trace: design.sv:90641:3
	wire le_1_le_39_qs;
	// Trace: design.sv:90642:3
	wire le_1_le_39_wd;
	// Trace: design.sv:90643:3
	wire le_1_le_39_we;
	// Trace: design.sv:90644:3
	wire le_1_le_40_qs;
	// Trace: design.sv:90645:3
	wire le_1_le_40_wd;
	// Trace: design.sv:90646:3
	wire le_1_le_40_we;
	// Trace: design.sv:90647:3
	wire le_1_le_41_qs;
	// Trace: design.sv:90648:3
	wire le_1_le_41_wd;
	// Trace: design.sv:90649:3
	wire le_1_le_41_we;
	// Trace: design.sv:90650:3
	wire le_1_le_42_qs;
	// Trace: design.sv:90651:3
	wire le_1_le_42_wd;
	// Trace: design.sv:90652:3
	wire le_1_le_42_we;
	// Trace: design.sv:90653:3
	wire le_1_le_43_qs;
	// Trace: design.sv:90654:3
	wire le_1_le_43_wd;
	// Trace: design.sv:90655:3
	wire le_1_le_43_we;
	// Trace: design.sv:90656:3
	wire le_1_le_44_qs;
	// Trace: design.sv:90657:3
	wire le_1_le_44_wd;
	// Trace: design.sv:90658:3
	wire le_1_le_44_we;
	// Trace: design.sv:90659:3
	wire le_1_le_45_qs;
	// Trace: design.sv:90660:3
	wire le_1_le_45_wd;
	// Trace: design.sv:90661:3
	wire le_1_le_45_we;
	// Trace: design.sv:90662:3
	wire le_1_le_46_qs;
	// Trace: design.sv:90663:3
	wire le_1_le_46_wd;
	// Trace: design.sv:90664:3
	wire le_1_le_46_we;
	// Trace: design.sv:90665:3
	wire le_1_le_47_qs;
	// Trace: design.sv:90666:3
	wire le_1_le_47_wd;
	// Trace: design.sv:90667:3
	wire le_1_le_47_we;
	// Trace: design.sv:90668:3
	wire le_1_le_48_qs;
	// Trace: design.sv:90669:3
	wire le_1_le_48_wd;
	// Trace: design.sv:90670:3
	wire le_1_le_48_we;
	// Trace: design.sv:90671:3
	wire le_1_le_49_qs;
	// Trace: design.sv:90672:3
	wire le_1_le_49_wd;
	// Trace: design.sv:90673:3
	wire le_1_le_49_we;
	// Trace: design.sv:90674:3
	wire le_1_le_50_qs;
	// Trace: design.sv:90675:3
	wire le_1_le_50_wd;
	// Trace: design.sv:90676:3
	wire le_1_le_50_we;
	// Trace: design.sv:90677:3
	wire le_1_le_51_qs;
	// Trace: design.sv:90678:3
	wire le_1_le_51_wd;
	// Trace: design.sv:90679:3
	wire le_1_le_51_we;
	// Trace: design.sv:90680:3
	wire le_1_le_52_qs;
	// Trace: design.sv:90681:3
	wire le_1_le_52_wd;
	// Trace: design.sv:90682:3
	wire le_1_le_52_we;
	// Trace: design.sv:90683:3
	wire le_1_le_53_qs;
	// Trace: design.sv:90684:3
	wire le_1_le_53_wd;
	// Trace: design.sv:90685:3
	wire le_1_le_53_we;
	// Trace: design.sv:90686:3
	wire le_1_le_54_qs;
	// Trace: design.sv:90687:3
	wire le_1_le_54_wd;
	// Trace: design.sv:90688:3
	wire le_1_le_54_we;
	// Trace: design.sv:90689:3
	wire le_1_le_55_qs;
	// Trace: design.sv:90690:3
	wire le_1_le_55_wd;
	// Trace: design.sv:90691:3
	wire le_1_le_55_we;
	// Trace: design.sv:90692:3
	wire le_1_le_56_qs;
	// Trace: design.sv:90693:3
	wire le_1_le_56_wd;
	// Trace: design.sv:90694:3
	wire le_1_le_56_we;
	// Trace: design.sv:90695:3
	wire le_1_le_57_qs;
	// Trace: design.sv:90696:3
	wire le_1_le_57_wd;
	// Trace: design.sv:90697:3
	wire le_1_le_57_we;
	// Trace: design.sv:90698:3
	wire le_1_le_58_qs;
	// Trace: design.sv:90699:3
	wire le_1_le_58_wd;
	// Trace: design.sv:90700:3
	wire le_1_le_58_we;
	// Trace: design.sv:90701:3
	wire le_1_le_59_qs;
	// Trace: design.sv:90702:3
	wire le_1_le_59_wd;
	// Trace: design.sv:90703:3
	wire le_1_le_59_we;
	// Trace: design.sv:90704:3
	wire le_1_le_60_qs;
	// Trace: design.sv:90705:3
	wire le_1_le_60_wd;
	// Trace: design.sv:90706:3
	wire le_1_le_60_we;
	// Trace: design.sv:90707:3
	wire le_1_le_61_qs;
	// Trace: design.sv:90708:3
	wire le_1_le_61_wd;
	// Trace: design.sv:90709:3
	wire le_1_le_61_we;
	// Trace: design.sv:90710:3
	wire le_1_le_62_qs;
	// Trace: design.sv:90711:3
	wire le_1_le_62_wd;
	// Trace: design.sv:90712:3
	wire le_1_le_62_we;
	// Trace: design.sv:90713:3
	wire le_1_le_63_qs;
	// Trace: design.sv:90714:3
	wire le_1_le_63_wd;
	// Trace: design.sv:90715:3
	wire le_1_le_63_we;
	// Trace: design.sv:90716:3
	wire [2:0] prio0_qs;
	// Trace: design.sv:90717:3
	wire [2:0] prio0_wd;
	// Trace: design.sv:90718:3
	wire prio0_we;
	// Trace: design.sv:90719:3
	wire [2:0] prio1_qs;
	// Trace: design.sv:90720:3
	wire [2:0] prio1_wd;
	// Trace: design.sv:90721:3
	wire prio1_we;
	// Trace: design.sv:90722:3
	wire [2:0] prio2_qs;
	// Trace: design.sv:90723:3
	wire [2:0] prio2_wd;
	// Trace: design.sv:90724:3
	wire prio2_we;
	// Trace: design.sv:90725:3
	wire [2:0] prio3_qs;
	// Trace: design.sv:90726:3
	wire [2:0] prio3_wd;
	// Trace: design.sv:90727:3
	wire prio3_we;
	// Trace: design.sv:90728:3
	wire [2:0] prio4_qs;
	// Trace: design.sv:90729:3
	wire [2:0] prio4_wd;
	// Trace: design.sv:90730:3
	wire prio4_we;
	// Trace: design.sv:90731:3
	wire [2:0] prio5_qs;
	// Trace: design.sv:90732:3
	wire [2:0] prio5_wd;
	// Trace: design.sv:90733:3
	wire prio5_we;
	// Trace: design.sv:90734:3
	wire [2:0] prio6_qs;
	// Trace: design.sv:90735:3
	wire [2:0] prio6_wd;
	// Trace: design.sv:90736:3
	wire prio6_we;
	// Trace: design.sv:90737:3
	wire [2:0] prio7_qs;
	// Trace: design.sv:90738:3
	wire [2:0] prio7_wd;
	// Trace: design.sv:90739:3
	wire prio7_we;
	// Trace: design.sv:90740:3
	wire [2:0] prio8_qs;
	// Trace: design.sv:90741:3
	wire [2:0] prio8_wd;
	// Trace: design.sv:90742:3
	wire prio8_we;
	// Trace: design.sv:90743:3
	wire [2:0] prio9_qs;
	// Trace: design.sv:90744:3
	wire [2:0] prio9_wd;
	// Trace: design.sv:90745:3
	wire prio9_we;
	// Trace: design.sv:90746:3
	wire [2:0] prio10_qs;
	// Trace: design.sv:90747:3
	wire [2:0] prio10_wd;
	// Trace: design.sv:90748:3
	wire prio10_we;
	// Trace: design.sv:90749:3
	wire [2:0] prio11_qs;
	// Trace: design.sv:90750:3
	wire [2:0] prio11_wd;
	// Trace: design.sv:90751:3
	wire prio11_we;
	// Trace: design.sv:90752:3
	wire [2:0] prio12_qs;
	// Trace: design.sv:90753:3
	wire [2:0] prio12_wd;
	// Trace: design.sv:90754:3
	wire prio12_we;
	// Trace: design.sv:90755:3
	wire [2:0] prio13_qs;
	// Trace: design.sv:90756:3
	wire [2:0] prio13_wd;
	// Trace: design.sv:90757:3
	wire prio13_we;
	// Trace: design.sv:90758:3
	wire [2:0] prio14_qs;
	// Trace: design.sv:90759:3
	wire [2:0] prio14_wd;
	// Trace: design.sv:90760:3
	wire prio14_we;
	// Trace: design.sv:90761:3
	wire [2:0] prio15_qs;
	// Trace: design.sv:90762:3
	wire [2:0] prio15_wd;
	// Trace: design.sv:90763:3
	wire prio15_we;
	// Trace: design.sv:90764:3
	wire [2:0] prio16_qs;
	// Trace: design.sv:90765:3
	wire [2:0] prio16_wd;
	// Trace: design.sv:90766:3
	wire prio16_we;
	// Trace: design.sv:90767:3
	wire [2:0] prio17_qs;
	// Trace: design.sv:90768:3
	wire [2:0] prio17_wd;
	// Trace: design.sv:90769:3
	wire prio17_we;
	// Trace: design.sv:90770:3
	wire [2:0] prio18_qs;
	// Trace: design.sv:90771:3
	wire [2:0] prio18_wd;
	// Trace: design.sv:90772:3
	wire prio18_we;
	// Trace: design.sv:90773:3
	wire [2:0] prio19_qs;
	// Trace: design.sv:90774:3
	wire [2:0] prio19_wd;
	// Trace: design.sv:90775:3
	wire prio19_we;
	// Trace: design.sv:90776:3
	wire [2:0] prio20_qs;
	// Trace: design.sv:90777:3
	wire [2:0] prio20_wd;
	// Trace: design.sv:90778:3
	wire prio20_we;
	// Trace: design.sv:90779:3
	wire [2:0] prio21_qs;
	// Trace: design.sv:90780:3
	wire [2:0] prio21_wd;
	// Trace: design.sv:90781:3
	wire prio21_we;
	// Trace: design.sv:90782:3
	wire [2:0] prio22_qs;
	// Trace: design.sv:90783:3
	wire [2:0] prio22_wd;
	// Trace: design.sv:90784:3
	wire prio22_we;
	// Trace: design.sv:90785:3
	wire [2:0] prio23_qs;
	// Trace: design.sv:90786:3
	wire [2:0] prio23_wd;
	// Trace: design.sv:90787:3
	wire prio23_we;
	// Trace: design.sv:90788:3
	wire [2:0] prio24_qs;
	// Trace: design.sv:90789:3
	wire [2:0] prio24_wd;
	// Trace: design.sv:90790:3
	wire prio24_we;
	// Trace: design.sv:90791:3
	wire [2:0] prio25_qs;
	// Trace: design.sv:90792:3
	wire [2:0] prio25_wd;
	// Trace: design.sv:90793:3
	wire prio25_we;
	// Trace: design.sv:90794:3
	wire [2:0] prio26_qs;
	// Trace: design.sv:90795:3
	wire [2:0] prio26_wd;
	// Trace: design.sv:90796:3
	wire prio26_we;
	// Trace: design.sv:90797:3
	wire [2:0] prio27_qs;
	// Trace: design.sv:90798:3
	wire [2:0] prio27_wd;
	// Trace: design.sv:90799:3
	wire prio27_we;
	// Trace: design.sv:90800:3
	wire [2:0] prio28_qs;
	// Trace: design.sv:90801:3
	wire [2:0] prio28_wd;
	// Trace: design.sv:90802:3
	wire prio28_we;
	// Trace: design.sv:90803:3
	wire [2:0] prio29_qs;
	// Trace: design.sv:90804:3
	wire [2:0] prio29_wd;
	// Trace: design.sv:90805:3
	wire prio29_we;
	// Trace: design.sv:90806:3
	wire [2:0] prio30_qs;
	// Trace: design.sv:90807:3
	wire [2:0] prio30_wd;
	// Trace: design.sv:90808:3
	wire prio30_we;
	// Trace: design.sv:90809:3
	wire [2:0] prio31_qs;
	// Trace: design.sv:90810:3
	wire [2:0] prio31_wd;
	// Trace: design.sv:90811:3
	wire prio31_we;
	// Trace: design.sv:90812:3
	wire [2:0] prio32_qs;
	// Trace: design.sv:90813:3
	wire [2:0] prio32_wd;
	// Trace: design.sv:90814:3
	wire prio32_we;
	// Trace: design.sv:90815:3
	wire [2:0] prio33_qs;
	// Trace: design.sv:90816:3
	wire [2:0] prio33_wd;
	// Trace: design.sv:90817:3
	wire prio33_we;
	// Trace: design.sv:90818:3
	wire [2:0] prio34_qs;
	// Trace: design.sv:90819:3
	wire [2:0] prio34_wd;
	// Trace: design.sv:90820:3
	wire prio34_we;
	// Trace: design.sv:90821:3
	wire [2:0] prio35_qs;
	// Trace: design.sv:90822:3
	wire [2:0] prio35_wd;
	// Trace: design.sv:90823:3
	wire prio35_we;
	// Trace: design.sv:90824:3
	wire [2:0] prio36_qs;
	// Trace: design.sv:90825:3
	wire [2:0] prio36_wd;
	// Trace: design.sv:90826:3
	wire prio36_we;
	// Trace: design.sv:90827:3
	wire [2:0] prio37_qs;
	// Trace: design.sv:90828:3
	wire [2:0] prio37_wd;
	// Trace: design.sv:90829:3
	wire prio37_we;
	// Trace: design.sv:90830:3
	wire [2:0] prio38_qs;
	// Trace: design.sv:90831:3
	wire [2:0] prio38_wd;
	// Trace: design.sv:90832:3
	wire prio38_we;
	// Trace: design.sv:90833:3
	wire [2:0] prio39_qs;
	// Trace: design.sv:90834:3
	wire [2:0] prio39_wd;
	// Trace: design.sv:90835:3
	wire prio39_we;
	// Trace: design.sv:90836:3
	wire [2:0] prio40_qs;
	// Trace: design.sv:90837:3
	wire [2:0] prio40_wd;
	// Trace: design.sv:90838:3
	wire prio40_we;
	// Trace: design.sv:90839:3
	wire [2:0] prio41_qs;
	// Trace: design.sv:90840:3
	wire [2:0] prio41_wd;
	// Trace: design.sv:90841:3
	wire prio41_we;
	// Trace: design.sv:90842:3
	wire [2:0] prio42_qs;
	// Trace: design.sv:90843:3
	wire [2:0] prio42_wd;
	// Trace: design.sv:90844:3
	wire prio42_we;
	// Trace: design.sv:90845:3
	wire [2:0] prio43_qs;
	// Trace: design.sv:90846:3
	wire [2:0] prio43_wd;
	// Trace: design.sv:90847:3
	wire prio43_we;
	// Trace: design.sv:90848:3
	wire [2:0] prio44_qs;
	// Trace: design.sv:90849:3
	wire [2:0] prio44_wd;
	// Trace: design.sv:90850:3
	wire prio44_we;
	// Trace: design.sv:90851:3
	wire [2:0] prio45_qs;
	// Trace: design.sv:90852:3
	wire [2:0] prio45_wd;
	// Trace: design.sv:90853:3
	wire prio45_we;
	// Trace: design.sv:90854:3
	wire [2:0] prio46_qs;
	// Trace: design.sv:90855:3
	wire [2:0] prio46_wd;
	// Trace: design.sv:90856:3
	wire prio46_we;
	// Trace: design.sv:90857:3
	wire [2:0] prio47_qs;
	// Trace: design.sv:90858:3
	wire [2:0] prio47_wd;
	// Trace: design.sv:90859:3
	wire prio47_we;
	// Trace: design.sv:90860:3
	wire [2:0] prio48_qs;
	// Trace: design.sv:90861:3
	wire [2:0] prio48_wd;
	// Trace: design.sv:90862:3
	wire prio48_we;
	// Trace: design.sv:90863:3
	wire [2:0] prio49_qs;
	// Trace: design.sv:90864:3
	wire [2:0] prio49_wd;
	// Trace: design.sv:90865:3
	wire prio49_we;
	// Trace: design.sv:90866:3
	wire [2:0] prio50_qs;
	// Trace: design.sv:90867:3
	wire [2:0] prio50_wd;
	// Trace: design.sv:90868:3
	wire prio50_we;
	// Trace: design.sv:90869:3
	wire [2:0] prio51_qs;
	// Trace: design.sv:90870:3
	wire [2:0] prio51_wd;
	// Trace: design.sv:90871:3
	wire prio51_we;
	// Trace: design.sv:90872:3
	wire [2:0] prio52_qs;
	// Trace: design.sv:90873:3
	wire [2:0] prio52_wd;
	// Trace: design.sv:90874:3
	wire prio52_we;
	// Trace: design.sv:90875:3
	wire [2:0] prio53_qs;
	// Trace: design.sv:90876:3
	wire [2:0] prio53_wd;
	// Trace: design.sv:90877:3
	wire prio53_we;
	// Trace: design.sv:90878:3
	wire [2:0] prio54_qs;
	// Trace: design.sv:90879:3
	wire [2:0] prio54_wd;
	// Trace: design.sv:90880:3
	wire prio54_we;
	// Trace: design.sv:90881:3
	wire [2:0] prio55_qs;
	// Trace: design.sv:90882:3
	wire [2:0] prio55_wd;
	// Trace: design.sv:90883:3
	wire prio55_we;
	// Trace: design.sv:90884:3
	wire [2:0] prio56_qs;
	// Trace: design.sv:90885:3
	wire [2:0] prio56_wd;
	// Trace: design.sv:90886:3
	wire prio56_we;
	// Trace: design.sv:90887:3
	wire [2:0] prio57_qs;
	// Trace: design.sv:90888:3
	wire [2:0] prio57_wd;
	// Trace: design.sv:90889:3
	wire prio57_we;
	// Trace: design.sv:90890:3
	wire [2:0] prio58_qs;
	// Trace: design.sv:90891:3
	wire [2:0] prio58_wd;
	// Trace: design.sv:90892:3
	wire prio58_we;
	// Trace: design.sv:90893:3
	wire [2:0] prio59_qs;
	// Trace: design.sv:90894:3
	wire [2:0] prio59_wd;
	// Trace: design.sv:90895:3
	wire prio59_we;
	// Trace: design.sv:90896:3
	wire [2:0] prio60_qs;
	// Trace: design.sv:90897:3
	wire [2:0] prio60_wd;
	// Trace: design.sv:90898:3
	wire prio60_we;
	// Trace: design.sv:90899:3
	wire [2:0] prio61_qs;
	// Trace: design.sv:90900:3
	wire [2:0] prio61_wd;
	// Trace: design.sv:90901:3
	wire prio61_we;
	// Trace: design.sv:90902:3
	wire [2:0] prio62_qs;
	// Trace: design.sv:90903:3
	wire [2:0] prio62_wd;
	// Trace: design.sv:90904:3
	wire prio62_we;
	// Trace: design.sv:90905:3
	wire [2:0] prio63_qs;
	// Trace: design.sv:90906:3
	wire [2:0] prio63_wd;
	// Trace: design.sv:90907:3
	wire prio63_we;
	// Trace: design.sv:90908:3
	wire ie0_0_e_0_qs;
	// Trace: design.sv:90909:3
	wire ie0_0_e_0_wd;
	// Trace: design.sv:90910:3
	wire ie0_0_e_0_we;
	// Trace: design.sv:90911:3
	wire ie0_0_e_1_qs;
	// Trace: design.sv:90912:3
	wire ie0_0_e_1_wd;
	// Trace: design.sv:90913:3
	wire ie0_0_e_1_we;
	// Trace: design.sv:90914:3
	wire ie0_0_e_2_qs;
	// Trace: design.sv:90915:3
	wire ie0_0_e_2_wd;
	// Trace: design.sv:90916:3
	wire ie0_0_e_2_we;
	// Trace: design.sv:90917:3
	wire ie0_0_e_3_qs;
	// Trace: design.sv:90918:3
	wire ie0_0_e_3_wd;
	// Trace: design.sv:90919:3
	wire ie0_0_e_3_we;
	// Trace: design.sv:90920:3
	wire ie0_0_e_4_qs;
	// Trace: design.sv:90921:3
	wire ie0_0_e_4_wd;
	// Trace: design.sv:90922:3
	wire ie0_0_e_4_we;
	// Trace: design.sv:90923:3
	wire ie0_0_e_5_qs;
	// Trace: design.sv:90924:3
	wire ie0_0_e_5_wd;
	// Trace: design.sv:90925:3
	wire ie0_0_e_5_we;
	// Trace: design.sv:90926:3
	wire ie0_0_e_6_qs;
	// Trace: design.sv:90927:3
	wire ie0_0_e_6_wd;
	// Trace: design.sv:90928:3
	wire ie0_0_e_6_we;
	// Trace: design.sv:90929:3
	wire ie0_0_e_7_qs;
	// Trace: design.sv:90930:3
	wire ie0_0_e_7_wd;
	// Trace: design.sv:90931:3
	wire ie0_0_e_7_we;
	// Trace: design.sv:90932:3
	wire ie0_0_e_8_qs;
	// Trace: design.sv:90933:3
	wire ie0_0_e_8_wd;
	// Trace: design.sv:90934:3
	wire ie0_0_e_8_we;
	// Trace: design.sv:90935:3
	wire ie0_0_e_9_qs;
	// Trace: design.sv:90936:3
	wire ie0_0_e_9_wd;
	// Trace: design.sv:90937:3
	wire ie0_0_e_9_we;
	// Trace: design.sv:90938:3
	wire ie0_0_e_10_qs;
	// Trace: design.sv:90939:3
	wire ie0_0_e_10_wd;
	// Trace: design.sv:90940:3
	wire ie0_0_e_10_we;
	// Trace: design.sv:90941:3
	wire ie0_0_e_11_qs;
	// Trace: design.sv:90942:3
	wire ie0_0_e_11_wd;
	// Trace: design.sv:90943:3
	wire ie0_0_e_11_we;
	// Trace: design.sv:90944:3
	wire ie0_0_e_12_qs;
	// Trace: design.sv:90945:3
	wire ie0_0_e_12_wd;
	// Trace: design.sv:90946:3
	wire ie0_0_e_12_we;
	// Trace: design.sv:90947:3
	wire ie0_0_e_13_qs;
	// Trace: design.sv:90948:3
	wire ie0_0_e_13_wd;
	// Trace: design.sv:90949:3
	wire ie0_0_e_13_we;
	// Trace: design.sv:90950:3
	wire ie0_0_e_14_qs;
	// Trace: design.sv:90951:3
	wire ie0_0_e_14_wd;
	// Trace: design.sv:90952:3
	wire ie0_0_e_14_we;
	// Trace: design.sv:90953:3
	wire ie0_0_e_15_qs;
	// Trace: design.sv:90954:3
	wire ie0_0_e_15_wd;
	// Trace: design.sv:90955:3
	wire ie0_0_e_15_we;
	// Trace: design.sv:90956:3
	wire ie0_0_e_16_qs;
	// Trace: design.sv:90957:3
	wire ie0_0_e_16_wd;
	// Trace: design.sv:90958:3
	wire ie0_0_e_16_we;
	// Trace: design.sv:90959:3
	wire ie0_0_e_17_qs;
	// Trace: design.sv:90960:3
	wire ie0_0_e_17_wd;
	// Trace: design.sv:90961:3
	wire ie0_0_e_17_we;
	// Trace: design.sv:90962:3
	wire ie0_0_e_18_qs;
	// Trace: design.sv:90963:3
	wire ie0_0_e_18_wd;
	// Trace: design.sv:90964:3
	wire ie0_0_e_18_we;
	// Trace: design.sv:90965:3
	wire ie0_0_e_19_qs;
	// Trace: design.sv:90966:3
	wire ie0_0_e_19_wd;
	// Trace: design.sv:90967:3
	wire ie0_0_e_19_we;
	// Trace: design.sv:90968:3
	wire ie0_0_e_20_qs;
	// Trace: design.sv:90969:3
	wire ie0_0_e_20_wd;
	// Trace: design.sv:90970:3
	wire ie0_0_e_20_we;
	// Trace: design.sv:90971:3
	wire ie0_0_e_21_qs;
	// Trace: design.sv:90972:3
	wire ie0_0_e_21_wd;
	// Trace: design.sv:90973:3
	wire ie0_0_e_21_we;
	// Trace: design.sv:90974:3
	wire ie0_0_e_22_qs;
	// Trace: design.sv:90975:3
	wire ie0_0_e_22_wd;
	// Trace: design.sv:90976:3
	wire ie0_0_e_22_we;
	// Trace: design.sv:90977:3
	wire ie0_0_e_23_qs;
	// Trace: design.sv:90978:3
	wire ie0_0_e_23_wd;
	// Trace: design.sv:90979:3
	wire ie0_0_e_23_we;
	// Trace: design.sv:90980:3
	wire ie0_0_e_24_qs;
	// Trace: design.sv:90981:3
	wire ie0_0_e_24_wd;
	// Trace: design.sv:90982:3
	wire ie0_0_e_24_we;
	// Trace: design.sv:90983:3
	wire ie0_0_e_25_qs;
	// Trace: design.sv:90984:3
	wire ie0_0_e_25_wd;
	// Trace: design.sv:90985:3
	wire ie0_0_e_25_we;
	// Trace: design.sv:90986:3
	wire ie0_0_e_26_qs;
	// Trace: design.sv:90987:3
	wire ie0_0_e_26_wd;
	// Trace: design.sv:90988:3
	wire ie0_0_e_26_we;
	// Trace: design.sv:90989:3
	wire ie0_0_e_27_qs;
	// Trace: design.sv:90990:3
	wire ie0_0_e_27_wd;
	// Trace: design.sv:90991:3
	wire ie0_0_e_27_we;
	// Trace: design.sv:90992:3
	wire ie0_0_e_28_qs;
	// Trace: design.sv:90993:3
	wire ie0_0_e_28_wd;
	// Trace: design.sv:90994:3
	wire ie0_0_e_28_we;
	// Trace: design.sv:90995:3
	wire ie0_0_e_29_qs;
	// Trace: design.sv:90996:3
	wire ie0_0_e_29_wd;
	// Trace: design.sv:90997:3
	wire ie0_0_e_29_we;
	// Trace: design.sv:90998:3
	wire ie0_0_e_30_qs;
	// Trace: design.sv:90999:3
	wire ie0_0_e_30_wd;
	// Trace: design.sv:91000:3
	wire ie0_0_e_30_we;
	// Trace: design.sv:91001:3
	wire ie0_0_e_31_qs;
	// Trace: design.sv:91002:3
	wire ie0_0_e_31_wd;
	// Trace: design.sv:91003:3
	wire ie0_0_e_31_we;
	// Trace: design.sv:91004:3
	wire ie0_1_e_32_qs;
	// Trace: design.sv:91005:3
	wire ie0_1_e_32_wd;
	// Trace: design.sv:91006:3
	wire ie0_1_e_32_we;
	// Trace: design.sv:91007:3
	wire ie0_1_e_33_qs;
	// Trace: design.sv:91008:3
	wire ie0_1_e_33_wd;
	// Trace: design.sv:91009:3
	wire ie0_1_e_33_we;
	// Trace: design.sv:91010:3
	wire ie0_1_e_34_qs;
	// Trace: design.sv:91011:3
	wire ie0_1_e_34_wd;
	// Trace: design.sv:91012:3
	wire ie0_1_e_34_we;
	// Trace: design.sv:91013:3
	wire ie0_1_e_35_qs;
	// Trace: design.sv:91014:3
	wire ie0_1_e_35_wd;
	// Trace: design.sv:91015:3
	wire ie0_1_e_35_we;
	// Trace: design.sv:91016:3
	wire ie0_1_e_36_qs;
	// Trace: design.sv:91017:3
	wire ie0_1_e_36_wd;
	// Trace: design.sv:91018:3
	wire ie0_1_e_36_we;
	// Trace: design.sv:91019:3
	wire ie0_1_e_37_qs;
	// Trace: design.sv:91020:3
	wire ie0_1_e_37_wd;
	// Trace: design.sv:91021:3
	wire ie0_1_e_37_we;
	// Trace: design.sv:91022:3
	wire ie0_1_e_38_qs;
	// Trace: design.sv:91023:3
	wire ie0_1_e_38_wd;
	// Trace: design.sv:91024:3
	wire ie0_1_e_38_we;
	// Trace: design.sv:91025:3
	wire ie0_1_e_39_qs;
	// Trace: design.sv:91026:3
	wire ie0_1_e_39_wd;
	// Trace: design.sv:91027:3
	wire ie0_1_e_39_we;
	// Trace: design.sv:91028:3
	wire ie0_1_e_40_qs;
	// Trace: design.sv:91029:3
	wire ie0_1_e_40_wd;
	// Trace: design.sv:91030:3
	wire ie0_1_e_40_we;
	// Trace: design.sv:91031:3
	wire ie0_1_e_41_qs;
	// Trace: design.sv:91032:3
	wire ie0_1_e_41_wd;
	// Trace: design.sv:91033:3
	wire ie0_1_e_41_we;
	// Trace: design.sv:91034:3
	wire ie0_1_e_42_qs;
	// Trace: design.sv:91035:3
	wire ie0_1_e_42_wd;
	// Trace: design.sv:91036:3
	wire ie0_1_e_42_we;
	// Trace: design.sv:91037:3
	wire ie0_1_e_43_qs;
	// Trace: design.sv:91038:3
	wire ie0_1_e_43_wd;
	// Trace: design.sv:91039:3
	wire ie0_1_e_43_we;
	// Trace: design.sv:91040:3
	wire ie0_1_e_44_qs;
	// Trace: design.sv:91041:3
	wire ie0_1_e_44_wd;
	// Trace: design.sv:91042:3
	wire ie0_1_e_44_we;
	// Trace: design.sv:91043:3
	wire ie0_1_e_45_qs;
	// Trace: design.sv:91044:3
	wire ie0_1_e_45_wd;
	// Trace: design.sv:91045:3
	wire ie0_1_e_45_we;
	// Trace: design.sv:91046:3
	wire ie0_1_e_46_qs;
	// Trace: design.sv:91047:3
	wire ie0_1_e_46_wd;
	// Trace: design.sv:91048:3
	wire ie0_1_e_46_we;
	// Trace: design.sv:91049:3
	wire ie0_1_e_47_qs;
	// Trace: design.sv:91050:3
	wire ie0_1_e_47_wd;
	// Trace: design.sv:91051:3
	wire ie0_1_e_47_we;
	// Trace: design.sv:91052:3
	wire ie0_1_e_48_qs;
	// Trace: design.sv:91053:3
	wire ie0_1_e_48_wd;
	// Trace: design.sv:91054:3
	wire ie0_1_e_48_we;
	// Trace: design.sv:91055:3
	wire ie0_1_e_49_qs;
	// Trace: design.sv:91056:3
	wire ie0_1_e_49_wd;
	// Trace: design.sv:91057:3
	wire ie0_1_e_49_we;
	// Trace: design.sv:91058:3
	wire ie0_1_e_50_qs;
	// Trace: design.sv:91059:3
	wire ie0_1_e_50_wd;
	// Trace: design.sv:91060:3
	wire ie0_1_e_50_we;
	// Trace: design.sv:91061:3
	wire ie0_1_e_51_qs;
	// Trace: design.sv:91062:3
	wire ie0_1_e_51_wd;
	// Trace: design.sv:91063:3
	wire ie0_1_e_51_we;
	// Trace: design.sv:91064:3
	wire ie0_1_e_52_qs;
	// Trace: design.sv:91065:3
	wire ie0_1_e_52_wd;
	// Trace: design.sv:91066:3
	wire ie0_1_e_52_we;
	// Trace: design.sv:91067:3
	wire ie0_1_e_53_qs;
	// Trace: design.sv:91068:3
	wire ie0_1_e_53_wd;
	// Trace: design.sv:91069:3
	wire ie0_1_e_53_we;
	// Trace: design.sv:91070:3
	wire ie0_1_e_54_qs;
	// Trace: design.sv:91071:3
	wire ie0_1_e_54_wd;
	// Trace: design.sv:91072:3
	wire ie0_1_e_54_we;
	// Trace: design.sv:91073:3
	wire ie0_1_e_55_qs;
	// Trace: design.sv:91074:3
	wire ie0_1_e_55_wd;
	// Trace: design.sv:91075:3
	wire ie0_1_e_55_we;
	// Trace: design.sv:91076:3
	wire ie0_1_e_56_qs;
	// Trace: design.sv:91077:3
	wire ie0_1_e_56_wd;
	// Trace: design.sv:91078:3
	wire ie0_1_e_56_we;
	// Trace: design.sv:91079:3
	wire ie0_1_e_57_qs;
	// Trace: design.sv:91080:3
	wire ie0_1_e_57_wd;
	// Trace: design.sv:91081:3
	wire ie0_1_e_57_we;
	// Trace: design.sv:91082:3
	wire ie0_1_e_58_qs;
	// Trace: design.sv:91083:3
	wire ie0_1_e_58_wd;
	// Trace: design.sv:91084:3
	wire ie0_1_e_58_we;
	// Trace: design.sv:91085:3
	wire ie0_1_e_59_qs;
	// Trace: design.sv:91086:3
	wire ie0_1_e_59_wd;
	// Trace: design.sv:91087:3
	wire ie0_1_e_59_we;
	// Trace: design.sv:91088:3
	wire ie0_1_e_60_qs;
	// Trace: design.sv:91089:3
	wire ie0_1_e_60_wd;
	// Trace: design.sv:91090:3
	wire ie0_1_e_60_we;
	// Trace: design.sv:91091:3
	wire ie0_1_e_61_qs;
	// Trace: design.sv:91092:3
	wire ie0_1_e_61_wd;
	// Trace: design.sv:91093:3
	wire ie0_1_e_61_we;
	// Trace: design.sv:91094:3
	wire ie0_1_e_62_qs;
	// Trace: design.sv:91095:3
	wire ie0_1_e_62_wd;
	// Trace: design.sv:91096:3
	wire ie0_1_e_62_we;
	// Trace: design.sv:91097:3
	wire ie0_1_e_63_qs;
	// Trace: design.sv:91098:3
	wire ie0_1_e_63_wd;
	// Trace: design.sv:91099:3
	wire ie0_1_e_63_we;
	// Trace: design.sv:91100:3
	wire [2:0] threshold0_qs;
	// Trace: design.sv:91101:3
	wire [2:0] threshold0_wd;
	// Trace: design.sv:91102:3
	wire threshold0_we;
	// Trace: design.sv:91103:3
	wire [5:0] cc0_qs;
	// Trace: design.sv:91104:3
	wire [5:0] cc0_wd;
	// Trace: design.sv:91105:3
	wire cc0_we;
	// Trace: design.sv:91106:3
	wire cc0_re;
	// Trace: design.sv:91107:3
	wire msip0_qs;
	// Trace: design.sv:91108:3
	wire msip0_wd;
	// Trace: design.sv:91109:3
	wire msip0_we;
	// Trace: design.sv:91117:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_0_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_0_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_0_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_0_ext_wd_0),
		.de(hw2reg[6]),
		.d(hw2reg[7]),
		.qe(),
		.q(),
		.qs(ip_0_p_0_qs)
	);
	// Trace: design.sv:91142:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_1_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_1_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_1_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_1_ext_wd_0),
		.de(hw2reg[8]),
		.d(hw2reg[9]),
		.qe(),
		.q(),
		.qs(ip_0_p_1_qs)
	);
	// Trace: design.sv:91167:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_2_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_2_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_2_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_2_ext_wd_0),
		.de(hw2reg[10]),
		.d(hw2reg[11]),
		.qe(),
		.q(),
		.qs(ip_0_p_2_qs)
	);
	// Trace: design.sv:91192:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_3_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_3_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_3_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_3_ext_wd_0),
		.de(hw2reg[12]),
		.d(hw2reg[13]),
		.qe(),
		.q(),
		.qs(ip_0_p_3_qs)
	);
	// Trace: design.sv:91217:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_4_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_4_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_4_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_4_ext_wd_0),
		.de(hw2reg[14]),
		.d(hw2reg[15]),
		.qe(),
		.q(),
		.qs(ip_0_p_4_qs)
	);
	// Trace: design.sv:91242:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_5_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_5_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_5_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_5_ext_wd_0),
		.de(hw2reg[16]),
		.d(hw2reg[17]),
		.qe(),
		.q(),
		.qs(ip_0_p_5_qs)
	);
	// Trace: design.sv:91267:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_6_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_6_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_6_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_6_ext_wd_0),
		.de(hw2reg[18]),
		.d(hw2reg[19]),
		.qe(),
		.q(),
		.qs(ip_0_p_6_qs)
	);
	// Trace: design.sv:91292:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_7_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_7_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_7_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_7_ext_wd_0),
		.de(hw2reg[20]),
		.d(hw2reg[21]),
		.qe(),
		.q(),
		.qs(ip_0_p_7_qs)
	);
	// Trace: design.sv:91317:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_8_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_8_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_8_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_8_ext_wd_0),
		.de(hw2reg[22]),
		.d(hw2reg[23]),
		.qe(),
		.q(),
		.qs(ip_0_p_8_qs)
	);
	// Trace: design.sv:91342:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_9_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_9_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_9_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_9_ext_wd_0),
		.de(hw2reg[24]),
		.d(hw2reg[25]),
		.qe(),
		.q(),
		.qs(ip_0_p_9_qs)
	);
	// Trace: design.sv:91367:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_10_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_10_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_10_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_10_ext_wd_0),
		.de(hw2reg[26]),
		.d(hw2reg[27]),
		.qe(),
		.q(),
		.qs(ip_0_p_10_qs)
	);
	// Trace: design.sv:91392:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_11_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_11_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_11_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_11_ext_wd_0),
		.de(hw2reg[28]),
		.d(hw2reg[29]),
		.qe(),
		.q(),
		.qs(ip_0_p_11_qs)
	);
	// Trace: design.sv:91417:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_12_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_12_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_12_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_12_ext_wd_0),
		.de(hw2reg[30]),
		.d(hw2reg[31]),
		.qe(),
		.q(),
		.qs(ip_0_p_12_qs)
	);
	// Trace: design.sv:91442:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_13_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_13_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_13_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_13_ext_wd_0),
		.de(hw2reg[32]),
		.d(hw2reg[33]),
		.qe(),
		.q(),
		.qs(ip_0_p_13_qs)
	);
	// Trace: design.sv:91467:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_14_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_14_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_14_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_14_ext_wd_0),
		.de(hw2reg[34]),
		.d(hw2reg[35]),
		.qe(),
		.q(),
		.qs(ip_0_p_14_qs)
	);
	// Trace: design.sv:91492:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_15_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_15_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_15_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_15_ext_wd_0),
		.de(hw2reg[36]),
		.d(hw2reg[37]),
		.qe(),
		.q(),
		.qs(ip_0_p_15_qs)
	);
	// Trace: design.sv:91517:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_16_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_16_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_16_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_16_ext_wd_0),
		.de(hw2reg[38]),
		.d(hw2reg[39]),
		.qe(),
		.q(),
		.qs(ip_0_p_16_qs)
	);
	// Trace: design.sv:91542:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_17_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_17_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_17_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_17_ext_wd_0),
		.de(hw2reg[40]),
		.d(hw2reg[41]),
		.qe(),
		.q(),
		.qs(ip_0_p_17_qs)
	);
	// Trace: design.sv:91567:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_18_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_18_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_18_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_18_ext_wd_0),
		.de(hw2reg[42]),
		.d(hw2reg[43]),
		.qe(),
		.q(),
		.qs(ip_0_p_18_qs)
	);
	// Trace: design.sv:91592:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_19_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_19_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_19_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_19_ext_wd_0),
		.de(hw2reg[44]),
		.d(hw2reg[45]),
		.qe(),
		.q(),
		.qs(ip_0_p_19_qs)
	);
	// Trace: design.sv:91617:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_20_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_20_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_20_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_20_ext_wd_0),
		.de(hw2reg[46]),
		.d(hw2reg[47]),
		.qe(),
		.q(),
		.qs(ip_0_p_20_qs)
	);
	// Trace: design.sv:91642:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_21_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_21_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_21_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_21_ext_wd_0),
		.de(hw2reg[48]),
		.d(hw2reg[49]),
		.qe(),
		.q(),
		.qs(ip_0_p_21_qs)
	);
	// Trace: design.sv:91667:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_22_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_22_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_22_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_22_ext_wd_0),
		.de(hw2reg[50]),
		.d(hw2reg[51]),
		.qe(),
		.q(),
		.qs(ip_0_p_22_qs)
	);
	// Trace: design.sv:91692:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_23_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_23_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_23_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_23_ext_wd_0),
		.de(hw2reg[52]),
		.d(hw2reg[53]),
		.qe(),
		.q(),
		.qs(ip_0_p_23_qs)
	);
	// Trace: design.sv:91717:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_24_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_24_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_24_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_24_ext_wd_0),
		.de(hw2reg[54]),
		.d(hw2reg[55]),
		.qe(),
		.q(),
		.qs(ip_0_p_24_qs)
	);
	// Trace: design.sv:91742:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_25_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_25_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_25_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_25_ext_wd_0),
		.de(hw2reg[56]),
		.d(hw2reg[57]),
		.qe(),
		.q(),
		.qs(ip_0_p_25_qs)
	);
	// Trace: design.sv:91767:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_26_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_26_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_26_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_26_ext_wd_0),
		.de(hw2reg[58]),
		.d(hw2reg[59]),
		.qe(),
		.q(),
		.qs(ip_0_p_26_qs)
	);
	// Trace: design.sv:91792:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_27_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_27_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_27_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_27_ext_wd_0),
		.de(hw2reg[60]),
		.d(hw2reg[61]),
		.qe(),
		.q(),
		.qs(ip_0_p_27_qs)
	);
	// Trace: design.sv:91817:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_28_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_28_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_28_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_28_ext_wd_0),
		.de(hw2reg[62]),
		.d(hw2reg[63]),
		.qe(),
		.q(),
		.qs(ip_0_p_28_qs)
	);
	// Trace: design.sv:91842:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_29_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_29_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_29_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_29_ext_wd_0),
		.de(hw2reg[64]),
		.d(hw2reg[65]),
		.qe(),
		.q(),
		.qs(ip_0_p_29_qs)
	);
	// Trace: design.sv:91867:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_30_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_30_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_30_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_30_ext_wd_0),
		.de(hw2reg[66]),
		.d(hw2reg[67]),
		.qe(),
		.q(),
		.qs(ip_0_p_30_qs)
	);
	// Trace: design.sv:91892:3
	localparam signed [31:0] sv2v_uu_u_ip_0_p_31_DW = 1;
	// removed localparam type sv2v_uu_u_ip_0_p_31_wd
	localparam [0:0] sv2v_uu_u_ip_0_p_31_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_0_p_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_0_p_31_ext_wd_0),
		.de(hw2reg[68]),
		.d(hw2reg[69]),
		.qe(),
		.q(),
		.qs(ip_0_p_31_qs)
	);
	// Trace: design.sv:91920:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_32_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_32_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_32_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_32(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_32_ext_wd_0),
		.de(hw2reg[70]),
		.d(hw2reg[71]),
		.qe(),
		.q(),
		.qs(ip_1_p_32_qs)
	);
	// Trace: design.sv:91945:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_33_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_33_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_33_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_33(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_33_ext_wd_0),
		.de(hw2reg[72]),
		.d(hw2reg[73]),
		.qe(),
		.q(),
		.qs(ip_1_p_33_qs)
	);
	// Trace: design.sv:91970:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_34_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_34_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_34_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_34(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_34_ext_wd_0),
		.de(hw2reg[74]),
		.d(hw2reg[75]),
		.qe(),
		.q(),
		.qs(ip_1_p_34_qs)
	);
	// Trace: design.sv:91995:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_35_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_35_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_35_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_35(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_35_ext_wd_0),
		.de(hw2reg[76]),
		.d(hw2reg[77]),
		.qe(),
		.q(),
		.qs(ip_1_p_35_qs)
	);
	// Trace: design.sv:92020:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_36_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_36_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_36_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_36(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_36_ext_wd_0),
		.de(hw2reg[78]),
		.d(hw2reg[79]),
		.qe(),
		.q(),
		.qs(ip_1_p_36_qs)
	);
	// Trace: design.sv:92045:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_37_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_37_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_37_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_37(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_37_ext_wd_0),
		.de(hw2reg[80]),
		.d(hw2reg[81]),
		.qe(),
		.q(),
		.qs(ip_1_p_37_qs)
	);
	// Trace: design.sv:92070:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_38_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_38_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_38_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_38(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_38_ext_wd_0),
		.de(hw2reg[82]),
		.d(hw2reg[83]),
		.qe(),
		.q(),
		.qs(ip_1_p_38_qs)
	);
	// Trace: design.sv:92095:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_39_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_39_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_39_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_39(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_39_ext_wd_0),
		.de(hw2reg[84]),
		.d(hw2reg[85]),
		.qe(),
		.q(),
		.qs(ip_1_p_39_qs)
	);
	// Trace: design.sv:92120:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_40_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_40_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_40_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_40(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_40_ext_wd_0),
		.de(hw2reg[86]),
		.d(hw2reg[87]),
		.qe(),
		.q(),
		.qs(ip_1_p_40_qs)
	);
	// Trace: design.sv:92145:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_41_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_41_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_41_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_41(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_41_ext_wd_0),
		.de(hw2reg[88]),
		.d(hw2reg[89]),
		.qe(),
		.q(),
		.qs(ip_1_p_41_qs)
	);
	// Trace: design.sv:92170:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_42_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_42_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_42_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_42(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_42_ext_wd_0),
		.de(hw2reg[90]),
		.d(hw2reg[91]),
		.qe(),
		.q(),
		.qs(ip_1_p_42_qs)
	);
	// Trace: design.sv:92195:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_43_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_43_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_43_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_43(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_43_ext_wd_0),
		.de(hw2reg[92]),
		.d(hw2reg[93]),
		.qe(),
		.q(),
		.qs(ip_1_p_43_qs)
	);
	// Trace: design.sv:92220:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_44_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_44_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_44_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_44(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_44_ext_wd_0),
		.de(hw2reg[94]),
		.d(hw2reg[95]),
		.qe(),
		.q(),
		.qs(ip_1_p_44_qs)
	);
	// Trace: design.sv:92245:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_45_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_45_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_45_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_45(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_45_ext_wd_0),
		.de(hw2reg[96]),
		.d(hw2reg[97]),
		.qe(),
		.q(),
		.qs(ip_1_p_45_qs)
	);
	// Trace: design.sv:92270:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_46_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_46_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_46_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_46(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_46_ext_wd_0),
		.de(hw2reg[98]),
		.d(hw2reg[99]),
		.qe(),
		.q(),
		.qs(ip_1_p_46_qs)
	);
	// Trace: design.sv:92295:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_47_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_47_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_47_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_47(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_47_ext_wd_0),
		.de(hw2reg[100]),
		.d(hw2reg[101]),
		.qe(),
		.q(),
		.qs(ip_1_p_47_qs)
	);
	// Trace: design.sv:92320:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_48_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_48_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_48_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_48(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_48_ext_wd_0),
		.de(hw2reg[102]),
		.d(hw2reg[103]),
		.qe(),
		.q(),
		.qs(ip_1_p_48_qs)
	);
	// Trace: design.sv:92345:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_49_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_49_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_49_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_49(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_49_ext_wd_0),
		.de(hw2reg[104]),
		.d(hw2reg[105]),
		.qe(),
		.q(),
		.qs(ip_1_p_49_qs)
	);
	// Trace: design.sv:92370:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_50_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_50_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_50_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_50(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_50_ext_wd_0),
		.de(hw2reg[106]),
		.d(hw2reg[107]),
		.qe(),
		.q(),
		.qs(ip_1_p_50_qs)
	);
	// Trace: design.sv:92395:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_51_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_51_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_51_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_51(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_51_ext_wd_0),
		.de(hw2reg[108]),
		.d(hw2reg[109]),
		.qe(),
		.q(),
		.qs(ip_1_p_51_qs)
	);
	// Trace: design.sv:92420:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_52_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_52_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_52_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_52(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_52_ext_wd_0),
		.de(hw2reg[110]),
		.d(hw2reg[111]),
		.qe(),
		.q(),
		.qs(ip_1_p_52_qs)
	);
	// Trace: design.sv:92445:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_53_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_53_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_53_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_53(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_53_ext_wd_0),
		.de(hw2reg[112]),
		.d(hw2reg[113]),
		.qe(),
		.q(),
		.qs(ip_1_p_53_qs)
	);
	// Trace: design.sv:92470:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_54_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_54_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_54_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_54(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_54_ext_wd_0),
		.de(hw2reg[114]),
		.d(hw2reg[115]),
		.qe(),
		.q(),
		.qs(ip_1_p_54_qs)
	);
	// Trace: design.sv:92495:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_55_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_55_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_55_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_55(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_55_ext_wd_0),
		.de(hw2reg[116]),
		.d(hw2reg[117]),
		.qe(),
		.q(),
		.qs(ip_1_p_55_qs)
	);
	// Trace: design.sv:92520:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_56_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_56_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_56_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_56(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_56_ext_wd_0),
		.de(hw2reg[118]),
		.d(hw2reg[119]),
		.qe(),
		.q(),
		.qs(ip_1_p_56_qs)
	);
	// Trace: design.sv:92545:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_57_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_57_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_57_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_57(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_57_ext_wd_0),
		.de(hw2reg[120]),
		.d(hw2reg[121]),
		.qe(),
		.q(),
		.qs(ip_1_p_57_qs)
	);
	// Trace: design.sv:92570:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_58_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_58_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_58_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_58(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_58_ext_wd_0),
		.de(hw2reg[122]),
		.d(hw2reg[123]),
		.qe(),
		.q(),
		.qs(ip_1_p_58_qs)
	);
	// Trace: design.sv:92595:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_59_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_59_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_59_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_59(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_59_ext_wd_0),
		.de(hw2reg[124]),
		.d(hw2reg[125]),
		.qe(),
		.q(),
		.qs(ip_1_p_59_qs)
	);
	// Trace: design.sv:92620:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_60_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_60_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_60_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_60(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_60_ext_wd_0),
		.de(hw2reg[126]),
		.d(hw2reg[127]),
		.qe(),
		.q(),
		.qs(ip_1_p_60_qs)
	);
	// Trace: design.sv:92645:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_61_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_61_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_61_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_61(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_61_ext_wd_0),
		.de(hw2reg[128]),
		.d(hw2reg[129]),
		.qe(),
		.q(),
		.qs(ip_1_p_61_qs)
	);
	// Trace: design.sv:92670:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_62_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_62_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_62_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_62(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_62_ext_wd_0),
		.de(hw2reg[130]),
		.d(hw2reg[131]),
		.qe(),
		.q(),
		.qs(ip_1_p_62_qs)
	);
	// Trace: design.sv:92695:3
	localparam signed [31:0] sv2v_uu_u_ip_1_p_63_DW = 1;
	// removed localparam type sv2v_uu_u_ip_1_p_63_wd
	localparam [0:0] sv2v_uu_u_ip_1_p_63_ext_wd_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RO"),
		.RESVAL(1'h0)
	) u_ip_1_p_63(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(sv2v_uu_u_ip_1_p_63_ext_wd_0),
		.de(hw2reg[132]),
		.d(hw2reg[133]),
		.qe(),
		.q(),
		.qs(ip_1_p_63_qs)
	);
	// Trace: design.sv:92725:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_0_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_0_d
	localparam [0:0] sv2v_uu_u_le_0_le_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_0_we),
		.wd(le_0_le_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_0_ext_d_0),
		.qe(),
		.q(reg2hw[268]),
		.qs(le_0_le_0_qs)
	);
	// Trace: design.sv:92751:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_1_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_1_d
	localparam [0:0] sv2v_uu_u_le_0_le_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_1_we),
		.wd(le_0_le_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_1_ext_d_0),
		.qe(),
		.q(reg2hw[269]),
		.qs(le_0_le_1_qs)
	);
	// Trace: design.sv:92777:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_2_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_2_d
	localparam [0:0] sv2v_uu_u_le_0_le_2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_2_we),
		.wd(le_0_le_2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_2_ext_d_0),
		.qe(),
		.q(reg2hw[270]),
		.qs(le_0_le_2_qs)
	);
	// Trace: design.sv:92803:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_3_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_3_d
	localparam [0:0] sv2v_uu_u_le_0_le_3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_3_we),
		.wd(le_0_le_3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_3_ext_d_0),
		.qe(),
		.q(reg2hw[271]),
		.qs(le_0_le_3_qs)
	);
	// Trace: design.sv:92829:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_4_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_4_d
	localparam [0:0] sv2v_uu_u_le_0_le_4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_4_we),
		.wd(le_0_le_4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_4_ext_d_0),
		.qe(),
		.q(reg2hw[272]),
		.qs(le_0_le_4_qs)
	);
	// Trace: design.sv:92855:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_5_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_5_d
	localparam [0:0] sv2v_uu_u_le_0_le_5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_5_we),
		.wd(le_0_le_5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_5_ext_d_0),
		.qe(),
		.q(reg2hw[273]),
		.qs(le_0_le_5_qs)
	);
	// Trace: design.sv:92881:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_6_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_6_d
	localparam [0:0] sv2v_uu_u_le_0_le_6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_6_we),
		.wd(le_0_le_6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_6_ext_d_0),
		.qe(),
		.q(reg2hw[274]),
		.qs(le_0_le_6_qs)
	);
	// Trace: design.sv:92907:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_7_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_7_d
	localparam [0:0] sv2v_uu_u_le_0_le_7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_7_we),
		.wd(le_0_le_7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_7_ext_d_0),
		.qe(),
		.q(reg2hw[275]),
		.qs(le_0_le_7_qs)
	);
	// Trace: design.sv:92933:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_8_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_8_d
	localparam [0:0] sv2v_uu_u_le_0_le_8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_8_we),
		.wd(le_0_le_8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_8_ext_d_0),
		.qe(),
		.q(reg2hw[276]),
		.qs(le_0_le_8_qs)
	);
	// Trace: design.sv:92959:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_9_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_9_d
	localparam [0:0] sv2v_uu_u_le_0_le_9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_9_we),
		.wd(le_0_le_9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_9_ext_d_0),
		.qe(),
		.q(reg2hw[277]),
		.qs(le_0_le_9_qs)
	);
	// Trace: design.sv:92985:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_10_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_10_d
	localparam [0:0] sv2v_uu_u_le_0_le_10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_10_we),
		.wd(le_0_le_10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_10_ext_d_0),
		.qe(),
		.q(reg2hw[278]),
		.qs(le_0_le_10_qs)
	);
	// Trace: design.sv:93011:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_11_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_11_d
	localparam [0:0] sv2v_uu_u_le_0_le_11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_11_we),
		.wd(le_0_le_11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_11_ext_d_0),
		.qe(),
		.q(reg2hw[279]),
		.qs(le_0_le_11_qs)
	);
	// Trace: design.sv:93037:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_12_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_12_d
	localparam [0:0] sv2v_uu_u_le_0_le_12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_12_we),
		.wd(le_0_le_12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_12_ext_d_0),
		.qe(),
		.q(reg2hw[280]),
		.qs(le_0_le_12_qs)
	);
	// Trace: design.sv:93063:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_13_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_13_d
	localparam [0:0] sv2v_uu_u_le_0_le_13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_13_we),
		.wd(le_0_le_13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_13_ext_d_0),
		.qe(),
		.q(reg2hw[281]),
		.qs(le_0_le_13_qs)
	);
	// Trace: design.sv:93089:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_14_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_14_d
	localparam [0:0] sv2v_uu_u_le_0_le_14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_14_we),
		.wd(le_0_le_14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_14_ext_d_0),
		.qe(),
		.q(reg2hw[282]),
		.qs(le_0_le_14_qs)
	);
	// Trace: design.sv:93115:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_15_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_15_d
	localparam [0:0] sv2v_uu_u_le_0_le_15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_15_we),
		.wd(le_0_le_15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_15_ext_d_0),
		.qe(),
		.q(reg2hw[283]),
		.qs(le_0_le_15_qs)
	);
	// Trace: design.sv:93141:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_16_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_16_d
	localparam [0:0] sv2v_uu_u_le_0_le_16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_16_we),
		.wd(le_0_le_16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_16_ext_d_0),
		.qe(),
		.q(reg2hw[284]),
		.qs(le_0_le_16_qs)
	);
	// Trace: design.sv:93167:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_17_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_17_d
	localparam [0:0] sv2v_uu_u_le_0_le_17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_17_we),
		.wd(le_0_le_17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_17_ext_d_0),
		.qe(),
		.q(reg2hw[285]),
		.qs(le_0_le_17_qs)
	);
	// Trace: design.sv:93193:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_18_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_18_d
	localparam [0:0] sv2v_uu_u_le_0_le_18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_18_we),
		.wd(le_0_le_18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_18_ext_d_0),
		.qe(),
		.q(reg2hw[286]),
		.qs(le_0_le_18_qs)
	);
	// Trace: design.sv:93219:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_19_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_19_d
	localparam [0:0] sv2v_uu_u_le_0_le_19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_19_we),
		.wd(le_0_le_19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_19_ext_d_0),
		.qe(),
		.q(reg2hw[287]),
		.qs(le_0_le_19_qs)
	);
	// Trace: design.sv:93245:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_20_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_20_d
	localparam [0:0] sv2v_uu_u_le_0_le_20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_20_we),
		.wd(le_0_le_20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_20_ext_d_0),
		.qe(),
		.q(reg2hw[288]),
		.qs(le_0_le_20_qs)
	);
	// Trace: design.sv:93271:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_21_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_21_d
	localparam [0:0] sv2v_uu_u_le_0_le_21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_21_we),
		.wd(le_0_le_21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_21_ext_d_0),
		.qe(),
		.q(reg2hw[289]),
		.qs(le_0_le_21_qs)
	);
	// Trace: design.sv:93297:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_22_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_22_d
	localparam [0:0] sv2v_uu_u_le_0_le_22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_22_we),
		.wd(le_0_le_22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_22_ext_d_0),
		.qe(),
		.q(reg2hw[290]),
		.qs(le_0_le_22_qs)
	);
	// Trace: design.sv:93323:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_23_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_23_d
	localparam [0:0] sv2v_uu_u_le_0_le_23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_23_we),
		.wd(le_0_le_23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_23_ext_d_0),
		.qe(),
		.q(reg2hw[291]),
		.qs(le_0_le_23_qs)
	);
	// Trace: design.sv:93349:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_24_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_24_d
	localparam [0:0] sv2v_uu_u_le_0_le_24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_24_we),
		.wd(le_0_le_24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_24_ext_d_0),
		.qe(),
		.q(reg2hw[292]),
		.qs(le_0_le_24_qs)
	);
	// Trace: design.sv:93375:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_25_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_25_d
	localparam [0:0] sv2v_uu_u_le_0_le_25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_25_we),
		.wd(le_0_le_25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_25_ext_d_0),
		.qe(),
		.q(reg2hw[293]),
		.qs(le_0_le_25_qs)
	);
	// Trace: design.sv:93401:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_26_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_26_d
	localparam [0:0] sv2v_uu_u_le_0_le_26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_26_we),
		.wd(le_0_le_26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_26_ext_d_0),
		.qe(),
		.q(reg2hw[294]),
		.qs(le_0_le_26_qs)
	);
	// Trace: design.sv:93427:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_27_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_27_d
	localparam [0:0] sv2v_uu_u_le_0_le_27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_27_we),
		.wd(le_0_le_27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_27_ext_d_0),
		.qe(),
		.q(reg2hw[295]),
		.qs(le_0_le_27_qs)
	);
	// Trace: design.sv:93453:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_28_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_28_d
	localparam [0:0] sv2v_uu_u_le_0_le_28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_28_we),
		.wd(le_0_le_28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_28_ext_d_0),
		.qe(),
		.q(reg2hw[296]),
		.qs(le_0_le_28_qs)
	);
	// Trace: design.sv:93479:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_29_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_29_d
	localparam [0:0] sv2v_uu_u_le_0_le_29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_29_we),
		.wd(le_0_le_29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_29_ext_d_0),
		.qe(),
		.q(reg2hw[297]),
		.qs(le_0_le_29_qs)
	);
	// Trace: design.sv:93505:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_30_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_30_d
	localparam [0:0] sv2v_uu_u_le_0_le_30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_30_we),
		.wd(le_0_le_30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_30_ext_d_0),
		.qe(),
		.q(reg2hw[298]),
		.qs(le_0_le_30_qs)
	);
	// Trace: design.sv:93531:3
	localparam signed [31:0] sv2v_uu_u_le_0_le_31_DW = 1;
	// removed localparam type sv2v_uu_u_le_0_le_31_d
	localparam [0:0] sv2v_uu_u_le_0_le_31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_0_le_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_0_le_31_we),
		.wd(le_0_le_31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_0_le_31_ext_d_0),
		.qe(),
		.q(reg2hw[299]),
		.qs(le_0_le_31_qs)
	);
	// Trace: design.sv:93560:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_32_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_32_d
	localparam [0:0] sv2v_uu_u_le_1_le_32_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_32(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_32_we),
		.wd(le_1_le_32_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_32_ext_d_0),
		.qe(),
		.q(reg2hw[300]),
		.qs(le_1_le_32_qs)
	);
	// Trace: design.sv:93586:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_33_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_33_d
	localparam [0:0] sv2v_uu_u_le_1_le_33_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_33(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_33_we),
		.wd(le_1_le_33_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_33_ext_d_0),
		.qe(),
		.q(reg2hw[301]),
		.qs(le_1_le_33_qs)
	);
	// Trace: design.sv:93612:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_34_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_34_d
	localparam [0:0] sv2v_uu_u_le_1_le_34_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_34(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_34_we),
		.wd(le_1_le_34_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_34_ext_d_0),
		.qe(),
		.q(reg2hw[302]),
		.qs(le_1_le_34_qs)
	);
	// Trace: design.sv:93638:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_35_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_35_d
	localparam [0:0] sv2v_uu_u_le_1_le_35_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_35(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_35_we),
		.wd(le_1_le_35_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_35_ext_d_0),
		.qe(),
		.q(reg2hw[303]),
		.qs(le_1_le_35_qs)
	);
	// Trace: design.sv:93664:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_36_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_36_d
	localparam [0:0] sv2v_uu_u_le_1_le_36_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_36(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_36_we),
		.wd(le_1_le_36_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_36_ext_d_0),
		.qe(),
		.q(reg2hw[304]),
		.qs(le_1_le_36_qs)
	);
	// Trace: design.sv:93690:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_37_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_37_d
	localparam [0:0] sv2v_uu_u_le_1_le_37_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_37(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_37_we),
		.wd(le_1_le_37_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_37_ext_d_0),
		.qe(),
		.q(reg2hw[305]),
		.qs(le_1_le_37_qs)
	);
	// Trace: design.sv:93716:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_38_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_38_d
	localparam [0:0] sv2v_uu_u_le_1_le_38_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_38(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_38_we),
		.wd(le_1_le_38_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_38_ext_d_0),
		.qe(),
		.q(reg2hw[306]),
		.qs(le_1_le_38_qs)
	);
	// Trace: design.sv:93742:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_39_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_39_d
	localparam [0:0] sv2v_uu_u_le_1_le_39_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_39(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_39_we),
		.wd(le_1_le_39_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_39_ext_d_0),
		.qe(),
		.q(reg2hw[307]),
		.qs(le_1_le_39_qs)
	);
	// Trace: design.sv:93768:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_40_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_40_d
	localparam [0:0] sv2v_uu_u_le_1_le_40_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_40(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_40_we),
		.wd(le_1_le_40_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_40_ext_d_0),
		.qe(),
		.q(reg2hw[308]),
		.qs(le_1_le_40_qs)
	);
	// Trace: design.sv:93794:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_41_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_41_d
	localparam [0:0] sv2v_uu_u_le_1_le_41_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_41(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_41_we),
		.wd(le_1_le_41_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_41_ext_d_0),
		.qe(),
		.q(reg2hw[309]),
		.qs(le_1_le_41_qs)
	);
	// Trace: design.sv:93820:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_42_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_42_d
	localparam [0:0] sv2v_uu_u_le_1_le_42_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_42(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_42_we),
		.wd(le_1_le_42_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_42_ext_d_0),
		.qe(),
		.q(reg2hw[310]),
		.qs(le_1_le_42_qs)
	);
	// Trace: design.sv:93846:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_43_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_43_d
	localparam [0:0] sv2v_uu_u_le_1_le_43_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_43(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_43_we),
		.wd(le_1_le_43_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_43_ext_d_0),
		.qe(),
		.q(reg2hw[311]),
		.qs(le_1_le_43_qs)
	);
	// Trace: design.sv:93872:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_44_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_44_d
	localparam [0:0] sv2v_uu_u_le_1_le_44_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_44(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_44_we),
		.wd(le_1_le_44_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_44_ext_d_0),
		.qe(),
		.q(reg2hw[312]),
		.qs(le_1_le_44_qs)
	);
	// Trace: design.sv:93898:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_45_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_45_d
	localparam [0:0] sv2v_uu_u_le_1_le_45_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_45(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_45_we),
		.wd(le_1_le_45_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_45_ext_d_0),
		.qe(),
		.q(reg2hw[313]),
		.qs(le_1_le_45_qs)
	);
	// Trace: design.sv:93924:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_46_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_46_d
	localparam [0:0] sv2v_uu_u_le_1_le_46_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_46(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_46_we),
		.wd(le_1_le_46_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_46_ext_d_0),
		.qe(),
		.q(reg2hw[314]),
		.qs(le_1_le_46_qs)
	);
	// Trace: design.sv:93950:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_47_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_47_d
	localparam [0:0] sv2v_uu_u_le_1_le_47_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_47(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_47_we),
		.wd(le_1_le_47_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_47_ext_d_0),
		.qe(),
		.q(reg2hw[315]),
		.qs(le_1_le_47_qs)
	);
	// Trace: design.sv:93976:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_48_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_48_d
	localparam [0:0] sv2v_uu_u_le_1_le_48_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_48(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_48_we),
		.wd(le_1_le_48_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_48_ext_d_0),
		.qe(),
		.q(reg2hw[316]),
		.qs(le_1_le_48_qs)
	);
	// Trace: design.sv:94002:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_49_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_49_d
	localparam [0:0] sv2v_uu_u_le_1_le_49_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_49(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_49_we),
		.wd(le_1_le_49_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_49_ext_d_0),
		.qe(),
		.q(reg2hw[317]),
		.qs(le_1_le_49_qs)
	);
	// Trace: design.sv:94028:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_50_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_50_d
	localparam [0:0] sv2v_uu_u_le_1_le_50_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_50(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_50_we),
		.wd(le_1_le_50_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_50_ext_d_0),
		.qe(),
		.q(reg2hw[318]),
		.qs(le_1_le_50_qs)
	);
	// Trace: design.sv:94054:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_51_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_51_d
	localparam [0:0] sv2v_uu_u_le_1_le_51_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_51(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_51_we),
		.wd(le_1_le_51_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_51_ext_d_0),
		.qe(),
		.q(reg2hw[319]),
		.qs(le_1_le_51_qs)
	);
	// Trace: design.sv:94080:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_52_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_52_d
	localparam [0:0] sv2v_uu_u_le_1_le_52_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_52(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_52_we),
		.wd(le_1_le_52_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_52_ext_d_0),
		.qe(),
		.q(reg2hw[320]),
		.qs(le_1_le_52_qs)
	);
	// Trace: design.sv:94106:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_53_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_53_d
	localparam [0:0] sv2v_uu_u_le_1_le_53_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_53(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_53_we),
		.wd(le_1_le_53_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_53_ext_d_0),
		.qe(),
		.q(reg2hw[321]),
		.qs(le_1_le_53_qs)
	);
	// Trace: design.sv:94132:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_54_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_54_d
	localparam [0:0] sv2v_uu_u_le_1_le_54_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_54(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_54_we),
		.wd(le_1_le_54_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_54_ext_d_0),
		.qe(),
		.q(reg2hw[322]),
		.qs(le_1_le_54_qs)
	);
	// Trace: design.sv:94158:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_55_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_55_d
	localparam [0:0] sv2v_uu_u_le_1_le_55_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_55(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_55_we),
		.wd(le_1_le_55_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_55_ext_d_0),
		.qe(),
		.q(reg2hw[323]),
		.qs(le_1_le_55_qs)
	);
	// Trace: design.sv:94184:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_56_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_56_d
	localparam [0:0] sv2v_uu_u_le_1_le_56_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_56(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_56_we),
		.wd(le_1_le_56_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_56_ext_d_0),
		.qe(),
		.q(reg2hw[324]),
		.qs(le_1_le_56_qs)
	);
	// Trace: design.sv:94210:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_57_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_57_d
	localparam [0:0] sv2v_uu_u_le_1_le_57_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_57(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_57_we),
		.wd(le_1_le_57_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_57_ext_d_0),
		.qe(),
		.q(reg2hw[325]),
		.qs(le_1_le_57_qs)
	);
	// Trace: design.sv:94236:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_58_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_58_d
	localparam [0:0] sv2v_uu_u_le_1_le_58_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_58(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_58_we),
		.wd(le_1_le_58_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_58_ext_d_0),
		.qe(),
		.q(reg2hw[326]),
		.qs(le_1_le_58_qs)
	);
	// Trace: design.sv:94262:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_59_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_59_d
	localparam [0:0] sv2v_uu_u_le_1_le_59_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_59(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_59_we),
		.wd(le_1_le_59_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_59_ext_d_0),
		.qe(),
		.q(reg2hw[327]),
		.qs(le_1_le_59_qs)
	);
	// Trace: design.sv:94288:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_60_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_60_d
	localparam [0:0] sv2v_uu_u_le_1_le_60_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_60(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_60_we),
		.wd(le_1_le_60_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_60_ext_d_0),
		.qe(),
		.q(reg2hw[328]),
		.qs(le_1_le_60_qs)
	);
	// Trace: design.sv:94314:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_61_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_61_d
	localparam [0:0] sv2v_uu_u_le_1_le_61_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_61(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_61_we),
		.wd(le_1_le_61_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_61_ext_d_0),
		.qe(),
		.q(reg2hw[329]),
		.qs(le_1_le_61_qs)
	);
	// Trace: design.sv:94340:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_62_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_62_d
	localparam [0:0] sv2v_uu_u_le_1_le_62_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_62(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_62_we),
		.wd(le_1_le_62_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_62_ext_d_0),
		.qe(),
		.q(reg2hw[330]),
		.qs(le_1_le_62_qs)
	);
	// Trace: design.sv:94366:3
	localparam signed [31:0] sv2v_uu_u_le_1_le_63_DW = 1;
	// removed localparam type sv2v_uu_u_le_1_le_63_d
	localparam [0:0] sv2v_uu_u_le_1_le_63_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_le_1_le_63(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(le_1_le_63_we),
		.wd(le_1_le_63_wd),
		.de(1'b0),
		.d(sv2v_uu_u_le_1_le_63_ext_d_0),
		.qe(),
		.q(reg2hw[331]),
		.qs(le_1_le_63_qs)
	);
	// Trace: design.sv:94394:3
	localparam signed [31:0] sv2v_uu_u_prio0_DW = 3;
	// removed localparam type sv2v_uu_u_prio0_d
	localparam [2:0] sv2v_uu_u_prio0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio0_we),
		.wd(prio0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio0_ext_d_0),
		.qe(),
		.q(reg2hw[267-:3]),
		.qs(prio0_qs)
	);
	// Trace: design.sv:94421:3
	localparam signed [31:0] sv2v_uu_u_prio1_DW = 3;
	// removed localparam type sv2v_uu_u_prio1_d
	localparam [2:0] sv2v_uu_u_prio1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio1_we),
		.wd(prio1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio1_ext_d_0),
		.qe(),
		.q(reg2hw[264-:3]),
		.qs(prio1_qs)
	);
	// Trace: design.sv:94448:3
	localparam signed [31:0] sv2v_uu_u_prio2_DW = 3;
	// removed localparam type sv2v_uu_u_prio2_d
	localparam [2:0] sv2v_uu_u_prio2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio2_we),
		.wd(prio2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio2_ext_d_0),
		.qe(),
		.q(reg2hw[261-:3]),
		.qs(prio2_qs)
	);
	// Trace: design.sv:94475:3
	localparam signed [31:0] sv2v_uu_u_prio3_DW = 3;
	// removed localparam type sv2v_uu_u_prio3_d
	localparam [2:0] sv2v_uu_u_prio3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio3_we),
		.wd(prio3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio3_ext_d_0),
		.qe(),
		.q(reg2hw[258-:3]),
		.qs(prio3_qs)
	);
	// Trace: design.sv:94502:3
	localparam signed [31:0] sv2v_uu_u_prio4_DW = 3;
	// removed localparam type sv2v_uu_u_prio4_d
	localparam [2:0] sv2v_uu_u_prio4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio4_we),
		.wd(prio4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio4_ext_d_0),
		.qe(),
		.q(reg2hw[255-:3]),
		.qs(prio4_qs)
	);
	// Trace: design.sv:94529:3
	localparam signed [31:0] sv2v_uu_u_prio5_DW = 3;
	// removed localparam type sv2v_uu_u_prio5_d
	localparam [2:0] sv2v_uu_u_prio5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio5_we),
		.wd(prio5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio5_ext_d_0),
		.qe(),
		.q(reg2hw[252-:3]),
		.qs(prio5_qs)
	);
	// Trace: design.sv:94556:3
	localparam signed [31:0] sv2v_uu_u_prio6_DW = 3;
	// removed localparam type sv2v_uu_u_prio6_d
	localparam [2:0] sv2v_uu_u_prio6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio6_we),
		.wd(prio6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio6_ext_d_0),
		.qe(),
		.q(reg2hw[249-:3]),
		.qs(prio6_qs)
	);
	// Trace: design.sv:94583:3
	localparam signed [31:0] sv2v_uu_u_prio7_DW = 3;
	// removed localparam type sv2v_uu_u_prio7_d
	localparam [2:0] sv2v_uu_u_prio7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio7_we),
		.wd(prio7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio7_ext_d_0),
		.qe(),
		.q(reg2hw[246-:3]),
		.qs(prio7_qs)
	);
	// Trace: design.sv:94610:3
	localparam signed [31:0] sv2v_uu_u_prio8_DW = 3;
	// removed localparam type sv2v_uu_u_prio8_d
	localparam [2:0] sv2v_uu_u_prio8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio8_we),
		.wd(prio8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio8_ext_d_0),
		.qe(),
		.q(reg2hw[243-:3]),
		.qs(prio8_qs)
	);
	// Trace: design.sv:94637:3
	localparam signed [31:0] sv2v_uu_u_prio9_DW = 3;
	// removed localparam type sv2v_uu_u_prio9_d
	localparam [2:0] sv2v_uu_u_prio9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio9_we),
		.wd(prio9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio9_ext_d_0),
		.qe(),
		.q(reg2hw[240-:3]),
		.qs(prio9_qs)
	);
	// Trace: design.sv:94664:3
	localparam signed [31:0] sv2v_uu_u_prio10_DW = 3;
	// removed localparam type sv2v_uu_u_prio10_d
	localparam [2:0] sv2v_uu_u_prio10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio10_we),
		.wd(prio10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio10_ext_d_0),
		.qe(),
		.q(reg2hw[237-:3]),
		.qs(prio10_qs)
	);
	// Trace: design.sv:94691:3
	localparam signed [31:0] sv2v_uu_u_prio11_DW = 3;
	// removed localparam type sv2v_uu_u_prio11_d
	localparam [2:0] sv2v_uu_u_prio11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio11_we),
		.wd(prio11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio11_ext_d_0),
		.qe(),
		.q(reg2hw[234-:3]),
		.qs(prio11_qs)
	);
	// Trace: design.sv:94718:3
	localparam signed [31:0] sv2v_uu_u_prio12_DW = 3;
	// removed localparam type sv2v_uu_u_prio12_d
	localparam [2:0] sv2v_uu_u_prio12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio12_we),
		.wd(prio12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio12_ext_d_0),
		.qe(),
		.q(reg2hw[231-:3]),
		.qs(prio12_qs)
	);
	// Trace: design.sv:94745:3
	localparam signed [31:0] sv2v_uu_u_prio13_DW = 3;
	// removed localparam type sv2v_uu_u_prio13_d
	localparam [2:0] sv2v_uu_u_prio13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio13_we),
		.wd(prio13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio13_ext_d_0),
		.qe(),
		.q(reg2hw[228-:3]),
		.qs(prio13_qs)
	);
	// Trace: design.sv:94772:3
	localparam signed [31:0] sv2v_uu_u_prio14_DW = 3;
	// removed localparam type sv2v_uu_u_prio14_d
	localparam [2:0] sv2v_uu_u_prio14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio14_we),
		.wd(prio14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio14_ext_d_0),
		.qe(),
		.q(reg2hw[225-:3]),
		.qs(prio14_qs)
	);
	// Trace: design.sv:94799:3
	localparam signed [31:0] sv2v_uu_u_prio15_DW = 3;
	// removed localparam type sv2v_uu_u_prio15_d
	localparam [2:0] sv2v_uu_u_prio15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio15_we),
		.wd(prio15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio15_ext_d_0),
		.qe(),
		.q(reg2hw[222-:3]),
		.qs(prio15_qs)
	);
	// Trace: design.sv:94826:3
	localparam signed [31:0] sv2v_uu_u_prio16_DW = 3;
	// removed localparam type sv2v_uu_u_prio16_d
	localparam [2:0] sv2v_uu_u_prio16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio16_we),
		.wd(prio16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio16_ext_d_0),
		.qe(),
		.q(reg2hw[219-:3]),
		.qs(prio16_qs)
	);
	// Trace: design.sv:94853:3
	localparam signed [31:0] sv2v_uu_u_prio17_DW = 3;
	// removed localparam type sv2v_uu_u_prio17_d
	localparam [2:0] sv2v_uu_u_prio17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio17_we),
		.wd(prio17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio17_ext_d_0),
		.qe(),
		.q(reg2hw[216-:3]),
		.qs(prio17_qs)
	);
	// Trace: design.sv:94880:3
	localparam signed [31:0] sv2v_uu_u_prio18_DW = 3;
	// removed localparam type sv2v_uu_u_prio18_d
	localparam [2:0] sv2v_uu_u_prio18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio18_we),
		.wd(prio18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio18_ext_d_0),
		.qe(),
		.q(reg2hw[213-:3]),
		.qs(prio18_qs)
	);
	// Trace: design.sv:94907:3
	localparam signed [31:0] sv2v_uu_u_prio19_DW = 3;
	// removed localparam type sv2v_uu_u_prio19_d
	localparam [2:0] sv2v_uu_u_prio19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio19_we),
		.wd(prio19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio19_ext_d_0),
		.qe(),
		.q(reg2hw[210-:3]),
		.qs(prio19_qs)
	);
	// Trace: design.sv:94934:3
	localparam signed [31:0] sv2v_uu_u_prio20_DW = 3;
	// removed localparam type sv2v_uu_u_prio20_d
	localparam [2:0] sv2v_uu_u_prio20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio20_we),
		.wd(prio20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio20_ext_d_0),
		.qe(),
		.q(reg2hw[207-:3]),
		.qs(prio20_qs)
	);
	// Trace: design.sv:94961:3
	localparam signed [31:0] sv2v_uu_u_prio21_DW = 3;
	// removed localparam type sv2v_uu_u_prio21_d
	localparam [2:0] sv2v_uu_u_prio21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio21_we),
		.wd(prio21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio21_ext_d_0),
		.qe(),
		.q(reg2hw[204-:3]),
		.qs(prio21_qs)
	);
	// Trace: design.sv:94988:3
	localparam signed [31:0] sv2v_uu_u_prio22_DW = 3;
	// removed localparam type sv2v_uu_u_prio22_d
	localparam [2:0] sv2v_uu_u_prio22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio22_we),
		.wd(prio22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio22_ext_d_0),
		.qe(),
		.q(reg2hw[201-:3]),
		.qs(prio22_qs)
	);
	// Trace: design.sv:95015:3
	localparam signed [31:0] sv2v_uu_u_prio23_DW = 3;
	// removed localparam type sv2v_uu_u_prio23_d
	localparam [2:0] sv2v_uu_u_prio23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio23_we),
		.wd(prio23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio23_ext_d_0),
		.qe(),
		.q(reg2hw[198-:3]),
		.qs(prio23_qs)
	);
	// Trace: design.sv:95042:3
	localparam signed [31:0] sv2v_uu_u_prio24_DW = 3;
	// removed localparam type sv2v_uu_u_prio24_d
	localparam [2:0] sv2v_uu_u_prio24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio24_we),
		.wd(prio24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio24_ext_d_0),
		.qe(),
		.q(reg2hw[195-:3]),
		.qs(prio24_qs)
	);
	// Trace: design.sv:95069:3
	localparam signed [31:0] sv2v_uu_u_prio25_DW = 3;
	// removed localparam type sv2v_uu_u_prio25_d
	localparam [2:0] sv2v_uu_u_prio25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio25_we),
		.wd(prio25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio25_ext_d_0),
		.qe(),
		.q(reg2hw[192-:3]),
		.qs(prio25_qs)
	);
	// Trace: design.sv:95096:3
	localparam signed [31:0] sv2v_uu_u_prio26_DW = 3;
	// removed localparam type sv2v_uu_u_prio26_d
	localparam [2:0] sv2v_uu_u_prio26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio26_we),
		.wd(prio26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio26_ext_d_0),
		.qe(),
		.q(reg2hw[189-:3]),
		.qs(prio26_qs)
	);
	// Trace: design.sv:95123:3
	localparam signed [31:0] sv2v_uu_u_prio27_DW = 3;
	// removed localparam type sv2v_uu_u_prio27_d
	localparam [2:0] sv2v_uu_u_prio27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio27_we),
		.wd(prio27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio27_ext_d_0),
		.qe(),
		.q(reg2hw[186-:3]),
		.qs(prio27_qs)
	);
	// Trace: design.sv:95150:3
	localparam signed [31:0] sv2v_uu_u_prio28_DW = 3;
	// removed localparam type sv2v_uu_u_prio28_d
	localparam [2:0] sv2v_uu_u_prio28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio28_we),
		.wd(prio28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio28_ext_d_0),
		.qe(),
		.q(reg2hw[183-:3]),
		.qs(prio28_qs)
	);
	// Trace: design.sv:95177:3
	localparam signed [31:0] sv2v_uu_u_prio29_DW = 3;
	// removed localparam type sv2v_uu_u_prio29_d
	localparam [2:0] sv2v_uu_u_prio29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio29_we),
		.wd(prio29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio29_ext_d_0),
		.qe(),
		.q(reg2hw[180-:3]),
		.qs(prio29_qs)
	);
	// Trace: design.sv:95204:3
	localparam signed [31:0] sv2v_uu_u_prio30_DW = 3;
	// removed localparam type sv2v_uu_u_prio30_d
	localparam [2:0] sv2v_uu_u_prio30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio30_we),
		.wd(prio30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio30_ext_d_0),
		.qe(),
		.q(reg2hw[177-:3]),
		.qs(prio30_qs)
	);
	// Trace: design.sv:95231:3
	localparam signed [31:0] sv2v_uu_u_prio31_DW = 3;
	// removed localparam type sv2v_uu_u_prio31_d
	localparam [2:0] sv2v_uu_u_prio31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio31_we),
		.wd(prio31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio31_ext_d_0),
		.qe(),
		.q(reg2hw[174-:3]),
		.qs(prio31_qs)
	);
	// Trace: design.sv:95258:3
	localparam signed [31:0] sv2v_uu_u_prio32_DW = 3;
	// removed localparam type sv2v_uu_u_prio32_d
	localparam [2:0] sv2v_uu_u_prio32_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio32(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio32_we),
		.wd(prio32_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio32_ext_d_0),
		.qe(),
		.q(reg2hw[171-:3]),
		.qs(prio32_qs)
	);
	// Trace: design.sv:95285:3
	localparam signed [31:0] sv2v_uu_u_prio33_DW = 3;
	// removed localparam type sv2v_uu_u_prio33_d
	localparam [2:0] sv2v_uu_u_prio33_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio33(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio33_we),
		.wd(prio33_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio33_ext_d_0),
		.qe(),
		.q(reg2hw[168-:3]),
		.qs(prio33_qs)
	);
	// Trace: design.sv:95312:3
	localparam signed [31:0] sv2v_uu_u_prio34_DW = 3;
	// removed localparam type sv2v_uu_u_prio34_d
	localparam [2:0] sv2v_uu_u_prio34_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio34(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio34_we),
		.wd(prio34_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio34_ext_d_0),
		.qe(),
		.q(reg2hw[165-:3]),
		.qs(prio34_qs)
	);
	// Trace: design.sv:95339:3
	localparam signed [31:0] sv2v_uu_u_prio35_DW = 3;
	// removed localparam type sv2v_uu_u_prio35_d
	localparam [2:0] sv2v_uu_u_prio35_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio35(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio35_we),
		.wd(prio35_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio35_ext_d_0),
		.qe(),
		.q(reg2hw[162-:3]),
		.qs(prio35_qs)
	);
	// Trace: design.sv:95366:3
	localparam signed [31:0] sv2v_uu_u_prio36_DW = 3;
	// removed localparam type sv2v_uu_u_prio36_d
	localparam [2:0] sv2v_uu_u_prio36_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio36(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio36_we),
		.wd(prio36_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio36_ext_d_0),
		.qe(),
		.q(reg2hw[159-:3]),
		.qs(prio36_qs)
	);
	// Trace: design.sv:95393:3
	localparam signed [31:0] sv2v_uu_u_prio37_DW = 3;
	// removed localparam type sv2v_uu_u_prio37_d
	localparam [2:0] sv2v_uu_u_prio37_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio37(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio37_we),
		.wd(prio37_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio37_ext_d_0),
		.qe(),
		.q(reg2hw[156-:3]),
		.qs(prio37_qs)
	);
	// Trace: design.sv:95420:3
	localparam signed [31:0] sv2v_uu_u_prio38_DW = 3;
	// removed localparam type sv2v_uu_u_prio38_d
	localparam [2:0] sv2v_uu_u_prio38_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio38(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio38_we),
		.wd(prio38_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio38_ext_d_0),
		.qe(),
		.q(reg2hw[153-:3]),
		.qs(prio38_qs)
	);
	// Trace: design.sv:95447:3
	localparam signed [31:0] sv2v_uu_u_prio39_DW = 3;
	// removed localparam type sv2v_uu_u_prio39_d
	localparam [2:0] sv2v_uu_u_prio39_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio39(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio39_we),
		.wd(prio39_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio39_ext_d_0),
		.qe(),
		.q(reg2hw[150-:3]),
		.qs(prio39_qs)
	);
	// Trace: design.sv:95474:3
	localparam signed [31:0] sv2v_uu_u_prio40_DW = 3;
	// removed localparam type sv2v_uu_u_prio40_d
	localparam [2:0] sv2v_uu_u_prio40_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio40(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio40_we),
		.wd(prio40_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio40_ext_d_0),
		.qe(),
		.q(reg2hw[147-:3]),
		.qs(prio40_qs)
	);
	// Trace: design.sv:95501:3
	localparam signed [31:0] sv2v_uu_u_prio41_DW = 3;
	// removed localparam type sv2v_uu_u_prio41_d
	localparam [2:0] sv2v_uu_u_prio41_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio41(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio41_we),
		.wd(prio41_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio41_ext_d_0),
		.qe(),
		.q(reg2hw[144-:3]),
		.qs(prio41_qs)
	);
	// Trace: design.sv:95528:3
	localparam signed [31:0] sv2v_uu_u_prio42_DW = 3;
	// removed localparam type sv2v_uu_u_prio42_d
	localparam [2:0] sv2v_uu_u_prio42_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio42(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio42_we),
		.wd(prio42_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio42_ext_d_0),
		.qe(),
		.q(reg2hw[141-:3]),
		.qs(prio42_qs)
	);
	// Trace: design.sv:95555:3
	localparam signed [31:0] sv2v_uu_u_prio43_DW = 3;
	// removed localparam type sv2v_uu_u_prio43_d
	localparam [2:0] sv2v_uu_u_prio43_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio43(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio43_we),
		.wd(prio43_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio43_ext_d_0),
		.qe(),
		.q(reg2hw[138-:3]),
		.qs(prio43_qs)
	);
	// Trace: design.sv:95582:3
	localparam signed [31:0] sv2v_uu_u_prio44_DW = 3;
	// removed localparam type sv2v_uu_u_prio44_d
	localparam [2:0] sv2v_uu_u_prio44_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio44(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio44_we),
		.wd(prio44_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio44_ext_d_0),
		.qe(),
		.q(reg2hw[135-:3]),
		.qs(prio44_qs)
	);
	// Trace: design.sv:95609:3
	localparam signed [31:0] sv2v_uu_u_prio45_DW = 3;
	// removed localparam type sv2v_uu_u_prio45_d
	localparam [2:0] sv2v_uu_u_prio45_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio45(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio45_we),
		.wd(prio45_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio45_ext_d_0),
		.qe(),
		.q(reg2hw[132-:3]),
		.qs(prio45_qs)
	);
	// Trace: design.sv:95636:3
	localparam signed [31:0] sv2v_uu_u_prio46_DW = 3;
	// removed localparam type sv2v_uu_u_prio46_d
	localparam [2:0] sv2v_uu_u_prio46_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio46(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio46_we),
		.wd(prio46_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio46_ext_d_0),
		.qe(),
		.q(reg2hw[129-:3]),
		.qs(prio46_qs)
	);
	// Trace: design.sv:95663:3
	localparam signed [31:0] sv2v_uu_u_prio47_DW = 3;
	// removed localparam type sv2v_uu_u_prio47_d
	localparam [2:0] sv2v_uu_u_prio47_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio47(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio47_we),
		.wd(prio47_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio47_ext_d_0),
		.qe(),
		.q(reg2hw[126-:3]),
		.qs(prio47_qs)
	);
	// Trace: design.sv:95690:3
	localparam signed [31:0] sv2v_uu_u_prio48_DW = 3;
	// removed localparam type sv2v_uu_u_prio48_d
	localparam [2:0] sv2v_uu_u_prio48_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio48(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio48_we),
		.wd(prio48_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio48_ext_d_0),
		.qe(),
		.q(reg2hw[123-:3]),
		.qs(prio48_qs)
	);
	// Trace: design.sv:95717:3
	localparam signed [31:0] sv2v_uu_u_prio49_DW = 3;
	// removed localparam type sv2v_uu_u_prio49_d
	localparam [2:0] sv2v_uu_u_prio49_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio49(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio49_we),
		.wd(prio49_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio49_ext_d_0),
		.qe(),
		.q(reg2hw[120-:3]),
		.qs(prio49_qs)
	);
	// Trace: design.sv:95744:3
	localparam signed [31:0] sv2v_uu_u_prio50_DW = 3;
	// removed localparam type sv2v_uu_u_prio50_d
	localparam [2:0] sv2v_uu_u_prio50_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio50(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio50_we),
		.wd(prio50_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio50_ext_d_0),
		.qe(),
		.q(reg2hw[117-:3]),
		.qs(prio50_qs)
	);
	// Trace: design.sv:95771:3
	localparam signed [31:0] sv2v_uu_u_prio51_DW = 3;
	// removed localparam type sv2v_uu_u_prio51_d
	localparam [2:0] sv2v_uu_u_prio51_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio51(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio51_we),
		.wd(prio51_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio51_ext_d_0),
		.qe(),
		.q(reg2hw[114-:3]),
		.qs(prio51_qs)
	);
	// Trace: design.sv:95798:3
	localparam signed [31:0] sv2v_uu_u_prio52_DW = 3;
	// removed localparam type sv2v_uu_u_prio52_d
	localparam [2:0] sv2v_uu_u_prio52_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio52(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio52_we),
		.wd(prio52_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio52_ext_d_0),
		.qe(),
		.q(reg2hw[111-:3]),
		.qs(prio52_qs)
	);
	// Trace: design.sv:95825:3
	localparam signed [31:0] sv2v_uu_u_prio53_DW = 3;
	// removed localparam type sv2v_uu_u_prio53_d
	localparam [2:0] sv2v_uu_u_prio53_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio53(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio53_we),
		.wd(prio53_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio53_ext_d_0),
		.qe(),
		.q(reg2hw[108-:3]),
		.qs(prio53_qs)
	);
	// Trace: design.sv:95852:3
	localparam signed [31:0] sv2v_uu_u_prio54_DW = 3;
	// removed localparam type sv2v_uu_u_prio54_d
	localparam [2:0] sv2v_uu_u_prio54_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio54(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio54_we),
		.wd(prio54_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio54_ext_d_0),
		.qe(),
		.q(reg2hw[105-:3]),
		.qs(prio54_qs)
	);
	// Trace: design.sv:95879:3
	localparam signed [31:0] sv2v_uu_u_prio55_DW = 3;
	// removed localparam type sv2v_uu_u_prio55_d
	localparam [2:0] sv2v_uu_u_prio55_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio55(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio55_we),
		.wd(prio55_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio55_ext_d_0),
		.qe(),
		.q(reg2hw[102-:3]),
		.qs(prio55_qs)
	);
	// Trace: design.sv:95906:3
	localparam signed [31:0] sv2v_uu_u_prio56_DW = 3;
	// removed localparam type sv2v_uu_u_prio56_d
	localparam [2:0] sv2v_uu_u_prio56_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio56(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio56_we),
		.wd(prio56_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio56_ext_d_0),
		.qe(),
		.q(reg2hw[99-:3]),
		.qs(prio56_qs)
	);
	// Trace: design.sv:95933:3
	localparam signed [31:0] sv2v_uu_u_prio57_DW = 3;
	// removed localparam type sv2v_uu_u_prio57_d
	localparam [2:0] sv2v_uu_u_prio57_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio57(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio57_we),
		.wd(prio57_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio57_ext_d_0),
		.qe(),
		.q(reg2hw[96-:3]),
		.qs(prio57_qs)
	);
	// Trace: design.sv:95960:3
	localparam signed [31:0] sv2v_uu_u_prio58_DW = 3;
	// removed localparam type sv2v_uu_u_prio58_d
	localparam [2:0] sv2v_uu_u_prio58_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio58(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio58_we),
		.wd(prio58_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio58_ext_d_0),
		.qe(),
		.q(reg2hw[93-:3]),
		.qs(prio58_qs)
	);
	// Trace: design.sv:95987:3
	localparam signed [31:0] sv2v_uu_u_prio59_DW = 3;
	// removed localparam type sv2v_uu_u_prio59_d
	localparam [2:0] sv2v_uu_u_prio59_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio59(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio59_we),
		.wd(prio59_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio59_ext_d_0),
		.qe(),
		.q(reg2hw[90-:3]),
		.qs(prio59_qs)
	);
	// Trace: design.sv:96014:3
	localparam signed [31:0] sv2v_uu_u_prio60_DW = 3;
	// removed localparam type sv2v_uu_u_prio60_d
	localparam [2:0] sv2v_uu_u_prio60_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio60(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio60_we),
		.wd(prio60_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio60_ext_d_0),
		.qe(),
		.q(reg2hw[87-:3]),
		.qs(prio60_qs)
	);
	// Trace: design.sv:96041:3
	localparam signed [31:0] sv2v_uu_u_prio61_DW = 3;
	// removed localparam type sv2v_uu_u_prio61_d
	localparam [2:0] sv2v_uu_u_prio61_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio61(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio61_we),
		.wd(prio61_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio61_ext_d_0),
		.qe(),
		.q(reg2hw[84-:3]),
		.qs(prio61_qs)
	);
	// Trace: design.sv:96068:3
	localparam signed [31:0] sv2v_uu_u_prio62_DW = 3;
	// removed localparam type sv2v_uu_u_prio62_d
	localparam [2:0] sv2v_uu_u_prio62_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio62(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio62_we),
		.wd(prio62_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio62_ext_d_0),
		.qe(),
		.q(reg2hw[81-:3]),
		.qs(prio62_qs)
	);
	// Trace: design.sv:96095:3
	localparam signed [31:0] sv2v_uu_u_prio63_DW = 3;
	// removed localparam type sv2v_uu_u_prio63_d
	localparam [2:0] sv2v_uu_u_prio63_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_prio63(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(prio63_we),
		.wd(prio63_wd),
		.de(1'b0),
		.d(sv2v_uu_u_prio63_ext_d_0),
		.qe(),
		.q(reg2hw[78-:3]),
		.qs(prio63_qs)
	);
	// Trace: design.sv:96125:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_0_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_0_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_0_we),
		.wd(ie0_0_e_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_0_ext_d_0),
		.qe(),
		.q(reg2hw[12]),
		.qs(ie0_0_e_0_qs)
	);
	// Trace: design.sv:96151:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_1_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_1_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_1_we),
		.wd(ie0_0_e_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_1_ext_d_0),
		.qe(),
		.q(reg2hw[13]),
		.qs(ie0_0_e_1_qs)
	);
	// Trace: design.sv:96177:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_2_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_2_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_2_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_2_we),
		.wd(ie0_0_e_2_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_2_ext_d_0),
		.qe(),
		.q(reg2hw[14]),
		.qs(ie0_0_e_2_qs)
	);
	// Trace: design.sv:96203:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_3_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_3_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_3_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_3_we),
		.wd(ie0_0_e_3_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_3_ext_d_0),
		.qe(),
		.q(reg2hw[15]),
		.qs(ie0_0_e_3_qs)
	);
	// Trace: design.sv:96229:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_4_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_4_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_4_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_4_we),
		.wd(ie0_0_e_4_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_4_ext_d_0),
		.qe(),
		.q(reg2hw[16]),
		.qs(ie0_0_e_4_qs)
	);
	// Trace: design.sv:96255:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_5_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_5_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_5_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_5_we),
		.wd(ie0_0_e_5_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_5_ext_d_0),
		.qe(),
		.q(reg2hw[17]),
		.qs(ie0_0_e_5_qs)
	);
	// Trace: design.sv:96281:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_6_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_6_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_6_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_6_we),
		.wd(ie0_0_e_6_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_6_ext_d_0),
		.qe(),
		.q(reg2hw[18]),
		.qs(ie0_0_e_6_qs)
	);
	// Trace: design.sv:96307:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_7_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_7_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_7_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_7_we),
		.wd(ie0_0_e_7_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_7_ext_d_0),
		.qe(),
		.q(reg2hw[19]),
		.qs(ie0_0_e_7_qs)
	);
	// Trace: design.sv:96333:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_8_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_8_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_8_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_8_we),
		.wd(ie0_0_e_8_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_8_ext_d_0),
		.qe(),
		.q(reg2hw[20]),
		.qs(ie0_0_e_8_qs)
	);
	// Trace: design.sv:96359:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_9_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_9_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_9_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_9_we),
		.wd(ie0_0_e_9_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_9_ext_d_0),
		.qe(),
		.q(reg2hw[21]),
		.qs(ie0_0_e_9_qs)
	);
	// Trace: design.sv:96385:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_10_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_10_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_10_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_10_we),
		.wd(ie0_0_e_10_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_10_ext_d_0),
		.qe(),
		.q(reg2hw[22]),
		.qs(ie0_0_e_10_qs)
	);
	// Trace: design.sv:96411:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_11_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_11_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_11_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_11_we),
		.wd(ie0_0_e_11_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_11_ext_d_0),
		.qe(),
		.q(reg2hw[23]),
		.qs(ie0_0_e_11_qs)
	);
	// Trace: design.sv:96437:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_12_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_12_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_12_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_12_we),
		.wd(ie0_0_e_12_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_12_ext_d_0),
		.qe(),
		.q(reg2hw[24]),
		.qs(ie0_0_e_12_qs)
	);
	// Trace: design.sv:96463:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_13_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_13_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_13_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_13_we),
		.wd(ie0_0_e_13_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_13_ext_d_0),
		.qe(),
		.q(reg2hw[25]),
		.qs(ie0_0_e_13_qs)
	);
	// Trace: design.sv:96489:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_14_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_14_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_14_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_14_we),
		.wd(ie0_0_e_14_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_14_ext_d_0),
		.qe(),
		.q(reg2hw[26]),
		.qs(ie0_0_e_14_qs)
	);
	// Trace: design.sv:96515:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_15_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_15_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_15_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_15_we),
		.wd(ie0_0_e_15_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_15_ext_d_0),
		.qe(),
		.q(reg2hw[27]),
		.qs(ie0_0_e_15_qs)
	);
	// Trace: design.sv:96541:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_16_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_16_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_16_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_16_we),
		.wd(ie0_0_e_16_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_16_ext_d_0),
		.qe(),
		.q(reg2hw[28]),
		.qs(ie0_0_e_16_qs)
	);
	// Trace: design.sv:96567:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_17_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_17_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_17_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_17_we),
		.wd(ie0_0_e_17_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_17_ext_d_0),
		.qe(),
		.q(reg2hw[29]),
		.qs(ie0_0_e_17_qs)
	);
	// Trace: design.sv:96593:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_18_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_18_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_18_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_18_we),
		.wd(ie0_0_e_18_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_18_ext_d_0),
		.qe(),
		.q(reg2hw[30]),
		.qs(ie0_0_e_18_qs)
	);
	// Trace: design.sv:96619:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_19_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_19_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_19_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_19_we),
		.wd(ie0_0_e_19_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_19_ext_d_0),
		.qe(),
		.q(reg2hw[31]),
		.qs(ie0_0_e_19_qs)
	);
	// Trace: design.sv:96645:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_20_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_20_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_20_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_20_we),
		.wd(ie0_0_e_20_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_20_ext_d_0),
		.qe(),
		.q(reg2hw[32]),
		.qs(ie0_0_e_20_qs)
	);
	// Trace: design.sv:96671:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_21_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_21_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_21_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_21_we),
		.wd(ie0_0_e_21_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_21_ext_d_0),
		.qe(),
		.q(reg2hw[33]),
		.qs(ie0_0_e_21_qs)
	);
	// Trace: design.sv:96697:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_22_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_22_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_22_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_22_we),
		.wd(ie0_0_e_22_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_22_ext_d_0),
		.qe(),
		.q(reg2hw[34]),
		.qs(ie0_0_e_22_qs)
	);
	// Trace: design.sv:96723:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_23_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_23_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_23_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_23_we),
		.wd(ie0_0_e_23_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_23_ext_d_0),
		.qe(),
		.q(reg2hw[35]),
		.qs(ie0_0_e_23_qs)
	);
	// Trace: design.sv:96749:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_24_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_24_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_24_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_24_we),
		.wd(ie0_0_e_24_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_24_ext_d_0),
		.qe(),
		.q(reg2hw[36]),
		.qs(ie0_0_e_24_qs)
	);
	// Trace: design.sv:96775:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_25_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_25_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_25_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_25_we),
		.wd(ie0_0_e_25_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_25_ext_d_0),
		.qe(),
		.q(reg2hw[37]),
		.qs(ie0_0_e_25_qs)
	);
	// Trace: design.sv:96801:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_26_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_26_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_26_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_26_we),
		.wd(ie0_0_e_26_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_26_ext_d_0),
		.qe(),
		.q(reg2hw[38]),
		.qs(ie0_0_e_26_qs)
	);
	// Trace: design.sv:96827:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_27_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_27_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_27_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_27_we),
		.wd(ie0_0_e_27_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_27_ext_d_0),
		.qe(),
		.q(reg2hw[39]),
		.qs(ie0_0_e_27_qs)
	);
	// Trace: design.sv:96853:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_28_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_28_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_28_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_28_we),
		.wd(ie0_0_e_28_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_28_ext_d_0),
		.qe(),
		.q(reg2hw[40]),
		.qs(ie0_0_e_28_qs)
	);
	// Trace: design.sv:96879:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_29_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_29_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_29_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_29_we),
		.wd(ie0_0_e_29_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_29_ext_d_0),
		.qe(),
		.q(reg2hw[41]),
		.qs(ie0_0_e_29_qs)
	);
	// Trace: design.sv:96905:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_30_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_30_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_30_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_30_we),
		.wd(ie0_0_e_30_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_30_ext_d_0),
		.qe(),
		.q(reg2hw[42]),
		.qs(ie0_0_e_30_qs)
	);
	// Trace: design.sv:96931:3
	localparam signed [31:0] sv2v_uu_u_ie0_0_e_31_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_0_e_31_d
	localparam [0:0] sv2v_uu_u_ie0_0_e_31_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_0_e_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_0_e_31_we),
		.wd(ie0_0_e_31_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_0_e_31_ext_d_0),
		.qe(),
		.q(reg2hw[43]),
		.qs(ie0_0_e_31_qs)
	);
	// Trace: design.sv:96960:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_32_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_32_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_32_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_32(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_32_we),
		.wd(ie0_1_e_32_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_32_ext_d_0),
		.qe(),
		.q(reg2hw[44]),
		.qs(ie0_1_e_32_qs)
	);
	// Trace: design.sv:96986:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_33_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_33_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_33_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_33(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_33_we),
		.wd(ie0_1_e_33_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_33_ext_d_0),
		.qe(),
		.q(reg2hw[45]),
		.qs(ie0_1_e_33_qs)
	);
	// Trace: design.sv:97012:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_34_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_34_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_34_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_34(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_34_we),
		.wd(ie0_1_e_34_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_34_ext_d_0),
		.qe(),
		.q(reg2hw[46]),
		.qs(ie0_1_e_34_qs)
	);
	// Trace: design.sv:97038:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_35_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_35_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_35_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_35(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_35_we),
		.wd(ie0_1_e_35_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_35_ext_d_0),
		.qe(),
		.q(reg2hw[47]),
		.qs(ie0_1_e_35_qs)
	);
	// Trace: design.sv:97064:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_36_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_36_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_36_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_36(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_36_we),
		.wd(ie0_1_e_36_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_36_ext_d_0),
		.qe(),
		.q(reg2hw[48]),
		.qs(ie0_1_e_36_qs)
	);
	// Trace: design.sv:97090:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_37_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_37_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_37_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_37(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_37_we),
		.wd(ie0_1_e_37_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_37_ext_d_0),
		.qe(),
		.q(reg2hw[49]),
		.qs(ie0_1_e_37_qs)
	);
	// Trace: design.sv:97116:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_38_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_38_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_38_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_38(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_38_we),
		.wd(ie0_1_e_38_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_38_ext_d_0),
		.qe(),
		.q(reg2hw[50]),
		.qs(ie0_1_e_38_qs)
	);
	// Trace: design.sv:97142:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_39_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_39_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_39_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_39(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_39_we),
		.wd(ie0_1_e_39_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_39_ext_d_0),
		.qe(),
		.q(reg2hw[51]),
		.qs(ie0_1_e_39_qs)
	);
	// Trace: design.sv:97168:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_40_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_40_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_40_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_40(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_40_we),
		.wd(ie0_1_e_40_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_40_ext_d_0),
		.qe(),
		.q(reg2hw[52]),
		.qs(ie0_1_e_40_qs)
	);
	// Trace: design.sv:97194:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_41_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_41_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_41_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_41(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_41_we),
		.wd(ie0_1_e_41_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_41_ext_d_0),
		.qe(),
		.q(reg2hw[53]),
		.qs(ie0_1_e_41_qs)
	);
	// Trace: design.sv:97220:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_42_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_42_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_42_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_42(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_42_we),
		.wd(ie0_1_e_42_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_42_ext_d_0),
		.qe(),
		.q(reg2hw[54]),
		.qs(ie0_1_e_42_qs)
	);
	// Trace: design.sv:97246:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_43_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_43_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_43_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_43(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_43_we),
		.wd(ie0_1_e_43_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_43_ext_d_0),
		.qe(),
		.q(reg2hw[55]),
		.qs(ie0_1_e_43_qs)
	);
	// Trace: design.sv:97272:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_44_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_44_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_44_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_44(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_44_we),
		.wd(ie0_1_e_44_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_44_ext_d_0),
		.qe(),
		.q(reg2hw[56]),
		.qs(ie0_1_e_44_qs)
	);
	// Trace: design.sv:97298:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_45_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_45_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_45_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_45(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_45_we),
		.wd(ie0_1_e_45_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_45_ext_d_0),
		.qe(),
		.q(reg2hw[57]),
		.qs(ie0_1_e_45_qs)
	);
	// Trace: design.sv:97324:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_46_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_46_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_46_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_46(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_46_we),
		.wd(ie0_1_e_46_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_46_ext_d_0),
		.qe(),
		.q(reg2hw[58]),
		.qs(ie0_1_e_46_qs)
	);
	// Trace: design.sv:97350:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_47_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_47_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_47_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_47(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_47_we),
		.wd(ie0_1_e_47_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_47_ext_d_0),
		.qe(),
		.q(reg2hw[59]),
		.qs(ie0_1_e_47_qs)
	);
	// Trace: design.sv:97376:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_48_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_48_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_48_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_48(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_48_we),
		.wd(ie0_1_e_48_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_48_ext_d_0),
		.qe(),
		.q(reg2hw[60]),
		.qs(ie0_1_e_48_qs)
	);
	// Trace: design.sv:97402:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_49_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_49_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_49_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_49(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_49_we),
		.wd(ie0_1_e_49_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_49_ext_d_0),
		.qe(),
		.q(reg2hw[61]),
		.qs(ie0_1_e_49_qs)
	);
	// Trace: design.sv:97428:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_50_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_50_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_50_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_50(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_50_we),
		.wd(ie0_1_e_50_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_50_ext_d_0),
		.qe(),
		.q(reg2hw[62]),
		.qs(ie0_1_e_50_qs)
	);
	// Trace: design.sv:97454:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_51_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_51_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_51_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_51(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_51_we),
		.wd(ie0_1_e_51_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_51_ext_d_0),
		.qe(),
		.q(reg2hw[63]),
		.qs(ie0_1_e_51_qs)
	);
	// Trace: design.sv:97480:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_52_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_52_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_52_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_52(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_52_we),
		.wd(ie0_1_e_52_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_52_ext_d_0),
		.qe(),
		.q(reg2hw[64]),
		.qs(ie0_1_e_52_qs)
	);
	// Trace: design.sv:97506:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_53_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_53_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_53_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_53(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_53_we),
		.wd(ie0_1_e_53_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_53_ext_d_0),
		.qe(),
		.q(reg2hw[65]),
		.qs(ie0_1_e_53_qs)
	);
	// Trace: design.sv:97532:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_54_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_54_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_54_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_54(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_54_we),
		.wd(ie0_1_e_54_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_54_ext_d_0),
		.qe(),
		.q(reg2hw[66]),
		.qs(ie0_1_e_54_qs)
	);
	// Trace: design.sv:97558:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_55_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_55_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_55_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_55(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_55_we),
		.wd(ie0_1_e_55_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_55_ext_d_0),
		.qe(),
		.q(reg2hw[67]),
		.qs(ie0_1_e_55_qs)
	);
	// Trace: design.sv:97584:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_56_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_56_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_56_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_56(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_56_we),
		.wd(ie0_1_e_56_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_56_ext_d_0),
		.qe(),
		.q(reg2hw[68]),
		.qs(ie0_1_e_56_qs)
	);
	// Trace: design.sv:97610:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_57_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_57_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_57_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_57(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_57_we),
		.wd(ie0_1_e_57_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_57_ext_d_0),
		.qe(),
		.q(reg2hw[69]),
		.qs(ie0_1_e_57_qs)
	);
	// Trace: design.sv:97636:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_58_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_58_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_58_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_58(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_58_we),
		.wd(ie0_1_e_58_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_58_ext_d_0),
		.qe(),
		.q(reg2hw[70]),
		.qs(ie0_1_e_58_qs)
	);
	// Trace: design.sv:97662:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_59_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_59_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_59_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_59(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_59_we),
		.wd(ie0_1_e_59_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_59_ext_d_0),
		.qe(),
		.q(reg2hw[71]),
		.qs(ie0_1_e_59_qs)
	);
	// Trace: design.sv:97688:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_60_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_60_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_60_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_60(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_60_we),
		.wd(ie0_1_e_60_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_60_ext_d_0),
		.qe(),
		.q(reg2hw[72]),
		.qs(ie0_1_e_60_qs)
	);
	// Trace: design.sv:97714:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_61_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_61_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_61_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_61(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_61_we),
		.wd(ie0_1_e_61_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_61_ext_d_0),
		.qe(),
		.q(reg2hw[73]),
		.qs(ie0_1_e_61_qs)
	);
	// Trace: design.sv:97740:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_62_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_62_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_62_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_62(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_62_we),
		.wd(ie0_1_e_62_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_62_ext_d_0),
		.qe(),
		.q(reg2hw[74]),
		.qs(ie0_1_e_62_qs)
	);
	// Trace: design.sv:97766:3
	localparam signed [31:0] sv2v_uu_u_ie0_1_e_63_DW = 1;
	// removed localparam type sv2v_uu_u_ie0_1_e_63_d
	localparam [0:0] sv2v_uu_u_ie0_1_e_63_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ie0_1_e_63(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ie0_1_e_63_we),
		.wd(ie0_1_e_63_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ie0_1_e_63_ext_d_0),
		.qe(),
		.q(reg2hw[75]),
		.qs(ie0_1_e_63_qs)
	);
	// Trace: design.sv:97794:3
	localparam signed [31:0] sv2v_uu_u_threshold0_DW = 3;
	// removed localparam type sv2v_uu_u_threshold0_d
	localparam [2:0] sv2v_uu_u_threshold0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_threshold0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(threshold0_we),
		.wd(threshold0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_threshold0_ext_d_0),
		.qe(),
		.q(reg2hw[11-:3]),
		.qs(threshold0_qs)
	);
	// Trace: design.sv:97821:3
	prim_subreg_ext #(.DW(6)) u_cc0(
		.re(cc0_re),
		.we(cc0_we),
		.wd(cc0_wd),
		.d(hw2reg[5-:6]),
		.qre(reg2hw[1]),
		.qe(reg2hw[2]),
		.q(reg2hw[8-:6]),
		.qs(cc0_qs)
	);
	// Trace: design.sv:97837:3
	localparam signed [31:0] sv2v_uu_u_msip0_DW = 1;
	// removed localparam type sv2v_uu_u_msip0_d
	localparam [0:0] sv2v_uu_u_msip0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_msip0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(msip0_we),
		.wd(msip0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_msip0_ext_d_0),
		.qe(),
		.q(reg2hw[-0]),
		.qs(msip0_qs)
	);
	// Trace: design.sv:97864:3
	reg [72:0] addr_hit;
	// Trace: design.sv:97865:3
	localparam signed [31:0] rv_plic_reg_pkg_BlockAw = 10;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_CC0_OFFSET = 10'h20c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_IE0_0_OFFSET = 10'h200;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_IE0_1_OFFSET = 10'h204;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_IP_0_OFFSET = 10'h000;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_IP_1_OFFSET = 10'h004;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_LE_0_OFFSET = 10'h008;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_LE_1_OFFSET = 10'h00c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_MSIP0_OFFSET = 10'h210;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO0_OFFSET = 10'h010;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO10_OFFSET = 10'h038;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO11_OFFSET = 10'h03c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO12_OFFSET = 10'h040;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO13_OFFSET = 10'h044;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO14_OFFSET = 10'h048;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO15_OFFSET = 10'h04c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO16_OFFSET = 10'h050;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO17_OFFSET = 10'h054;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO18_OFFSET = 10'h058;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO19_OFFSET = 10'h05c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO1_OFFSET = 10'h014;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO20_OFFSET = 10'h060;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO21_OFFSET = 10'h064;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO22_OFFSET = 10'h068;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO23_OFFSET = 10'h06c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO24_OFFSET = 10'h070;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO25_OFFSET = 10'h074;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO26_OFFSET = 10'h078;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO27_OFFSET = 10'h07c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO28_OFFSET = 10'h080;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO29_OFFSET = 10'h084;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO2_OFFSET = 10'h018;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO30_OFFSET = 10'h088;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO31_OFFSET = 10'h08c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO32_OFFSET = 10'h090;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO33_OFFSET = 10'h094;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO34_OFFSET = 10'h098;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO35_OFFSET = 10'h09c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO36_OFFSET = 10'h0a0;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO37_OFFSET = 10'h0a4;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO38_OFFSET = 10'h0a8;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO39_OFFSET = 10'h0ac;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO3_OFFSET = 10'h01c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO40_OFFSET = 10'h0b0;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO41_OFFSET = 10'h0b4;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO42_OFFSET = 10'h0b8;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO43_OFFSET = 10'h0bc;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO44_OFFSET = 10'h0c0;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO45_OFFSET = 10'h0c4;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO46_OFFSET = 10'h0c8;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO47_OFFSET = 10'h0cc;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO48_OFFSET = 10'h0d0;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO49_OFFSET = 10'h0d4;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO4_OFFSET = 10'h020;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO50_OFFSET = 10'h0d8;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO51_OFFSET = 10'h0dc;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO52_OFFSET = 10'h0e0;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO53_OFFSET = 10'h0e4;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO54_OFFSET = 10'h0e8;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO55_OFFSET = 10'h0ec;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO56_OFFSET = 10'h0f0;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO57_OFFSET = 10'h0f4;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO58_OFFSET = 10'h0f8;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO59_OFFSET = 10'h0fc;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO5_OFFSET = 10'h024;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO60_OFFSET = 10'h100;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO61_OFFSET = 10'h104;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO62_OFFSET = 10'h108;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO63_OFFSET = 10'h10c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO6_OFFSET = 10'h028;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO7_OFFSET = 10'h02c;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO8_OFFSET = 10'h030;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_PRIO9_OFFSET = 10'h034;
	localparam [9:0] rv_plic_reg_pkg_RV_PLIC_THRESHOLD0_OFFSET = 10'h208;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:97866:5
		addr_hit = 1'sb0;
		// Trace: design.sv:97867:5
		addr_hit[0] = reg_addr == rv_plic_reg_pkg_RV_PLIC_IP_0_OFFSET;
		// Trace: design.sv:97868:5
		addr_hit[1] = reg_addr == rv_plic_reg_pkg_RV_PLIC_IP_1_OFFSET;
		// Trace: design.sv:97869:5
		addr_hit[2] = reg_addr == rv_plic_reg_pkg_RV_PLIC_LE_0_OFFSET;
		// Trace: design.sv:97870:5
		addr_hit[3] = reg_addr == rv_plic_reg_pkg_RV_PLIC_LE_1_OFFSET;
		// Trace: design.sv:97871:5
		addr_hit[4] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO0_OFFSET;
		// Trace: design.sv:97872:5
		addr_hit[5] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO1_OFFSET;
		// Trace: design.sv:97873:5
		addr_hit[6] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO2_OFFSET;
		// Trace: design.sv:97874:5
		addr_hit[7] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO3_OFFSET;
		// Trace: design.sv:97875:5
		addr_hit[8] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO4_OFFSET;
		// Trace: design.sv:97876:5
		addr_hit[9] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO5_OFFSET;
		// Trace: design.sv:97877:5
		addr_hit[10] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO6_OFFSET;
		// Trace: design.sv:97878:5
		addr_hit[11] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO7_OFFSET;
		// Trace: design.sv:97879:5
		addr_hit[12] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO8_OFFSET;
		// Trace: design.sv:97880:5
		addr_hit[13] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO9_OFFSET;
		// Trace: design.sv:97881:5
		addr_hit[14] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO10_OFFSET;
		// Trace: design.sv:97882:5
		addr_hit[15] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO11_OFFSET;
		// Trace: design.sv:97883:5
		addr_hit[16] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO12_OFFSET;
		// Trace: design.sv:97884:5
		addr_hit[17] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO13_OFFSET;
		// Trace: design.sv:97885:5
		addr_hit[18] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO14_OFFSET;
		// Trace: design.sv:97886:5
		addr_hit[19] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO15_OFFSET;
		// Trace: design.sv:97887:5
		addr_hit[20] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO16_OFFSET;
		// Trace: design.sv:97888:5
		addr_hit[21] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO17_OFFSET;
		// Trace: design.sv:97889:5
		addr_hit[22] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO18_OFFSET;
		// Trace: design.sv:97890:5
		addr_hit[23] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO19_OFFSET;
		// Trace: design.sv:97891:5
		addr_hit[24] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO20_OFFSET;
		// Trace: design.sv:97892:5
		addr_hit[25] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO21_OFFSET;
		// Trace: design.sv:97893:5
		addr_hit[26] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO22_OFFSET;
		// Trace: design.sv:97894:5
		addr_hit[27] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO23_OFFSET;
		// Trace: design.sv:97895:5
		addr_hit[28] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO24_OFFSET;
		// Trace: design.sv:97896:5
		addr_hit[29] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO25_OFFSET;
		// Trace: design.sv:97897:5
		addr_hit[30] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO26_OFFSET;
		// Trace: design.sv:97898:5
		addr_hit[31] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO27_OFFSET;
		// Trace: design.sv:97899:5
		addr_hit[32] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO28_OFFSET;
		// Trace: design.sv:97900:5
		addr_hit[33] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO29_OFFSET;
		// Trace: design.sv:97901:5
		addr_hit[34] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO30_OFFSET;
		// Trace: design.sv:97902:5
		addr_hit[35] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO31_OFFSET;
		// Trace: design.sv:97903:5
		addr_hit[36] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO32_OFFSET;
		// Trace: design.sv:97904:5
		addr_hit[37] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO33_OFFSET;
		// Trace: design.sv:97905:5
		addr_hit[38] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO34_OFFSET;
		// Trace: design.sv:97906:5
		addr_hit[39] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO35_OFFSET;
		// Trace: design.sv:97907:5
		addr_hit[40] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO36_OFFSET;
		// Trace: design.sv:97908:5
		addr_hit[41] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO37_OFFSET;
		// Trace: design.sv:97909:5
		addr_hit[42] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO38_OFFSET;
		// Trace: design.sv:97910:5
		addr_hit[43] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO39_OFFSET;
		// Trace: design.sv:97911:5
		addr_hit[44] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO40_OFFSET;
		// Trace: design.sv:97912:5
		addr_hit[45] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO41_OFFSET;
		// Trace: design.sv:97913:5
		addr_hit[46] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO42_OFFSET;
		// Trace: design.sv:97914:5
		addr_hit[47] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO43_OFFSET;
		// Trace: design.sv:97915:5
		addr_hit[48] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO44_OFFSET;
		// Trace: design.sv:97916:5
		addr_hit[49] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO45_OFFSET;
		// Trace: design.sv:97917:5
		addr_hit[50] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO46_OFFSET;
		// Trace: design.sv:97918:5
		addr_hit[51] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO47_OFFSET;
		// Trace: design.sv:97919:5
		addr_hit[52] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO48_OFFSET;
		// Trace: design.sv:97920:5
		addr_hit[53] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO49_OFFSET;
		// Trace: design.sv:97921:5
		addr_hit[54] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO50_OFFSET;
		// Trace: design.sv:97922:5
		addr_hit[55] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO51_OFFSET;
		// Trace: design.sv:97923:5
		addr_hit[56] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO52_OFFSET;
		// Trace: design.sv:97924:5
		addr_hit[57] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO53_OFFSET;
		// Trace: design.sv:97925:5
		addr_hit[58] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO54_OFFSET;
		// Trace: design.sv:97926:5
		addr_hit[59] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO55_OFFSET;
		// Trace: design.sv:97927:5
		addr_hit[60] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO56_OFFSET;
		// Trace: design.sv:97928:5
		addr_hit[61] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO57_OFFSET;
		// Trace: design.sv:97929:5
		addr_hit[62] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO58_OFFSET;
		// Trace: design.sv:97930:5
		addr_hit[63] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO59_OFFSET;
		// Trace: design.sv:97931:5
		addr_hit[64] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO60_OFFSET;
		// Trace: design.sv:97932:5
		addr_hit[65] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO61_OFFSET;
		// Trace: design.sv:97933:5
		addr_hit[66] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO62_OFFSET;
		// Trace: design.sv:97934:5
		addr_hit[67] = reg_addr == rv_plic_reg_pkg_RV_PLIC_PRIO63_OFFSET;
		// Trace: design.sv:97935:5
		addr_hit[68] = reg_addr == rv_plic_reg_pkg_RV_PLIC_IE0_0_OFFSET;
		// Trace: design.sv:97936:5
		addr_hit[69] = reg_addr == rv_plic_reg_pkg_RV_PLIC_IE0_1_OFFSET;
		// Trace: design.sv:97937:5
		addr_hit[70] = reg_addr == rv_plic_reg_pkg_RV_PLIC_THRESHOLD0_OFFSET;
		// Trace: design.sv:97938:5
		addr_hit[71] = reg_addr == rv_plic_reg_pkg_RV_PLIC_CC0_OFFSET;
		// Trace: design.sv:97939:5
		addr_hit[72] = reg_addr == rv_plic_reg_pkg_RV_PLIC_MSIP0_OFFSET;
	end
	// Trace: design.sv:97942:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:97945:3
	localparam [291:0] rv_plic_reg_pkg_RV_PLIC_PERMIT = 292'b1111111111111111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000111111111000100010001;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:97946:5
		wr_err = reg_we & (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((addr_hit[0] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[288+:4] & ~reg_be)) | (addr_hit[1] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[284+:4] & ~reg_be))) | (addr_hit[2] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[280+:4] & ~reg_be))) | (addr_hit[3] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[276+:4] & ~reg_be))) | (addr_hit[4] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[272+:4] & ~reg_be))) | (addr_hit[5] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[268+:4] & ~reg_be))) | (addr_hit[6] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[264+:4] & ~reg_be))) | (addr_hit[7] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[260+:4] & ~reg_be))) | (addr_hit[8] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[256+:4] & ~reg_be))) | (addr_hit[9] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[252+:4] & ~reg_be))) | (addr_hit[10] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[248+:4] & ~reg_be))) | (addr_hit[11] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[244+:4] & ~reg_be))) | (addr_hit[12] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[240+:4] & ~reg_be))) | (addr_hit[13] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[236+:4] & ~reg_be))) | (addr_hit[14] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[232+:4] & ~reg_be))) | (addr_hit[15] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[228+:4] & ~reg_be))) | (addr_hit[16] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[224+:4] & ~reg_be))) | (addr_hit[17] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[220+:4] & ~reg_be))) | (addr_hit[18] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[216+:4] & ~reg_be))) | (addr_hit[19] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[212+:4] & ~reg_be))) | (addr_hit[20] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[208+:4] & ~reg_be))) | (addr_hit[21] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[204+:4] & ~reg_be))) | (addr_hit[22] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[200+:4] & ~reg_be))) | (addr_hit[23] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[196+:4] & ~reg_be))) | (addr_hit[24] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[192+:4] & ~reg_be))) | (addr_hit[25] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[188+:4] & ~reg_be))) | (addr_hit[26] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[184+:4] & ~reg_be))) | (addr_hit[27] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[180+:4] & ~reg_be))) | (addr_hit[28] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[176+:4] & ~reg_be))) | (addr_hit[29] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[172+:4] & ~reg_be))) | (addr_hit[30] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[168+:4] & ~reg_be))) | (addr_hit[31] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[164+:4] & ~reg_be))) | (addr_hit[32] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[160+:4] & ~reg_be))) | (addr_hit[33] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[156+:4] & ~reg_be))) | (addr_hit[34] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[152+:4] & ~reg_be))) | (addr_hit[35] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[148+:4] & ~reg_be))) | (addr_hit[36] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[144+:4] & ~reg_be))) | (addr_hit[37] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[140+:4] & ~reg_be))) | (addr_hit[38] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[136+:4] & ~reg_be))) | (addr_hit[39] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[132+:4] & ~reg_be))) | (addr_hit[40] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[128+:4] & ~reg_be))) | (addr_hit[41] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[124+:4] & ~reg_be))) | (addr_hit[42] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[120+:4] & ~reg_be))) | (addr_hit[43] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[116+:4] & ~reg_be))) | (addr_hit[44] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[112+:4] & ~reg_be))) | (addr_hit[45] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[108+:4] & ~reg_be))) | (addr_hit[46] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[104+:4] & ~reg_be))) | (addr_hit[47] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[100+:4] & ~reg_be))) | (addr_hit[48] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[96+:4] & ~reg_be))) | (addr_hit[49] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[92+:4] & ~reg_be))) | (addr_hit[50] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[88+:4] & ~reg_be))) | (addr_hit[51] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[84+:4] & ~reg_be))) | (addr_hit[52] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[80+:4] & ~reg_be))) | (addr_hit[53] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[76+:4] & ~reg_be))) | (addr_hit[54] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[72+:4] & ~reg_be))) | (addr_hit[55] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[68+:4] & ~reg_be))) | (addr_hit[56] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[64+:4] & ~reg_be))) | (addr_hit[57] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[60+:4] & ~reg_be))) | (addr_hit[58] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[56+:4] & ~reg_be))) | (addr_hit[59] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[52+:4] & ~reg_be))) | (addr_hit[60] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[48+:4] & ~reg_be))) | (addr_hit[61] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[44+:4] & ~reg_be))) | (addr_hit[62] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[40+:4] & ~reg_be))) | (addr_hit[63] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[36+:4] & ~reg_be))) | (addr_hit[64] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[32+:4] & ~reg_be))) | (addr_hit[65] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[28+:4] & ~reg_be))) | (addr_hit[66] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[24+:4] & ~reg_be))) | (addr_hit[67] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[20+:4] & ~reg_be))) | (addr_hit[68] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[16+:4] & ~reg_be))) | (addr_hit[69] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[12+:4] & ~reg_be))) | (addr_hit[70] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[8+:4] & ~reg_be))) | (addr_hit[71] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[4+:4] & ~reg_be))) | (addr_hit[72] & |(rv_plic_reg_pkg_RV_PLIC_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:98022:3
	assign le_0_le_0_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98023:3
	assign le_0_le_0_wd = reg_wdata[0];
	// Trace: design.sv:98025:3
	assign le_0_le_1_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98026:3
	assign le_0_le_1_wd = reg_wdata[1];
	// Trace: design.sv:98028:3
	assign le_0_le_2_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98029:3
	assign le_0_le_2_wd = reg_wdata[2];
	// Trace: design.sv:98031:3
	assign le_0_le_3_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98032:3
	assign le_0_le_3_wd = reg_wdata[3];
	// Trace: design.sv:98034:3
	assign le_0_le_4_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98035:3
	assign le_0_le_4_wd = reg_wdata[4];
	// Trace: design.sv:98037:3
	assign le_0_le_5_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98038:3
	assign le_0_le_5_wd = reg_wdata[5];
	// Trace: design.sv:98040:3
	assign le_0_le_6_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98041:3
	assign le_0_le_6_wd = reg_wdata[6];
	// Trace: design.sv:98043:3
	assign le_0_le_7_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98044:3
	assign le_0_le_7_wd = reg_wdata[7];
	// Trace: design.sv:98046:3
	assign le_0_le_8_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98047:3
	assign le_0_le_8_wd = reg_wdata[8];
	// Trace: design.sv:98049:3
	assign le_0_le_9_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98050:3
	assign le_0_le_9_wd = reg_wdata[9];
	// Trace: design.sv:98052:3
	assign le_0_le_10_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98053:3
	assign le_0_le_10_wd = reg_wdata[10];
	// Trace: design.sv:98055:3
	assign le_0_le_11_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98056:3
	assign le_0_le_11_wd = reg_wdata[11];
	// Trace: design.sv:98058:3
	assign le_0_le_12_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98059:3
	assign le_0_le_12_wd = reg_wdata[12];
	// Trace: design.sv:98061:3
	assign le_0_le_13_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98062:3
	assign le_0_le_13_wd = reg_wdata[13];
	// Trace: design.sv:98064:3
	assign le_0_le_14_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98065:3
	assign le_0_le_14_wd = reg_wdata[14];
	// Trace: design.sv:98067:3
	assign le_0_le_15_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98068:3
	assign le_0_le_15_wd = reg_wdata[15];
	// Trace: design.sv:98070:3
	assign le_0_le_16_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98071:3
	assign le_0_le_16_wd = reg_wdata[16];
	// Trace: design.sv:98073:3
	assign le_0_le_17_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98074:3
	assign le_0_le_17_wd = reg_wdata[17];
	// Trace: design.sv:98076:3
	assign le_0_le_18_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98077:3
	assign le_0_le_18_wd = reg_wdata[18];
	// Trace: design.sv:98079:3
	assign le_0_le_19_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98080:3
	assign le_0_le_19_wd = reg_wdata[19];
	// Trace: design.sv:98082:3
	assign le_0_le_20_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98083:3
	assign le_0_le_20_wd = reg_wdata[20];
	// Trace: design.sv:98085:3
	assign le_0_le_21_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98086:3
	assign le_0_le_21_wd = reg_wdata[21];
	// Trace: design.sv:98088:3
	assign le_0_le_22_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98089:3
	assign le_0_le_22_wd = reg_wdata[22];
	// Trace: design.sv:98091:3
	assign le_0_le_23_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98092:3
	assign le_0_le_23_wd = reg_wdata[23];
	// Trace: design.sv:98094:3
	assign le_0_le_24_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98095:3
	assign le_0_le_24_wd = reg_wdata[24];
	// Trace: design.sv:98097:3
	assign le_0_le_25_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98098:3
	assign le_0_le_25_wd = reg_wdata[25];
	// Trace: design.sv:98100:3
	assign le_0_le_26_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98101:3
	assign le_0_le_26_wd = reg_wdata[26];
	// Trace: design.sv:98103:3
	assign le_0_le_27_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98104:3
	assign le_0_le_27_wd = reg_wdata[27];
	// Trace: design.sv:98106:3
	assign le_0_le_28_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98107:3
	assign le_0_le_28_wd = reg_wdata[28];
	// Trace: design.sv:98109:3
	assign le_0_le_29_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98110:3
	assign le_0_le_29_wd = reg_wdata[29];
	// Trace: design.sv:98112:3
	assign le_0_le_30_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98113:3
	assign le_0_le_30_wd = reg_wdata[30];
	// Trace: design.sv:98115:3
	assign le_0_le_31_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:98116:3
	assign le_0_le_31_wd = reg_wdata[31];
	// Trace: design.sv:98118:3
	assign le_1_le_32_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98119:3
	assign le_1_le_32_wd = reg_wdata[0];
	// Trace: design.sv:98121:3
	assign le_1_le_33_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98122:3
	assign le_1_le_33_wd = reg_wdata[1];
	// Trace: design.sv:98124:3
	assign le_1_le_34_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98125:3
	assign le_1_le_34_wd = reg_wdata[2];
	// Trace: design.sv:98127:3
	assign le_1_le_35_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98128:3
	assign le_1_le_35_wd = reg_wdata[3];
	// Trace: design.sv:98130:3
	assign le_1_le_36_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98131:3
	assign le_1_le_36_wd = reg_wdata[4];
	// Trace: design.sv:98133:3
	assign le_1_le_37_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98134:3
	assign le_1_le_37_wd = reg_wdata[5];
	// Trace: design.sv:98136:3
	assign le_1_le_38_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98137:3
	assign le_1_le_38_wd = reg_wdata[6];
	// Trace: design.sv:98139:3
	assign le_1_le_39_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98140:3
	assign le_1_le_39_wd = reg_wdata[7];
	// Trace: design.sv:98142:3
	assign le_1_le_40_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98143:3
	assign le_1_le_40_wd = reg_wdata[8];
	// Trace: design.sv:98145:3
	assign le_1_le_41_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98146:3
	assign le_1_le_41_wd = reg_wdata[9];
	// Trace: design.sv:98148:3
	assign le_1_le_42_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98149:3
	assign le_1_le_42_wd = reg_wdata[10];
	// Trace: design.sv:98151:3
	assign le_1_le_43_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98152:3
	assign le_1_le_43_wd = reg_wdata[11];
	// Trace: design.sv:98154:3
	assign le_1_le_44_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98155:3
	assign le_1_le_44_wd = reg_wdata[12];
	// Trace: design.sv:98157:3
	assign le_1_le_45_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98158:3
	assign le_1_le_45_wd = reg_wdata[13];
	// Trace: design.sv:98160:3
	assign le_1_le_46_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98161:3
	assign le_1_le_46_wd = reg_wdata[14];
	// Trace: design.sv:98163:3
	assign le_1_le_47_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98164:3
	assign le_1_le_47_wd = reg_wdata[15];
	// Trace: design.sv:98166:3
	assign le_1_le_48_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98167:3
	assign le_1_le_48_wd = reg_wdata[16];
	// Trace: design.sv:98169:3
	assign le_1_le_49_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98170:3
	assign le_1_le_49_wd = reg_wdata[17];
	// Trace: design.sv:98172:3
	assign le_1_le_50_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98173:3
	assign le_1_le_50_wd = reg_wdata[18];
	// Trace: design.sv:98175:3
	assign le_1_le_51_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98176:3
	assign le_1_le_51_wd = reg_wdata[19];
	// Trace: design.sv:98178:3
	assign le_1_le_52_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98179:3
	assign le_1_le_52_wd = reg_wdata[20];
	// Trace: design.sv:98181:3
	assign le_1_le_53_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98182:3
	assign le_1_le_53_wd = reg_wdata[21];
	// Trace: design.sv:98184:3
	assign le_1_le_54_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98185:3
	assign le_1_le_54_wd = reg_wdata[22];
	// Trace: design.sv:98187:3
	assign le_1_le_55_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98188:3
	assign le_1_le_55_wd = reg_wdata[23];
	// Trace: design.sv:98190:3
	assign le_1_le_56_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98191:3
	assign le_1_le_56_wd = reg_wdata[24];
	// Trace: design.sv:98193:3
	assign le_1_le_57_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98194:3
	assign le_1_le_57_wd = reg_wdata[25];
	// Trace: design.sv:98196:3
	assign le_1_le_58_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98197:3
	assign le_1_le_58_wd = reg_wdata[26];
	// Trace: design.sv:98199:3
	assign le_1_le_59_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98200:3
	assign le_1_le_59_wd = reg_wdata[27];
	// Trace: design.sv:98202:3
	assign le_1_le_60_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98203:3
	assign le_1_le_60_wd = reg_wdata[28];
	// Trace: design.sv:98205:3
	assign le_1_le_61_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98206:3
	assign le_1_le_61_wd = reg_wdata[29];
	// Trace: design.sv:98208:3
	assign le_1_le_62_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98209:3
	assign le_1_le_62_wd = reg_wdata[30];
	// Trace: design.sv:98211:3
	assign le_1_le_63_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:98212:3
	assign le_1_le_63_wd = reg_wdata[31];
	// Trace: design.sv:98214:3
	assign prio0_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:98215:3
	assign prio0_wd = reg_wdata[2:0];
	// Trace: design.sv:98217:3
	assign prio1_we = (addr_hit[5] & reg_we) & !reg_error;
	// Trace: design.sv:98218:3
	assign prio1_wd = reg_wdata[2:0];
	// Trace: design.sv:98220:3
	assign prio2_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:98221:3
	assign prio2_wd = reg_wdata[2:0];
	// Trace: design.sv:98223:3
	assign prio3_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:98224:3
	assign prio3_wd = reg_wdata[2:0];
	// Trace: design.sv:98226:3
	assign prio4_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:98227:3
	assign prio4_wd = reg_wdata[2:0];
	// Trace: design.sv:98229:3
	assign prio5_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:98230:3
	assign prio5_wd = reg_wdata[2:0];
	// Trace: design.sv:98232:3
	assign prio6_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:98233:3
	assign prio6_wd = reg_wdata[2:0];
	// Trace: design.sv:98235:3
	assign prio7_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:98236:3
	assign prio7_wd = reg_wdata[2:0];
	// Trace: design.sv:98238:3
	assign prio8_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:98239:3
	assign prio8_wd = reg_wdata[2:0];
	// Trace: design.sv:98241:3
	assign prio9_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:98242:3
	assign prio9_wd = reg_wdata[2:0];
	// Trace: design.sv:98244:3
	assign prio10_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:98245:3
	assign prio10_wd = reg_wdata[2:0];
	// Trace: design.sv:98247:3
	assign prio11_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:98248:3
	assign prio11_wd = reg_wdata[2:0];
	// Trace: design.sv:98250:3
	assign prio12_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:98251:3
	assign prio12_wd = reg_wdata[2:0];
	// Trace: design.sv:98253:3
	assign prio13_we = (addr_hit[17] & reg_we) & !reg_error;
	// Trace: design.sv:98254:3
	assign prio13_wd = reg_wdata[2:0];
	// Trace: design.sv:98256:3
	assign prio14_we = (addr_hit[18] & reg_we) & !reg_error;
	// Trace: design.sv:98257:3
	assign prio14_wd = reg_wdata[2:0];
	// Trace: design.sv:98259:3
	assign prio15_we = (addr_hit[19] & reg_we) & !reg_error;
	// Trace: design.sv:98260:3
	assign prio15_wd = reg_wdata[2:0];
	// Trace: design.sv:98262:3
	assign prio16_we = (addr_hit[20] & reg_we) & !reg_error;
	// Trace: design.sv:98263:3
	assign prio16_wd = reg_wdata[2:0];
	// Trace: design.sv:98265:3
	assign prio17_we = (addr_hit[21] & reg_we) & !reg_error;
	// Trace: design.sv:98266:3
	assign prio17_wd = reg_wdata[2:0];
	// Trace: design.sv:98268:3
	assign prio18_we = (addr_hit[22] & reg_we) & !reg_error;
	// Trace: design.sv:98269:3
	assign prio18_wd = reg_wdata[2:0];
	// Trace: design.sv:98271:3
	assign prio19_we = (addr_hit[23] & reg_we) & !reg_error;
	// Trace: design.sv:98272:3
	assign prio19_wd = reg_wdata[2:0];
	// Trace: design.sv:98274:3
	assign prio20_we = (addr_hit[24] & reg_we) & !reg_error;
	// Trace: design.sv:98275:3
	assign prio20_wd = reg_wdata[2:0];
	// Trace: design.sv:98277:3
	assign prio21_we = (addr_hit[25] & reg_we) & !reg_error;
	// Trace: design.sv:98278:3
	assign prio21_wd = reg_wdata[2:0];
	// Trace: design.sv:98280:3
	assign prio22_we = (addr_hit[26] & reg_we) & !reg_error;
	// Trace: design.sv:98281:3
	assign prio22_wd = reg_wdata[2:0];
	// Trace: design.sv:98283:3
	assign prio23_we = (addr_hit[27] & reg_we) & !reg_error;
	// Trace: design.sv:98284:3
	assign prio23_wd = reg_wdata[2:0];
	// Trace: design.sv:98286:3
	assign prio24_we = (addr_hit[28] & reg_we) & !reg_error;
	// Trace: design.sv:98287:3
	assign prio24_wd = reg_wdata[2:0];
	// Trace: design.sv:98289:3
	assign prio25_we = (addr_hit[29] & reg_we) & !reg_error;
	// Trace: design.sv:98290:3
	assign prio25_wd = reg_wdata[2:0];
	// Trace: design.sv:98292:3
	assign prio26_we = (addr_hit[30] & reg_we) & !reg_error;
	// Trace: design.sv:98293:3
	assign prio26_wd = reg_wdata[2:0];
	// Trace: design.sv:98295:3
	assign prio27_we = (addr_hit[31] & reg_we) & !reg_error;
	// Trace: design.sv:98296:3
	assign prio27_wd = reg_wdata[2:0];
	// Trace: design.sv:98298:3
	assign prio28_we = (addr_hit[32] & reg_we) & !reg_error;
	// Trace: design.sv:98299:3
	assign prio28_wd = reg_wdata[2:0];
	// Trace: design.sv:98301:3
	assign prio29_we = (addr_hit[33] & reg_we) & !reg_error;
	// Trace: design.sv:98302:3
	assign prio29_wd = reg_wdata[2:0];
	// Trace: design.sv:98304:3
	assign prio30_we = (addr_hit[34] & reg_we) & !reg_error;
	// Trace: design.sv:98305:3
	assign prio30_wd = reg_wdata[2:0];
	// Trace: design.sv:98307:3
	assign prio31_we = (addr_hit[35] & reg_we) & !reg_error;
	// Trace: design.sv:98308:3
	assign prio31_wd = reg_wdata[2:0];
	// Trace: design.sv:98310:3
	assign prio32_we = (addr_hit[36] & reg_we) & !reg_error;
	// Trace: design.sv:98311:3
	assign prio32_wd = reg_wdata[2:0];
	// Trace: design.sv:98313:3
	assign prio33_we = (addr_hit[37] & reg_we) & !reg_error;
	// Trace: design.sv:98314:3
	assign prio33_wd = reg_wdata[2:0];
	// Trace: design.sv:98316:3
	assign prio34_we = (addr_hit[38] & reg_we) & !reg_error;
	// Trace: design.sv:98317:3
	assign prio34_wd = reg_wdata[2:0];
	// Trace: design.sv:98319:3
	assign prio35_we = (addr_hit[39] & reg_we) & !reg_error;
	// Trace: design.sv:98320:3
	assign prio35_wd = reg_wdata[2:0];
	// Trace: design.sv:98322:3
	assign prio36_we = (addr_hit[40] & reg_we) & !reg_error;
	// Trace: design.sv:98323:3
	assign prio36_wd = reg_wdata[2:0];
	// Trace: design.sv:98325:3
	assign prio37_we = (addr_hit[41] & reg_we) & !reg_error;
	// Trace: design.sv:98326:3
	assign prio37_wd = reg_wdata[2:0];
	// Trace: design.sv:98328:3
	assign prio38_we = (addr_hit[42] & reg_we) & !reg_error;
	// Trace: design.sv:98329:3
	assign prio38_wd = reg_wdata[2:0];
	// Trace: design.sv:98331:3
	assign prio39_we = (addr_hit[43] & reg_we) & !reg_error;
	// Trace: design.sv:98332:3
	assign prio39_wd = reg_wdata[2:0];
	// Trace: design.sv:98334:3
	assign prio40_we = (addr_hit[44] & reg_we) & !reg_error;
	// Trace: design.sv:98335:3
	assign prio40_wd = reg_wdata[2:0];
	// Trace: design.sv:98337:3
	assign prio41_we = (addr_hit[45] & reg_we) & !reg_error;
	// Trace: design.sv:98338:3
	assign prio41_wd = reg_wdata[2:0];
	// Trace: design.sv:98340:3
	assign prio42_we = (addr_hit[46] & reg_we) & !reg_error;
	// Trace: design.sv:98341:3
	assign prio42_wd = reg_wdata[2:0];
	// Trace: design.sv:98343:3
	assign prio43_we = (addr_hit[47] & reg_we) & !reg_error;
	// Trace: design.sv:98344:3
	assign prio43_wd = reg_wdata[2:0];
	// Trace: design.sv:98346:3
	assign prio44_we = (addr_hit[48] & reg_we) & !reg_error;
	// Trace: design.sv:98347:3
	assign prio44_wd = reg_wdata[2:0];
	// Trace: design.sv:98349:3
	assign prio45_we = (addr_hit[49] & reg_we) & !reg_error;
	// Trace: design.sv:98350:3
	assign prio45_wd = reg_wdata[2:0];
	// Trace: design.sv:98352:3
	assign prio46_we = (addr_hit[50] & reg_we) & !reg_error;
	// Trace: design.sv:98353:3
	assign prio46_wd = reg_wdata[2:0];
	// Trace: design.sv:98355:3
	assign prio47_we = (addr_hit[51] & reg_we) & !reg_error;
	// Trace: design.sv:98356:3
	assign prio47_wd = reg_wdata[2:0];
	// Trace: design.sv:98358:3
	assign prio48_we = (addr_hit[52] & reg_we) & !reg_error;
	// Trace: design.sv:98359:3
	assign prio48_wd = reg_wdata[2:0];
	// Trace: design.sv:98361:3
	assign prio49_we = (addr_hit[53] & reg_we) & !reg_error;
	// Trace: design.sv:98362:3
	assign prio49_wd = reg_wdata[2:0];
	// Trace: design.sv:98364:3
	assign prio50_we = (addr_hit[54] & reg_we) & !reg_error;
	// Trace: design.sv:98365:3
	assign prio50_wd = reg_wdata[2:0];
	// Trace: design.sv:98367:3
	assign prio51_we = (addr_hit[55] & reg_we) & !reg_error;
	// Trace: design.sv:98368:3
	assign prio51_wd = reg_wdata[2:0];
	// Trace: design.sv:98370:3
	assign prio52_we = (addr_hit[56] & reg_we) & !reg_error;
	// Trace: design.sv:98371:3
	assign prio52_wd = reg_wdata[2:0];
	// Trace: design.sv:98373:3
	assign prio53_we = (addr_hit[57] & reg_we) & !reg_error;
	// Trace: design.sv:98374:3
	assign prio53_wd = reg_wdata[2:0];
	// Trace: design.sv:98376:3
	assign prio54_we = (addr_hit[58] & reg_we) & !reg_error;
	// Trace: design.sv:98377:3
	assign prio54_wd = reg_wdata[2:0];
	// Trace: design.sv:98379:3
	assign prio55_we = (addr_hit[59] & reg_we) & !reg_error;
	// Trace: design.sv:98380:3
	assign prio55_wd = reg_wdata[2:0];
	// Trace: design.sv:98382:3
	assign prio56_we = (addr_hit[60] & reg_we) & !reg_error;
	// Trace: design.sv:98383:3
	assign prio56_wd = reg_wdata[2:0];
	// Trace: design.sv:98385:3
	assign prio57_we = (addr_hit[61] & reg_we) & !reg_error;
	// Trace: design.sv:98386:3
	assign prio57_wd = reg_wdata[2:0];
	// Trace: design.sv:98388:3
	assign prio58_we = (addr_hit[62] & reg_we) & !reg_error;
	// Trace: design.sv:98389:3
	assign prio58_wd = reg_wdata[2:0];
	// Trace: design.sv:98391:3
	assign prio59_we = (addr_hit[63] & reg_we) & !reg_error;
	// Trace: design.sv:98392:3
	assign prio59_wd = reg_wdata[2:0];
	// Trace: design.sv:98394:3
	assign prio60_we = (addr_hit[64] & reg_we) & !reg_error;
	// Trace: design.sv:98395:3
	assign prio60_wd = reg_wdata[2:0];
	// Trace: design.sv:98397:3
	assign prio61_we = (addr_hit[65] & reg_we) & !reg_error;
	// Trace: design.sv:98398:3
	assign prio61_wd = reg_wdata[2:0];
	// Trace: design.sv:98400:3
	assign prio62_we = (addr_hit[66] & reg_we) & !reg_error;
	// Trace: design.sv:98401:3
	assign prio62_wd = reg_wdata[2:0];
	// Trace: design.sv:98403:3
	assign prio63_we = (addr_hit[67] & reg_we) & !reg_error;
	// Trace: design.sv:98404:3
	assign prio63_wd = reg_wdata[2:0];
	// Trace: design.sv:98406:3
	assign ie0_0_e_0_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98407:3
	assign ie0_0_e_0_wd = reg_wdata[0];
	// Trace: design.sv:98409:3
	assign ie0_0_e_1_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98410:3
	assign ie0_0_e_1_wd = reg_wdata[1];
	// Trace: design.sv:98412:3
	assign ie0_0_e_2_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98413:3
	assign ie0_0_e_2_wd = reg_wdata[2];
	// Trace: design.sv:98415:3
	assign ie0_0_e_3_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98416:3
	assign ie0_0_e_3_wd = reg_wdata[3];
	// Trace: design.sv:98418:3
	assign ie0_0_e_4_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98419:3
	assign ie0_0_e_4_wd = reg_wdata[4];
	// Trace: design.sv:98421:3
	assign ie0_0_e_5_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98422:3
	assign ie0_0_e_5_wd = reg_wdata[5];
	// Trace: design.sv:98424:3
	assign ie0_0_e_6_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98425:3
	assign ie0_0_e_6_wd = reg_wdata[6];
	// Trace: design.sv:98427:3
	assign ie0_0_e_7_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98428:3
	assign ie0_0_e_7_wd = reg_wdata[7];
	// Trace: design.sv:98430:3
	assign ie0_0_e_8_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98431:3
	assign ie0_0_e_8_wd = reg_wdata[8];
	// Trace: design.sv:98433:3
	assign ie0_0_e_9_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98434:3
	assign ie0_0_e_9_wd = reg_wdata[9];
	// Trace: design.sv:98436:3
	assign ie0_0_e_10_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98437:3
	assign ie0_0_e_10_wd = reg_wdata[10];
	// Trace: design.sv:98439:3
	assign ie0_0_e_11_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98440:3
	assign ie0_0_e_11_wd = reg_wdata[11];
	// Trace: design.sv:98442:3
	assign ie0_0_e_12_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98443:3
	assign ie0_0_e_12_wd = reg_wdata[12];
	// Trace: design.sv:98445:3
	assign ie0_0_e_13_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98446:3
	assign ie0_0_e_13_wd = reg_wdata[13];
	// Trace: design.sv:98448:3
	assign ie0_0_e_14_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98449:3
	assign ie0_0_e_14_wd = reg_wdata[14];
	// Trace: design.sv:98451:3
	assign ie0_0_e_15_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98452:3
	assign ie0_0_e_15_wd = reg_wdata[15];
	// Trace: design.sv:98454:3
	assign ie0_0_e_16_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98455:3
	assign ie0_0_e_16_wd = reg_wdata[16];
	// Trace: design.sv:98457:3
	assign ie0_0_e_17_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98458:3
	assign ie0_0_e_17_wd = reg_wdata[17];
	// Trace: design.sv:98460:3
	assign ie0_0_e_18_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98461:3
	assign ie0_0_e_18_wd = reg_wdata[18];
	// Trace: design.sv:98463:3
	assign ie0_0_e_19_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98464:3
	assign ie0_0_e_19_wd = reg_wdata[19];
	// Trace: design.sv:98466:3
	assign ie0_0_e_20_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98467:3
	assign ie0_0_e_20_wd = reg_wdata[20];
	// Trace: design.sv:98469:3
	assign ie0_0_e_21_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98470:3
	assign ie0_0_e_21_wd = reg_wdata[21];
	// Trace: design.sv:98472:3
	assign ie0_0_e_22_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98473:3
	assign ie0_0_e_22_wd = reg_wdata[22];
	// Trace: design.sv:98475:3
	assign ie0_0_e_23_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98476:3
	assign ie0_0_e_23_wd = reg_wdata[23];
	// Trace: design.sv:98478:3
	assign ie0_0_e_24_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98479:3
	assign ie0_0_e_24_wd = reg_wdata[24];
	// Trace: design.sv:98481:3
	assign ie0_0_e_25_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98482:3
	assign ie0_0_e_25_wd = reg_wdata[25];
	// Trace: design.sv:98484:3
	assign ie0_0_e_26_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98485:3
	assign ie0_0_e_26_wd = reg_wdata[26];
	// Trace: design.sv:98487:3
	assign ie0_0_e_27_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98488:3
	assign ie0_0_e_27_wd = reg_wdata[27];
	// Trace: design.sv:98490:3
	assign ie0_0_e_28_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98491:3
	assign ie0_0_e_28_wd = reg_wdata[28];
	// Trace: design.sv:98493:3
	assign ie0_0_e_29_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98494:3
	assign ie0_0_e_29_wd = reg_wdata[29];
	// Trace: design.sv:98496:3
	assign ie0_0_e_30_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98497:3
	assign ie0_0_e_30_wd = reg_wdata[30];
	// Trace: design.sv:98499:3
	assign ie0_0_e_31_we = (addr_hit[68] & reg_we) & !reg_error;
	// Trace: design.sv:98500:3
	assign ie0_0_e_31_wd = reg_wdata[31];
	// Trace: design.sv:98502:3
	assign ie0_1_e_32_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98503:3
	assign ie0_1_e_32_wd = reg_wdata[0];
	// Trace: design.sv:98505:3
	assign ie0_1_e_33_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98506:3
	assign ie0_1_e_33_wd = reg_wdata[1];
	// Trace: design.sv:98508:3
	assign ie0_1_e_34_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98509:3
	assign ie0_1_e_34_wd = reg_wdata[2];
	// Trace: design.sv:98511:3
	assign ie0_1_e_35_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98512:3
	assign ie0_1_e_35_wd = reg_wdata[3];
	// Trace: design.sv:98514:3
	assign ie0_1_e_36_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98515:3
	assign ie0_1_e_36_wd = reg_wdata[4];
	// Trace: design.sv:98517:3
	assign ie0_1_e_37_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98518:3
	assign ie0_1_e_37_wd = reg_wdata[5];
	// Trace: design.sv:98520:3
	assign ie0_1_e_38_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98521:3
	assign ie0_1_e_38_wd = reg_wdata[6];
	// Trace: design.sv:98523:3
	assign ie0_1_e_39_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98524:3
	assign ie0_1_e_39_wd = reg_wdata[7];
	// Trace: design.sv:98526:3
	assign ie0_1_e_40_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98527:3
	assign ie0_1_e_40_wd = reg_wdata[8];
	// Trace: design.sv:98529:3
	assign ie0_1_e_41_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98530:3
	assign ie0_1_e_41_wd = reg_wdata[9];
	// Trace: design.sv:98532:3
	assign ie0_1_e_42_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98533:3
	assign ie0_1_e_42_wd = reg_wdata[10];
	// Trace: design.sv:98535:3
	assign ie0_1_e_43_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98536:3
	assign ie0_1_e_43_wd = reg_wdata[11];
	// Trace: design.sv:98538:3
	assign ie0_1_e_44_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98539:3
	assign ie0_1_e_44_wd = reg_wdata[12];
	// Trace: design.sv:98541:3
	assign ie0_1_e_45_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98542:3
	assign ie0_1_e_45_wd = reg_wdata[13];
	// Trace: design.sv:98544:3
	assign ie0_1_e_46_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98545:3
	assign ie0_1_e_46_wd = reg_wdata[14];
	// Trace: design.sv:98547:3
	assign ie0_1_e_47_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98548:3
	assign ie0_1_e_47_wd = reg_wdata[15];
	// Trace: design.sv:98550:3
	assign ie0_1_e_48_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98551:3
	assign ie0_1_e_48_wd = reg_wdata[16];
	// Trace: design.sv:98553:3
	assign ie0_1_e_49_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98554:3
	assign ie0_1_e_49_wd = reg_wdata[17];
	// Trace: design.sv:98556:3
	assign ie0_1_e_50_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98557:3
	assign ie0_1_e_50_wd = reg_wdata[18];
	// Trace: design.sv:98559:3
	assign ie0_1_e_51_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98560:3
	assign ie0_1_e_51_wd = reg_wdata[19];
	// Trace: design.sv:98562:3
	assign ie0_1_e_52_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98563:3
	assign ie0_1_e_52_wd = reg_wdata[20];
	// Trace: design.sv:98565:3
	assign ie0_1_e_53_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98566:3
	assign ie0_1_e_53_wd = reg_wdata[21];
	// Trace: design.sv:98568:3
	assign ie0_1_e_54_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98569:3
	assign ie0_1_e_54_wd = reg_wdata[22];
	// Trace: design.sv:98571:3
	assign ie0_1_e_55_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98572:3
	assign ie0_1_e_55_wd = reg_wdata[23];
	// Trace: design.sv:98574:3
	assign ie0_1_e_56_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98575:3
	assign ie0_1_e_56_wd = reg_wdata[24];
	// Trace: design.sv:98577:3
	assign ie0_1_e_57_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98578:3
	assign ie0_1_e_57_wd = reg_wdata[25];
	// Trace: design.sv:98580:3
	assign ie0_1_e_58_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98581:3
	assign ie0_1_e_58_wd = reg_wdata[26];
	// Trace: design.sv:98583:3
	assign ie0_1_e_59_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98584:3
	assign ie0_1_e_59_wd = reg_wdata[27];
	// Trace: design.sv:98586:3
	assign ie0_1_e_60_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98587:3
	assign ie0_1_e_60_wd = reg_wdata[28];
	// Trace: design.sv:98589:3
	assign ie0_1_e_61_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98590:3
	assign ie0_1_e_61_wd = reg_wdata[29];
	// Trace: design.sv:98592:3
	assign ie0_1_e_62_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98593:3
	assign ie0_1_e_62_wd = reg_wdata[30];
	// Trace: design.sv:98595:3
	assign ie0_1_e_63_we = (addr_hit[69] & reg_we) & !reg_error;
	// Trace: design.sv:98596:3
	assign ie0_1_e_63_wd = reg_wdata[31];
	// Trace: design.sv:98598:3
	assign threshold0_we = (addr_hit[70] & reg_we) & !reg_error;
	// Trace: design.sv:98599:3
	assign threshold0_wd = reg_wdata[2:0];
	// Trace: design.sv:98601:3
	assign cc0_we = (addr_hit[71] & reg_we) & !reg_error;
	// Trace: design.sv:98602:3
	assign cc0_wd = reg_wdata[5:0];
	// Trace: design.sv:98603:3
	assign cc0_re = (addr_hit[71] & reg_re) & !reg_error;
	// Trace: design.sv:98605:3
	assign msip0_we = (addr_hit[72] & reg_we) & !reg_error;
	// Trace: design.sv:98606:3
	assign msip0_wd = reg_wdata[0];
	// Trace: design.sv:98609:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:98610:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:98611:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]: begin
				// Trace: design.sv:98613:9
				reg_rdata_next[0] = ip_0_p_0_qs;
				// Trace: design.sv:98614:9
				reg_rdata_next[1] = ip_0_p_1_qs;
				// Trace: design.sv:98615:9
				reg_rdata_next[2] = ip_0_p_2_qs;
				// Trace: design.sv:98616:9
				reg_rdata_next[3] = ip_0_p_3_qs;
				// Trace: design.sv:98617:9
				reg_rdata_next[4] = ip_0_p_4_qs;
				// Trace: design.sv:98618:9
				reg_rdata_next[5] = ip_0_p_5_qs;
				// Trace: design.sv:98619:9
				reg_rdata_next[6] = ip_0_p_6_qs;
				// Trace: design.sv:98620:9
				reg_rdata_next[7] = ip_0_p_7_qs;
				// Trace: design.sv:98621:9
				reg_rdata_next[8] = ip_0_p_8_qs;
				// Trace: design.sv:98622:9
				reg_rdata_next[9] = ip_0_p_9_qs;
				// Trace: design.sv:98623:9
				reg_rdata_next[10] = ip_0_p_10_qs;
				// Trace: design.sv:98624:9
				reg_rdata_next[11] = ip_0_p_11_qs;
				// Trace: design.sv:98625:9
				reg_rdata_next[12] = ip_0_p_12_qs;
				// Trace: design.sv:98626:9
				reg_rdata_next[13] = ip_0_p_13_qs;
				// Trace: design.sv:98627:9
				reg_rdata_next[14] = ip_0_p_14_qs;
				// Trace: design.sv:98628:9
				reg_rdata_next[15] = ip_0_p_15_qs;
				// Trace: design.sv:98629:9
				reg_rdata_next[16] = ip_0_p_16_qs;
				// Trace: design.sv:98630:9
				reg_rdata_next[17] = ip_0_p_17_qs;
				// Trace: design.sv:98631:9
				reg_rdata_next[18] = ip_0_p_18_qs;
				// Trace: design.sv:98632:9
				reg_rdata_next[19] = ip_0_p_19_qs;
				// Trace: design.sv:98633:9
				reg_rdata_next[20] = ip_0_p_20_qs;
				// Trace: design.sv:98634:9
				reg_rdata_next[21] = ip_0_p_21_qs;
				// Trace: design.sv:98635:9
				reg_rdata_next[22] = ip_0_p_22_qs;
				// Trace: design.sv:98636:9
				reg_rdata_next[23] = ip_0_p_23_qs;
				// Trace: design.sv:98637:9
				reg_rdata_next[24] = ip_0_p_24_qs;
				// Trace: design.sv:98638:9
				reg_rdata_next[25] = ip_0_p_25_qs;
				// Trace: design.sv:98639:9
				reg_rdata_next[26] = ip_0_p_26_qs;
				// Trace: design.sv:98640:9
				reg_rdata_next[27] = ip_0_p_27_qs;
				// Trace: design.sv:98641:9
				reg_rdata_next[28] = ip_0_p_28_qs;
				// Trace: design.sv:98642:9
				reg_rdata_next[29] = ip_0_p_29_qs;
				// Trace: design.sv:98643:9
				reg_rdata_next[30] = ip_0_p_30_qs;
				// Trace: design.sv:98644:9
				reg_rdata_next[31] = ip_0_p_31_qs;
			end
			addr_hit[1]: begin
				// Trace: design.sv:98648:9
				reg_rdata_next[0] = ip_1_p_32_qs;
				// Trace: design.sv:98649:9
				reg_rdata_next[1] = ip_1_p_33_qs;
				// Trace: design.sv:98650:9
				reg_rdata_next[2] = ip_1_p_34_qs;
				// Trace: design.sv:98651:9
				reg_rdata_next[3] = ip_1_p_35_qs;
				// Trace: design.sv:98652:9
				reg_rdata_next[4] = ip_1_p_36_qs;
				// Trace: design.sv:98653:9
				reg_rdata_next[5] = ip_1_p_37_qs;
				// Trace: design.sv:98654:9
				reg_rdata_next[6] = ip_1_p_38_qs;
				// Trace: design.sv:98655:9
				reg_rdata_next[7] = ip_1_p_39_qs;
				// Trace: design.sv:98656:9
				reg_rdata_next[8] = ip_1_p_40_qs;
				// Trace: design.sv:98657:9
				reg_rdata_next[9] = ip_1_p_41_qs;
				// Trace: design.sv:98658:9
				reg_rdata_next[10] = ip_1_p_42_qs;
				// Trace: design.sv:98659:9
				reg_rdata_next[11] = ip_1_p_43_qs;
				// Trace: design.sv:98660:9
				reg_rdata_next[12] = ip_1_p_44_qs;
				// Trace: design.sv:98661:9
				reg_rdata_next[13] = ip_1_p_45_qs;
				// Trace: design.sv:98662:9
				reg_rdata_next[14] = ip_1_p_46_qs;
				// Trace: design.sv:98663:9
				reg_rdata_next[15] = ip_1_p_47_qs;
				// Trace: design.sv:98664:9
				reg_rdata_next[16] = ip_1_p_48_qs;
				// Trace: design.sv:98665:9
				reg_rdata_next[17] = ip_1_p_49_qs;
				// Trace: design.sv:98666:9
				reg_rdata_next[18] = ip_1_p_50_qs;
				// Trace: design.sv:98667:9
				reg_rdata_next[19] = ip_1_p_51_qs;
				// Trace: design.sv:98668:9
				reg_rdata_next[20] = ip_1_p_52_qs;
				// Trace: design.sv:98669:9
				reg_rdata_next[21] = ip_1_p_53_qs;
				// Trace: design.sv:98670:9
				reg_rdata_next[22] = ip_1_p_54_qs;
				// Trace: design.sv:98671:9
				reg_rdata_next[23] = ip_1_p_55_qs;
				// Trace: design.sv:98672:9
				reg_rdata_next[24] = ip_1_p_56_qs;
				// Trace: design.sv:98673:9
				reg_rdata_next[25] = ip_1_p_57_qs;
				// Trace: design.sv:98674:9
				reg_rdata_next[26] = ip_1_p_58_qs;
				// Trace: design.sv:98675:9
				reg_rdata_next[27] = ip_1_p_59_qs;
				// Trace: design.sv:98676:9
				reg_rdata_next[28] = ip_1_p_60_qs;
				// Trace: design.sv:98677:9
				reg_rdata_next[29] = ip_1_p_61_qs;
				// Trace: design.sv:98678:9
				reg_rdata_next[30] = ip_1_p_62_qs;
				// Trace: design.sv:98679:9
				reg_rdata_next[31] = ip_1_p_63_qs;
			end
			addr_hit[2]: begin
				// Trace: design.sv:98683:9
				reg_rdata_next[0] = le_0_le_0_qs;
				// Trace: design.sv:98684:9
				reg_rdata_next[1] = le_0_le_1_qs;
				// Trace: design.sv:98685:9
				reg_rdata_next[2] = le_0_le_2_qs;
				// Trace: design.sv:98686:9
				reg_rdata_next[3] = le_0_le_3_qs;
				// Trace: design.sv:98687:9
				reg_rdata_next[4] = le_0_le_4_qs;
				// Trace: design.sv:98688:9
				reg_rdata_next[5] = le_0_le_5_qs;
				// Trace: design.sv:98689:9
				reg_rdata_next[6] = le_0_le_6_qs;
				// Trace: design.sv:98690:9
				reg_rdata_next[7] = le_0_le_7_qs;
				// Trace: design.sv:98691:9
				reg_rdata_next[8] = le_0_le_8_qs;
				// Trace: design.sv:98692:9
				reg_rdata_next[9] = le_0_le_9_qs;
				// Trace: design.sv:98693:9
				reg_rdata_next[10] = le_0_le_10_qs;
				// Trace: design.sv:98694:9
				reg_rdata_next[11] = le_0_le_11_qs;
				// Trace: design.sv:98695:9
				reg_rdata_next[12] = le_0_le_12_qs;
				// Trace: design.sv:98696:9
				reg_rdata_next[13] = le_0_le_13_qs;
				// Trace: design.sv:98697:9
				reg_rdata_next[14] = le_0_le_14_qs;
				// Trace: design.sv:98698:9
				reg_rdata_next[15] = le_0_le_15_qs;
				// Trace: design.sv:98699:9
				reg_rdata_next[16] = le_0_le_16_qs;
				// Trace: design.sv:98700:9
				reg_rdata_next[17] = le_0_le_17_qs;
				// Trace: design.sv:98701:9
				reg_rdata_next[18] = le_0_le_18_qs;
				// Trace: design.sv:98702:9
				reg_rdata_next[19] = le_0_le_19_qs;
				// Trace: design.sv:98703:9
				reg_rdata_next[20] = le_0_le_20_qs;
				// Trace: design.sv:98704:9
				reg_rdata_next[21] = le_0_le_21_qs;
				// Trace: design.sv:98705:9
				reg_rdata_next[22] = le_0_le_22_qs;
				// Trace: design.sv:98706:9
				reg_rdata_next[23] = le_0_le_23_qs;
				// Trace: design.sv:98707:9
				reg_rdata_next[24] = le_0_le_24_qs;
				// Trace: design.sv:98708:9
				reg_rdata_next[25] = le_0_le_25_qs;
				// Trace: design.sv:98709:9
				reg_rdata_next[26] = le_0_le_26_qs;
				// Trace: design.sv:98710:9
				reg_rdata_next[27] = le_0_le_27_qs;
				// Trace: design.sv:98711:9
				reg_rdata_next[28] = le_0_le_28_qs;
				// Trace: design.sv:98712:9
				reg_rdata_next[29] = le_0_le_29_qs;
				// Trace: design.sv:98713:9
				reg_rdata_next[30] = le_0_le_30_qs;
				// Trace: design.sv:98714:9
				reg_rdata_next[31] = le_0_le_31_qs;
			end
			addr_hit[3]: begin
				// Trace: design.sv:98718:9
				reg_rdata_next[0] = le_1_le_32_qs;
				// Trace: design.sv:98719:9
				reg_rdata_next[1] = le_1_le_33_qs;
				// Trace: design.sv:98720:9
				reg_rdata_next[2] = le_1_le_34_qs;
				// Trace: design.sv:98721:9
				reg_rdata_next[3] = le_1_le_35_qs;
				// Trace: design.sv:98722:9
				reg_rdata_next[4] = le_1_le_36_qs;
				// Trace: design.sv:98723:9
				reg_rdata_next[5] = le_1_le_37_qs;
				// Trace: design.sv:98724:9
				reg_rdata_next[6] = le_1_le_38_qs;
				// Trace: design.sv:98725:9
				reg_rdata_next[7] = le_1_le_39_qs;
				// Trace: design.sv:98726:9
				reg_rdata_next[8] = le_1_le_40_qs;
				// Trace: design.sv:98727:9
				reg_rdata_next[9] = le_1_le_41_qs;
				// Trace: design.sv:98728:9
				reg_rdata_next[10] = le_1_le_42_qs;
				// Trace: design.sv:98729:9
				reg_rdata_next[11] = le_1_le_43_qs;
				// Trace: design.sv:98730:9
				reg_rdata_next[12] = le_1_le_44_qs;
				// Trace: design.sv:98731:9
				reg_rdata_next[13] = le_1_le_45_qs;
				// Trace: design.sv:98732:9
				reg_rdata_next[14] = le_1_le_46_qs;
				// Trace: design.sv:98733:9
				reg_rdata_next[15] = le_1_le_47_qs;
				// Trace: design.sv:98734:9
				reg_rdata_next[16] = le_1_le_48_qs;
				// Trace: design.sv:98735:9
				reg_rdata_next[17] = le_1_le_49_qs;
				// Trace: design.sv:98736:9
				reg_rdata_next[18] = le_1_le_50_qs;
				// Trace: design.sv:98737:9
				reg_rdata_next[19] = le_1_le_51_qs;
				// Trace: design.sv:98738:9
				reg_rdata_next[20] = le_1_le_52_qs;
				// Trace: design.sv:98739:9
				reg_rdata_next[21] = le_1_le_53_qs;
				// Trace: design.sv:98740:9
				reg_rdata_next[22] = le_1_le_54_qs;
				// Trace: design.sv:98741:9
				reg_rdata_next[23] = le_1_le_55_qs;
				// Trace: design.sv:98742:9
				reg_rdata_next[24] = le_1_le_56_qs;
				// Trace: design.sv:98743:9
				reg_rdata_next[25] = le_1_le_57_qs;
				// Trace: design.sv:98744:9
				reg_rdata_next[26] = le_1_le_58_qs;
				// Trace: design.sv:98745:9
				reg_rdata_next[27] = le_1_le_59_qs;
				// Trace: design.sv:98746:9
				reg_rdata_next[28] = le_1_le_60_qs;
				// Trace: design.sv:98747:9
				reg_rdata_next[29] = le_1_le_61_qs;
				// Trace: design.sv:98748:9
				reg_rdata_next[30] = le_1_le_62_qs;
				// Trace: design.sv:98749:9
				reg_rdata_next[31] = le_1_le_63_qs;
			end
			addr_hit[4]:
				// Trace: design.sv:98753:9
				reg_rdata_next[2:0] = prio0_qs;
			addr_hit[5]:
				// Trace: design.sv:98757:9
				reg_rdata_next[2:0] = prio1_qs;
			addr_hit[6]:
				// Trace: design.sv:98761:9
				reg_rdata_next[2:0] = prio2_qs;
			addr_hit[7]:
				// Trace: design.sv:98765:9
				reg_rdata_next[2:0] = prio3_qs;
			addr_hit[8]:
				// Trace: design.sv:98769:9
				reg_rdata_next[2:0] = prio4_qs;
			addr_hit[9]:
				// Trace: design.sv:98773:9
				reg_rdata_next[2:0] = prio5_qs;
			addr_hit[10]:
				// Trace: design.sv:98777:9
				reg_rdata_next[2:0] = prio6_qs;
			addr_hit[11]:
				// Trace: design.sv:98781:9
				reg_rdata_next[2:0] = prio7_qs;
			addr_hit[12]:
				// Trace: design.sv:98785:9
				reg_rdata_next[2:0] = prio8_qs;
			addr_hit[13]:
				// Trace: design.sv:98789:9
				reg_rdata_next[2:0] = prio9_qs;
			addr_hit[14]:
				// Trace: design.sv:98793:9
				reg_rdata_next[2:0] = prio10_qs;
			addr_hit[15]:
				// Trace: design.sv:98797:9
				reg_rdata_next[2:0] = prio11_qs;
			addr_hit[16]:
				// Trace: design.sv:98801:9
				reg_rdata_next[2:0] = prio12_qs;
			addr_hit[17]:
				// Trace: design.sv:98805:9
				reg_rdata_next[2:0] = prio13_qs;
			addr_hit[18]:
				// Trace: design.sv:98809:9
				reg_rdata_next[2:0] = prio14_qs;
			addr_hit[19]:
				// Trace: design.sv:98813:9
				reg_rdata_next[2:0] = prio15_qs;
			addr_hit[20]:
				// Trace: design.sv:98817:9
				reg_rdata_next[2:0] = prio16_qs;
			addr_hit[21]:
				// Trace: design.sv:98821:9
				reg_rdata_next[2:0] = prio17_qs;
			addr_hit[22]:
				// Trace: design.sv:98825:9
				reg_rdata_next[2:0] = prio18_qs;
			addr_hit[23]:
				// Trace: design.sv:98829:9
				reg_rdata_next[2:0] = prio19_qs;
			addr_hit[24]:
				// Trace: design.sv:98833:9
				reg_rdata_next[2:0] = prio20_qs;
			addr_hit[25]:
				// Trace: design.sv:98837:9
				reg_rdata_next[2:0] = prio21_qs;
			addr_hit[26]:
				// Trace: design.sv:98841:9
				reg_rdata_next[2:0] = prio22_qs;
			addr_hit[27]:
				// Trace: design.sv:98845:9
				reg_rdata_next[2:0] = prio23_qs;
			addr_hit[28]:
				// Trace: design.sv:98849:9
				reg_rdata_next[2:0] = prio24_qs;
			addr_hit[29]:
				// Trace: design.sv:98853:9
				reg_rdata_next[2:0] = prio25_qs;
			addr_hit[30]:
				// Trace: design.sv:98857:9
				reg_rdata_next[2:0] = prio26_qs;
			addr_hit[31]:
				// Trace: design.sv:98861:9
				reg_rdata_next[2:0] = prio27_qs;
			addr_hit[32]:
				// Trace: design.sv:98865:9
				reg_rdata_next[2:0] = prio28_qs;
			addr_hit[33]:
				// Trace: design.sv:98869:9
				reg_rdata_next[2:0] = prio29_qs;
			addr_hit[34]:
				// Trace: design.sv:98873:9
				reg_rdata_next[2:0] = prio30_qs;
			addr_hit[35]:
				// Trace: design.sv:98877:9
				reg_rdata_next[2:0] = prio31_qs;
			addr_hit[36]:
				// Trace: design.sv:98881:9
				reg_rdata_next[2:0] = prio32_qs;
			addr_hit[37]:
				// Trace: design.sv:98885:9
				reg_rdata_next[2:0] = prio33_qs;
			addr_hit[38]:
				// Trace: design.sv:98889:9
				reg_rdata_next[2:0] = prio34_qs;
			addr_hit[39]:
				// Trace: design.sv:98893:9
				reg_rdata_next[2:0] = prio35_qs;
			addr_hit[40]:
				// Trace: design.sv:98897:9
				reg_rdata_next[2:0] = prio36_qs;
			addr_hit[41]:
				// Trace: design.sv:98901:9
				reg_rdata_next[2:0] = prio37_qs;
			addr_hit[42]:
				// Trace: design.sv:98905:9
				reg_rdata_next[2:0] = prio38_qs;
			addr_hit[43]:
				// Trace: design.sv:98909:9
				reg_rdata_next[2:0] = prio39_qs;
			addr_hit[44]:
				// Trace: design.sv:98913:9
				reg_rdata_next[2:0] = prio40_qs;
			addr_hit[45]:
				// Trace: design.sv:98917:9
				reg_rdata_next[2:0] = prio41_qs;
			addr_hit[46]:
				// Trace: design.sv:98921:9
				reg_rdata_next[2:0] = prio42_qs;
			addr_hit[47]:
				// Trace: design.sv:98925:9
				reg_rdata_next[2:0] = prio43_qs;
			addr_hit[48]:
				// Trace: design.sv:98929:9
				reg_rdata_next[2:0] = prio44_qs;
			addr_hit[49]:
				// Trace: design.sv:98933:9
				reg_rdata_next[2:0] = prio45_qs;
			addr_hit[50]:
				// Trace: design.sv:98937:9
				reg_rdata_next[2:0] = prio46_qs;
			addr_hit[51]:
				// Trace: design.sv:98941:9
				reg_rdata_next[2:0] = prio47_qs;
			addr_hit[52]:
				// Trace: design.sv:98945:9
				reg_rdata_next[2:0] = prio48_qs;
			addr_hit[53]:
				// Trace: design.sv:98949:9
				reg_rdata_next[2:0] = prio49_qs;
			addr_hit[54]:
				// Trace: design.sv:98953:9
				reg_rdata_next[2:0] = prio50_qs;
			addr_hit[55]:
				// Trace: design.sv:98957:9
				reg_rdata_next[2:0] = prio51_qs;
			addr_hit[56]:
				// Trace: design.sv:98961:9
				reg_rdata_next[2:0] = prio52_qs;
			addr_hit[57]:
				// Trace: design.sv:98965:9
				reg_rdata_next[2:0] = prio53_qs;
			addr_hit[58]:
				// Trace: design.sv:98969:9
				reg_rdata_next[2:0] = prio54_qs;
			addr_hit[59]:
				// Trace: design.sv:98973:9
				reg_rdata_next[2:0] = prio55_qs;
			addr_hit[60]:
				// Trace: design.sv:98977:9
				reg_rdata_next[2:0] = prio56_qs;
			addr_hit[61]:
				// Trace: design.sv:98981:9
				reg_rdata_next[2:0] = prio57_qs;
			addr_hit[62]:
				// Trace: design.sv:98985:9
				reg_rdata_next[2:0] = prio58_qs;
			addr_hit[63]:
				// Trace: design.sv:98989:9
				reg_rdata_next[2:0] = prio59_qs;
			addr_hit[64]:
				// Trace: design.sv:98993:9
				reg_rdata_next[2:0] = prio60_qs;
			addr_hit[65]:
				// Trace: design.sv:98997:9
				reg_rdata_next[2:0] = prio61_qs;
			addr_hit[66]:
				// Trace: design.sv:99001:9
				reg_rdata_next[2:0] = prio62_qs;
			addr_hit[67]:
				// Trace: design.sv:99005:9
				reg_rdata_next[2:0] = prio63_qs;
			addr_hit[68]: begin
				// Trace: design.sv:99009:9
				reg_rdata_next[0] = ie0_0_e_0_qs;
				// Trace: design.sv:99010:9
				reg_rdata_next[1] = ie0_0_e_1_qs;
				// Trace: design.sv:99011:9
				reg_rdata_next[2] = ie0_0_e_2_qs;
				// Trace: design.sv:99012:9
				reg_rdata_next[3] = ie0_0_e_3_qs;
				// Trace: design.sv:99013:9
				reg_rdata_next[4] = ie0_0_e_4_qs;
				// Trace: design.sv:99014:9
				reg_rdata_next[5] = ie0_0_e_5_qs;
				// Trace: design.sv:99015:9
				reg_rdata_next[6] = ie0_0_e_6_qs;
				// Trace: design.sv:99016:9
				reg_rdata_next[7] = ie0_0_e_7_qs;
				// Trace: design.sv:99017:9
				reg_rdata_next[8] = ie0_0_e_8_qs;
				// Trace: design.sv:99018:9
				reg_rdata_next[9] = ie0_0_e_9_qs;
				// Trace: design.sv:99019:9
				reg_rdata_next[10] = ie0_0_e_10_qs;
				// Trace: design.sv:99020:9
				reg_rdata_next[11] = ie0_0_e_11_qs;
				// Trace: design.sv:99021:9
				reg_rdata_next[12] = ie0_0_e_12_qs;
				// Trace: design.sv:99022:9
				reg_rdata_next[13] = ie0_0_e_13_qs;
				// Trace: design.sv:99023:9
				reg_rdata_next[14] = ie0_0_e_14_qs;
				// Trace: design.sv:99024:9
				reg_rdata_next[15] = ie0_0_e_15_qs;
				// Trace: design.sv:99025:9
				reg_rdata_next[16] = ie0_0_e_16_qs;
				// Trace: design.sv:99026:9
				reg_rdata_next[17] = ie0_0_e_17_qs;
				// Trace: design.sv:99027:9
				reg_rdata_next[18] = ie0_0_e_18_qs;
				// Trace: design.sv:99028:9
				reg_rdata_next[19] = ie0_0_e_19_qs;
				// Trace: design.sv:99029:9
				reg_rdata_next[20] = ie0_0_e_20_qs;
				// Trace: design.sv:99030:9
				reg_rdata_next[21] = ie0_0_e_21_qs;
				// Trace: design.sv:99031:9
				reg_rdata_next[22] = ie0_0_e_22_qs;
				// Trace: design.sv:99032:9
				reg_rdata_next[23] = ie0_0_e_23_qs;
				// Trace: design.sv:99033:9
				reg_rdata_next[24] = ie0_0_e_24_qs;
				// Trace: design.sv:99034:9
				reg_rdata_next[25] = ie0_0_e_25_qs;
				// Trace: design.sv:99035:9
				reg_rdata_next[26] = ie0_0_e_26_qs;
				// Trace: design.sv:99036:9
				reg_rdata_next[27] = ie0_0_e_27_qs;
				// Trace: design.sv:99037:9
				reg_rdata_next[28] = ie0_0_e_28_qs;
				// Trace: design.sv:99038:9
				reg_rdata_next[29] = ie0_0_e_29_qs;
				// Trace: design.sv:99039:9
				reg_rdata_next[30] = ie0_0_e_30_qs;
				// Trace: design.sv:99040:9
				reg_rdata_next[31] = ie0_0_e_31_qs;
			end
			addr_hit[69]: begin
				// Trace: design.sv:99044:9
				reg_rdata_next[0] = ie0_1_e_32_qs;
				// Trace: design.sv:99045:9
				reg_rdata_next[1] = ie0_1_e_33_qs;
				// Trace: design.sv:99046:9
				reg_rdata_next[2] = ie0_1_e_34_qs;
				// Trace: design.sv:99047:9
				reg_rdata_next[3] = ie0_1_e_35_qs;
				// Trace: design.sv:99048:9
				reg_rdata_next[4] = ie0_1_e_36_qs;
				// Trace: design.sv:99049:9
				reg_rdata_next[5] = ie0_1_e_37_qs;
				// Trace: design.sv:99050:9
				reg_rdata_next[6] = ie0_1_e_38_qs;
				// Trace: design.sv:99051:9
				reg_rdata_next[7] = ie0_1_e_39_qs;
				// Trace: design.sv:99052:9
				reg_rdata_next[8] = ie0_1_e_40_qs;
				// Trace: design.sv:99053:9
				reg_rdata_next[9] = ie0_1_e_41_qs;
				// Trace: design.sv:99054:9
				reg_rdata_next[10] = ie0_1_e_42_qs;
				// Trace: design.sv:99055:9
				reg_rdata_next[11] = ie0_1_e_43_qs;
				// Trace: design.sv:99056:9
				reg_rdata_next[12] = ie0_1_e_44_qs;
				// Trace: design.sv:99057:9
				reg_rdata_next[13] = ie0_1_e_45_qs;
				// Trace: design.sv:99058:9
				reg_rdata_next[14] = ie0_1_e_46_qs;
				// Trace: design.sv:99059:9
				reg_rdata_next[15] = ie0_1_e_47_qs;
				// Trace: design.sv:99060:9
				reg_rdata_next[16] = ie0_1_e_48_qs;
				// Trace: design.sv:99061:9
				reg_rdata_next[17] = ie0_1_e_49_qs;
				// Trace: design.sv:99062:9
				reg_rdata_next[18] = ie0_1_e_50_qs;
				// Trace: design.sv:99063:9
				reg_rdata_next[19] = ie0_1_e_51_qs;
				// Trace: design.sv:99064:9
				reg_rdata_next[20] = ie0_1_e_52_qs;
				// Trace: design.sv:99065:9
				reg_rdata_next[21] = ie0_1_e_53_qs;
				// Trace: design.sv:99066:9
				reg_rdata_next[22] = ie0_1_e_54_qs;
				// Trace: design.sv:99067:9
				reg_rdata_next[23] = ie0_1_e_55_qs;
				// Trace: design.sv:99068:9
				reg_rdata_next[24] = ie0_1_e_56_qs;
				// Trace: design.sv:99069:9
				reg_rdata_next[25] = ie0_1_e_57_qs;
				// Trace: design.sv:99070:9
				reg_rdata_next[26] = ie0_1_e_58_qs;
				// Trace: design.sv:99071:9
				reg_rdata_next[27] = ie0_1_e_59_qs;
				// Trace: design.sv:99072:9
				reg_rdata_next[28] = ie0_1_e_60_qs;
				// Trace: design.sv:99073:9
				reg_rdata_next[29] = ie0_1_e_61_qs;
				// Trace: design.sv:99074:9
				reg_rdata_next[30] = ie0_1_e_62_qs;
				// Trace: design.sv:99075:9
				reg_rdata_next[31] = ie0_1_e_63_qs;
			end
			addr_hit[70]:
				// Trace: design.sv:99079:9
				reg_rdata_next[2:0] = threshold0_qs;
			addr_hit[71]:
				// Trace: design.sv:99083:9
				reg_rdata_next[5:0] = cc0_qs;
			addr_hit[72]:
				// Trace: design.sv:99087:9
				reg_rdata_next[0] = msip0_qs;
			default:
				// Trace: design.sv:99091:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:99100:3
	wire unused_wdata;
	// Trace: design.sv:99101:3
	wire unused_be;
	// Trace: design.sv:99102:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:99103:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module rv_plic (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	intr_src_i,
	irq_o,
	irq_id_o,
	msip_o
);
	reg _sv2v_0;
	// removed import rv_plic_reg_pkg::*;
	// Trace: design.sv:99137:14
	localparam signed [31:0] rv_plic_reg_pkg_NumSrc = 64;
	localparam signed [31:0] SRCW = 6;
	// Trace: design.sv:99139:3
	input clk_i;
	// Trace: design.sv:99140:3
	input rst_ni;
	// Trace: design.sv:99143:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:99144:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:99147:3
	input [63:0] intr_src_i;
	// Trace: design.sv:99150:3
	localparam signed [31:0] rv_plic_reg_pkg_NumTarget = 1;
	output wire [0:0] irq_o;
	// Trace: design.sv:99151:3
	output wire [(rv_plic_reg_pkg_NumTarget * SRCW) - 1:0] irq_id_o;
	// Trace: design.sv:99153:3
	output wire [0:0] msip_o;
	// Trace: design.sv:99156:3
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_cc0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_ie0_mreg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_le_mreg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_msip0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio10_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio11_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio12_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio13_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio14_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio15_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio16_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio17_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio18_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio19_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio1_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio20_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio21_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio22_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio23_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio24_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio25_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio26_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio27_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio28_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio29_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio2_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio30_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio31_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio32_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio33_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio34_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio35_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio36_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio37_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio38_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio39_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio3_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio40_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio41_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio42_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio43_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio44_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio45_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio46_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio47_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio48_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio49_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio4_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio50_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio51_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio52_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio53_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio54_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio55_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio56_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio57_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio58_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio59_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio5_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio60_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio61_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio62_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio63_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio6_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio7_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio8_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_prio9_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_threshold0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_reg2hw_t
	wire [331:0] reg2hw;
	// Trace: design.sv:99157:3
	// removed localparam type rv_plic_reg_pkg_rv_plic_hw2reg_cc0_reg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_hw2reg_ip_mreg_t
	// removed localparam type rv_plic_reg_pkg_rv_plic_hw2reg_t
	wire [133:0] hw2reg;
	// Trace: design.sv:99159:3
	localparam signed [31:0] MAX_PRIO = 7;
	// Trace: design.sv:99160:3
	localparam signed [31:0] PRIOW = 3;
	// Trace: design.sv:99162:3
	wire [63:0] le;
	// Trace: design.sv:99163:3
	wire [63:0] ip;
	// Trace: design.sv:99165:3
	wire [63:0] ie [0:0];
	// Trace: design.sv:99167:3
	wire [0:0] claim_re;
	// Trace: design.sv:99168:3
	wire [5:0] claim_id [0:0];
	// Trace: design.sv:99169:3
	reg [63:0] claim;
	// Trace: design.sv:99171:3
	wire [0:0] complete_we;
	// Trace: design.sv:99172:3
	wire [5:0] complete_id [0:0];
	// Trace: design.sv:99173:3
	reg [63:0] complete;
	// Trace: design.sv:99175:3
	wire [(rv_plic_reg_pkg_NumTarget * SRCW) - 1:0] cc_id;
	// Trace: design.sv:99177:3
	wire [(rv_plic_reg_pkg_NumSrc * PRIOW) - 1:0] prio;
	// Trace: design.sv:99179:3
	wire [2:0] threshold [0:0];
	// Trace: design.sv:99182:3
	assign cc_id = irq_id_o;
	// Trace: design.sv:99184:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:99185:5
		claim = 1'sb0;
		// Trace: design.sv:99186:5
		begin : sv2v_autoblock_1
			// Trace: design.sv:99186:10
			reg signed [31:0] i;
			// Trace: design.sv:99186:10
			for (i = 0; i < rv_plic_reg_pkg_NumTarget; i = i + 1)
				begin
					// Trace: design.sv:99187:7
					if (claim_re[i])
						// Trace: design.sv:99187:24
						claim[claim_id[i]] = 1'b1;
				end
		end
	end
	// Trace: design.sv:99190:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:99191:5
		complete = 1'sb0;
		// Trace: design.sv:99192:5
		begin : sv2v_autoblock_2
			// Trace: design.sv:99192:10
			reg signed [31:0] i;
			// Trace: design.sv:99192:10
			for (i = 0; i < rv_plic_reg_pkg_NumTarget; i = i + 1)
				begin
					// Trace: design.sv:99193:7
					if (complete_we[i])
						// Trace: design.sv:99193:27
						complete[complete_id[i]] = 1'b1;
				end
		end
	end
	// Trace: design.sv:99207:3
	assign prio[189+:PRIOW] = reg2hw[267-:3];
	// Trace: design.sv:99208:3
	assign prio[186+:PRIOW] = reg2hw[264-:3];
	// Trace: design.sv:99209:3
	assign prio[183+:PRIOW] = reg2hw[261-:3];
	// Trace: design.sv:99210:3
	assign prio[180+:PRIOW] = reg2hw[258-:3];
	// Trace: design.sv:99211:3
	assign prio[177+:PRIOW] = reg2hw[255-:3];
	// Trace: design.sv:99212:3
	assign prio[174+:PRIOW] = reg2hw[252-:3];
	// Trace: design.sv:99213:3
	assign prio[171+:PRIOW] = reg2hw[249-:3];
	// Trace: design.sv:99214:3
	assign prio[168+:PRIOW] = reg2hw[246-:3];
	// Trace: design.sv:99215:3
	assign prio[165+:PRIOW] = reg2hw[243-:3];
	// Trace: design.sv:99216:3
	assign prio[162+:PRIOW] = reg2hw[240-:3];
	// Trace: design.sv:99217:3
	assign prio[159+:PRIOW] = reg2hw[237-:3];
	// Trace: design.sv:99218:3
	assign prio[156+:PRIOW] = reg2hw[234-:3];
	// Trace: design.sv:99219:3
	assign prio[153+:PRIOW] = reg2hw[231-:3];
	// Trace: design.sv:99220:3
	assign prio[150+:PRIOW] = reg2hw[228-:3];
	// Trace: design.sv:99221:3
	assign prio[147+:PRIOW] = reg2hw[225-:3];
	// Trace: design.sv:99222:3
	assign prio[144+:PRIOW] = reg2hw[222-:3];
	// Trace: design.sv:99223:3
	assign prio[141+:PRIOW] = reg2hw[219-:3];
	// Trace: design.sv:99224:3
	assign prio[138+:PRIOW] = reg2hw[216-:3];
	// Trace: design.sv:99225:3
	assign prio[135+:PRIOW] = reg2hw[213-:3];
	// Trace: design.sv:99226:3
	assign prio[132+:PRIOW] = reg2hw[210-:3];
	// Trace: design.sv:99227:3
	assign prio[129+:PRIOW] = reg2hw[207-:3];
	// Trace: design.sv:99228:3
	assign prio[126+:PRIOW] = reg2hw[204-:3];
	// Trace: design.sv:99229:3
	assign prio[123+:PRIOW] = reg2hw[201-:3];
	// Trace: design.sv:99230:3
	assign prio[120+:PRIOW] = reg2hw[198-:3];
	// Trace: design.sv:99231:3
	assign prio[117+:PRIOW] = reg2hw[195-:3];
	// Trace: design.sv:99232:3
	assign prio[114+:PRIOW] = reg2hw[192-:3];
	// Trace: design.sv:99233:3
	assign prio[111+:PRIOW] = reg2hw[189-:3];
	// Trace: design.sv:99234:3
	assign prio[108+:PRIOW] = reg2hw[186-:3];
	// Trace: design.sv:99235:3
	assign prio[105+:PRIOW] = reg2hw[183-:3];
	// Trace: design.sv:99236:3
	assign prio[102+:PRIOW] = reg2hw[180-:3];
	// Trace: design.sv:99237:3
	assign prio[99+:PRIOW] = reg2hw[177-:3];
	// Trace: design.sv:99238:3
	assign prio[96+:PRIOW] = reg2hw[174-:3];
	// Trace: design.sv:99239:3
	assign prio[93+:PRIOW] = reg2hw[171-:3];
	// Trace: design.sv:99240:3
	assign prio[90+:PRIOW] = reg2hw[168-:3];
	// Trace: design.sv:99241:3
	assign prio[87+:PRIOW] = reg2hw[165-:3];
	// Trace: design.sv:99242:3
	assign prio[84+:PRIOW] = reg2hw[162-:3];
	// Trace: design.sv:99243:3
	assign prio[81+:PRIOW] = reg2hw[159-:3];
	// Trace: design.sv:99244:3
	assign prio[78+:PRIOW] = reg2hw[156-:3];
	// Trace: design.sv:99245:3
	assign prio[75+:PRIOW] = reg2hw[153-:3];
	// Trace: design.sv:99246:3
	assign prio[72+:PRIOW] = reg2hw[150-:3];
	// Trace: design.sv:99247:3
	assign prio[69+:PRIOW] = reg2hw[147-:3];
	// Trace: design.sv:99248:3
	assign prio[66+:PRIOW] = reg2hw[144-:3];
	// Trace: design.sv:99249:3
	assign prio[63+:PRIOW] = reg2hw[141-:3];
	// Trace: design.sv:99250:3
	assign prio[60+:PRIOW] = reg2hw[138-:3];
	// Trace: design.sv:99251:3
	assign prio[57+:PRIOW] = reg2hw[135-:3];
	// Trace: design.sv:99252:3
	assign prio[54+:PRIOW] = reg2hw[132-:3];
	// Trace: design.sv:99253:3
	assign prio[51+:PRIOW] = reg2hw[129-:3];
	// Trace: design.sv:99254:3
	assign prio[48+:PRIOW] = reg2hw[126-:3];
	// Trace: design.sv:99255:3
	assign prio[45+:PRIOW] = reg2hw[123-:3];
	// Trace: design.sv:99256:3
	assign prio[42+:PRIOW] = reg2hw[120-:3];
	// Trace: design.sv:99257:3
	assign prio[39+:PRIOW] = reg2hw[117-:3];
	// Trace: design.sv:99258:3
	assign prio[36+:PRIOW] = reg2hw[114-:3];
	// Trace: design.sv:99259:3
	assign prio[33+:PRIOW] = reg2hw[111-:3];
	// Trace: design.sv:99260:3
	assign prio[30+:PRIOW] = reg2hw[108-:3];
	// Trace: design.sv:99261:3
	assign prio[27+:PRIOW] = reg2hw[105-:3];
	// Trace: design.sv:99262:3
	assign prio[24+:PRIOW] = reg2hw[102-:3];
	// Trace: design.sv:99263:3
	assign prio[21+:PRIOW] = reg2hw[99-:3];
	// Trace: design.sv:99264:3
	assign prio[18+:PRIOW] = reg2hw[96-:3];
	// Trace: design.sv:99265:3
	assign prio[15+:PRIOW] = reg2hw[93-:3];
	// Trace: design.sv:99266:3
	assign prio[12+:PRIOW] = reg2hw[90-:3];
	// Trace: design.sv:99267:3
	assign prio[9+:PRIOW] = reg2hw[87-:3];
	// Trace: design.sv:99268:3
	assign prio[6+:PRIOW] = reg2hw[84-:3];
	// Trace: design.sv:99269:3
	assign prio[3+:PRIOW] = reg2hw[81-:3];
	// Trace: design.sv:99270:3
	assign prio[0+:PRIOW] = reg2hw[78-:3];
	// Trace: design.sv:99275:3
	genvar _gv_s_1;
	generate
		for (_gv_s_1 = 0; _gv_s_1 < 64; _gv_s_1 = _gv_s_1 + 1) begin : gen_ie0
			localparam s = _gv_s_1;
			// Trace: design.sv:99276:5
			assign ie[0][s] = reg2hw[12 + s];
		end
	endgenerate
	// Trace: design.sv:99282:3
	assign threshold[0] = reg2hw[11-:3];
	// Trace: design.sv:99287:3
	assign claim_re[0] = reg2hw[1];
	// Trace: design.sv:99288:3
	assign claim_id[0] = irq_id_o[0+:SRCW];
	// Trace: design.sv:99289:3
	assign complete_we[0] = reg2hw[2];
	// Trace: design.sv:99290:3
	assign complete_id[0] = reg2hw[8-:6];
	// Trace: design.sv:99291:3
	assign hw2reg[5-:6] = cc_id[0+:SRCW];
	// Trace: design.sv:99296:3
	assign msip_o[0] = reg2hw[-0];
	// Trace: design.sv:99301:3
	genvar _gv_s_2;
	generate
		for (_gv_s_2 = 0; _gv_s_2 < 64; _gv_s_2 = _gv_s_2 + 1) begin : gen_ip
			localparam s = _gv_s_2;
			// Trace: design.sv:99302:5
			assign hw2reg[6 + (s * 2)] = 1'b1;
			// Trace: design.sv:99303:5
			assign hw2reg[6 + ((s * 2) + 1)] = ip[s];
		end
	endgenerate
	// Trace: design.sv:99309:3
	genvar _gv_s_3;
	generate
		for (_gv_s_3 = 0; _gv_s_3 < 64; _gv_s_3 = _gv_s_3 + 1) begin : gen_le
			localparam s = _gv_s_3;
			// Trace: design.sv:99310:5
			assign le[s] = reg2hw[268 + s];
		end
	endgenerate
	// Trace: design.sv:99316:3
	rv_plic_gateway #(.N_SOURCE(rv_plic_reg_pkg_NumSrc)) u_gateway(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.src_i(intr_src_i),
		.le_i(le),
		.claim_i(claim),
		.complete_i(complete),
		.ip_o(ip)
	);
	// Trace: design.sv:99334:3
	genvar _gv_i_92;
	generate
		for (_gv_i_92 = 0; _gv_i_92 < rv_plic_reg_pkg_NumTarget; _gv_i_92 = _gv_i_92 + 1) begin : gen_target
			localparam i = _gv_i_92;
			// Trace: design.sv:99335:5
			rv_plic_target #(
				.N_SOURCE(rv_plic_reg_pkg_NumSrc),
				.MAX_PRIO(MAX_PRIO)
			) u_target(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.ip_i(ip),
				.ie_i(ie[i]),
				.prio_i(prio),
				.threshold_i(threshold[i]),
				.irq_o(irq_o[i]),
				.irq_id_o(irq_id_o[-i * SRCW+:SRCW])
			);
		end
	endgenerate
	// Trace: design.sv:99359:3
	rv_plic_reg_top u_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.tl_o(tl_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.intg_err_o(),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:99378:3
	genvar _gv_k_15;
	initial _sv2v_0 = 0;
endmodule
// removed package "rv_timer_reg_pkg"
module rv_timer_reg_top (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	reg2hw,
	hw2reg,
	intg_err_o,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:99627:3
	input clk_i;
	// Trace: design.sv:99628:3
	input rst_ni;
	// Trace: design.sv:99630:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:99631:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:99633:3
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_cfg0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_cfg1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_compare_lower0_0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_compare_lower1_0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_compare_upper0_0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_compare_upper1_0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_ctrl_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_enable0_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_enable1_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_state0_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_state1_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_test0_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_test1_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_timer_v_lower0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_timer_v_lower1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_timer_v_upper0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_timer_v_upper1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_t
	output wire [309:0] reg2hw;
	// Trace: design.sv:99634:3
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_intr_state0_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_intr_state1_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_timer_v_lower0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_timer_v_lower1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_timer_v_upper0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_timer_v_upper1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_t
	input wire [135:0] hw2reg;
	// Trace: design.sv:99637:3
	output wire intg_err_o;
	// Trace: design.sv:99640:3
	input devmode_i;
	// Trace: design.sv:99643:3
	// removed import rv_timer_reg_pkg::*;
	// Trace: design.sv:99645:3
	localparam signed [31:0] AW = 10;
	// Trace: design.sv:99646:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:99647:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:99650:3
	wire reg_we;
	// Trace: design.sv:99651:3
	wire reg_re;
	// Trace: design.sv:99652:3
	wire [9:0] reg_addr;
	// Trace: design.sv:99653:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:99654:3
	wire [3:0] reg_be;
	// Trace: design.sv:99655:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:99656:3
	wire reg_error;
	// Trace: design.sv:99658:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:99660:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:99662:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_reg_h2d;
	// Trace: design.sv:99663:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_reg_d2h;
	// Trace: design.sv:99665:3
	assign intg_err_o = 1'sb0;
	// Trace: design.sv:99667:3
	assign tl_reg_h2d = tl_i;
	// Trace: design.sv:99668:3
	assign tl_o = tl_reg_d2h;
	// Trace: design.sv:99670:3
	tlul_adapter_reg #(
		.RegAw(AW),
		.RegDw(DW),
		.EnableDataIntgGen(0)
	) u_reg_if(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_reg_h2d),
		.tl_o(tl_reg_d2h),
		.we_o(reg_we),
		.re_o(reg_re),
		.addr_o(reg_addr),
		.wdata_o(reg_wdata),
		.be_o(reg_be),
		.rdata_i(reg_rdata),
		.error_i(reg_error)
	);
	// Trace: design.sv:99690:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:99691:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:99696:3
	wire ctrl_active_0_qs;
	// Trace: design.sv:99697:3
	wire ctrl_active_0_wd;
	// Trace: design.sv:99698:3
	wire ctrl_active_0_we;
	// Trace: design.sv:99699:3
	wire ctrl_active_1_qs;
	// Trace: design.sv:99700:3
	wire ctrl_active_1_wd;
	// Trace: design.sv:99701:3
	wire ctrl_active_1_we;
	// Trace: design.sv:99702:3
	wire [11:0] cfg0_prescale_qs;
	// Trace: design.sv:99703:3
	wire [11:0] cfg0_prescale_wd;
	// Trace: design.sv:99704:3
	wire cfg0_prescale_we;
	// Trace: design.sv:99705:3
	wire [7:0] cfg0_step_qs;
	// Trace: design.sv:99706:3
	wire [7:0] cfg0_step_wd;
	// Trace: design.sv:99707:3
	wire cfg0_step_we;
	// Trace: design.sv:99708:3
	wire [31:0] timer_v_lower0_qs;
	// Trace: design.sv:99709:3
	wire [31:0] timer_v_lower0_wd;
	// Trace: design.sv:99710:3
	wire timer_v_lower0_we;
	// Trace: design.sv:99711:3
	wire [31:0] timer_v_upper0_qs;
	// Trace: design.sv:99712:3
	wire [31:0] timer_v_upper0_wd;
	// Trace: design.sv:99713:3
	wire timer_v_upper0_we;
	// Trace: design.sv:99714:3
	wire [31:0] compare_lower0_0_qs;
	// Trace: design.sv:99715:3
	wire [31:0] compare_lower0_0_wd;
	// Trace: design.sv:99716:3
	wire compare_lower0_0_we;
	// Trace: design.sv:99717:3
	wire [31:0] compare_upper0_0_qs;
	// Trace: design.sv:99718:3
	wire [31:0] compare_upper0_0_wd;
	// Trace: design.sv:99719:3
	wire compare_upper0_0_we;
	// Trace: design.sv:99720:3
	wire intr_enable0_qs;
	// Trace: design.sv:99721:3
	wire intr_enable0_wd;
	// Trace: design.sv:99722:3
	wire intr_enable0_we;
	// Trace: design.sv:99723:3
	wire intr_state0_qs;
	// Trace: design.sv:99724:3
	wire intr_state0_wd;
	// Trace: design.sv:99725:3
	wire intr_state0_we;
	// Trace: design.sv:99726:3
	wire intr_test0_wd;
	// Trace: design.sv:99727:3
	wire intr_test0_we;
	// Trace: design.sv:99728:3
	wire [11:0] cfg1_prescale_qs;
	// Trace: design.sv:99729:3
	wire [11:0] cfg1_prescale_wd;
	// Trace: design.sv:99730:3
	wire cfg1_prescale_we;
	// Trace: design.sv:99731:3
	wire [7:0] cfg1_step_qs;
	// Trace: design.sv:99732:3
	wire [7:0] cfg1_step_wd;
	// Trace: design.sv:99733:3
	wire cfg1_step_we;
	// Trace: design.sv:99734:3
	wire [31:0] timer_v_lower1_qs;
	// Trace: design.sv:99735:3
	wire [31:0] timer_v_lower1_wd;
	// Trace: design.sv:99736:3
	wire timer_v_lower1_we;
	// Trace: design.sv:99737:3
	wire [31:0] timer_v_upper1_qs;
	// Trace: design.sv:99738:3
	wire [31:0] timer_v_upper1_wd;
	// Trace: design.sv:99739:3
	wire timer_v_upper1_we;
	// Trace: design.sv:99740:3
	wire [31:0] compare_lower1_0_qs;
	// Trace: design.sv:99741:3
	wire [31:0] compare_lower1_0_wd;
	// Trace: design.sv:99742:3
	wire compare_lower1_0_we;
	// Trace: design.sv:99743:3
	wire [31:0] compare_upper1_0_qs;
	// Trace: design.sv:99744:3
	wire [31:0] compare_upper1_0_wd;
	// Trace: design.sv:99745:3
	wire compare_upper1_0_we;
	// Trace: design.sv:99746:3
	wire intr_enable1_qs;
	// Trace: design.sv:99747:3
	wire intr_enable1_wd;
	// Trace: design.sv:99748:3
	wire intr_enable1_we;
	// Trace: design.sv:99749:3
	wire intr_state1_qs;
	// Trace: design.sv:99750:3
	wire intr_state1_wd;
	// Trace: design.sv:99751:3
	wire intr_state1_we;
	// Trace: design.sv:99752:3
	wire intr_test1_wd;
	// Trace: design.sv:99753:3
	wire intr_test1_we;
	// Trace: design.sv:99761:3
	localparam signed [31:0] sv2v_uu_u_ctrl_active_0_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_active_0_d
	localparam [0:0] sv2v_uu_u_ctrl_active_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_active_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_active_0_we),
		.wd(ctrl_active_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_active_0_ext_d_0),
		.qe(),
		.q(reg2hw[308]),
		.qs(ctrl_active_0_qs)
	);
	// Trace: design.sv:99787:3
	localparam signed [31:0] sv2v_uu_u_ctrl_active_1_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_active_1_d
	localparam [0:0] sv2v_uu_u_ctrl_active_1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_active_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_active_1_we),
		.wd(ctrl_active_1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_active_1_ext_d_0),
		.qe(),
		.q(reg2hw[309]),
		.qs(ctrl_active_1_qs)
	);
	// Trace: design.sv:99816:3
	localparam signed [31:0] sv2v_uu_u_cfg0_prescale_DW = 12;
	// removed localparam type sv2v_uu_u_cfg0_prescale_d
	localparam [11:0] sv2v_uu_u_cfg0_prescale_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(12),
		.SWACCESS("RW"),
		.RESVAL(12'h000)
	) u_cfg0_prescale(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cfg0_prescale_we),
		.wd(cfg0_prescale_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cfg0_prescale_ext_d_0),
		.qe(),
		.q(reg2hw[307-:12]),
		.qs(cfg0_prescale_qs)
	);
	// Trace: design.sv:99842:3
	localparam signed [31:0] sv2v_uu_u_cfg0_step_DW = 8;
	// removed localparam type sv2v_uu_u_cfg0_step_d
	localparam [7:0] sv2v_uu_u_cfg0_step_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("RW"),
		.RESVAL(8'h01)
	) u_cfg0_step(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cfg0_step_we),
		.wd(cfg0_step_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cfg0_step_ext_d_0),
		.qe(),
		.q(reg2hw[295-:8]),
		.qs(cfg0_step_qs)
	);
	// Trace: design.sv:99869:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_timer_v_lower0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timer_v_lower0_we),
		.wd(timer_v_lower0_wd),
		.de(hw2reg[103]),
		.d(hw2reg[135-:32]),
		.qe(),
		.q(reg2hw[287-:32]),
		.qs(timer_v_lower0_qs)
	);
	// Trace: design.sv:99896:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_timer_v_upper0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timer_v_upper0_we),
		.wd(timer_v_upper0_wd),
		.de(hw2reg[70]),
		.d(hw2reg[102-:32]),
		.qe(),
		.q(reg2hw[255-:32]),
		.qs(timer_v_upper0_qs)
	);
	// Trace: design.sv:99923:3
	localparam signed [31:0] sv2v_uu_u_compare_lower0_0_DW = 32;
	// removed localparam type sv2v_uu_u_compare_lower0_0_d
	localparam [31:0] sv2v_uu_u_compare_lower0_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'hffffffff)
	) u_compare_lower0_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(compare_lower0_0_we),
		.wd(compare_lower0_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_compare_lower0_0_ext_d_0),
		.qe(reg2hw[191]),
		.q(reg2hw[223-:32]),
		.qs(compare_lower0_0_qs)
	);
	// Trace: design.sv:99950:3
	localparam signed [31:0] sv2v_uu_u_compare_upper0_0_DW = 32;
	// removed localparam type sv2v_uu_u_compare_upper0_0_d
	localparam [31:0] sv2v_uu_u_compare_upper0_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'hffffffff)
	) u_compare_upper0_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(compare_upper0_0_we),
		.wd(compare_upper0_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_compare_upper0_0_ext_d_0),
		.qe(reg2hw[158]),
		.q(reg2hw[190-:32]),
		.qs(compare_upper0_0_qs)
	);
	// Trace: design.sv:99979:3
	localparam signed [31:0] sv2v_uu_u_intr_enable0_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable0_d
	localparam [0:0] sv2v_uu_u_intr_enable0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable0_we),
		.wd(intr_enable0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable0_ext_d_0),
		.qe(),
		.q(reg2hw[157]),
		.qs(intr_enable0_qs)
	);
	// Trace: design.sv:100008:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state0_we),
		.wd(intr_state0_wd),
		.de(hw2reg[68]),
		.d(hw2reg[69]),
		.qe(),
		.q(reg2hw[156]),
		.qs(intr_state0_qs)
	);
	// Trace: design.sv:100037:3
	localparam [31:0] sv2v_uu_u_intr_test0_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test0_d
	localparam [0:0] sv2v_uu_u_intr_test0_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test0(
		.re(1'b0),
		.we(intr_test0_we),
		.wd(intr_test0_wd),
		.d(sv2v_uu_u_intr_test0_ext_d_0),
		.qre(),
		.qe(reg2hw[154]),
		.q(reg2hw[155]),
		.qs()
	);
	// Trace: design.sv:100054:3
	localparam signed [31:0] sv2v_uu_u_cfg1_prescale_DW = 12;
	// removed localparam type sv2v_uu_u_cfg1_prescale_d
	localparam [11:0] sv2v_uu_u_cfg1_prescale_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(12),
		.SWACCESS("RW"),
		.RESVAL(12'h000)
	) u_cfg1_prescale(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cfg1_prescale_we),
		.wd(cfg1_prescale_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cfg1_prescale_ext_d_0),
		.qe(),
		.q(reg2hw[153-:12]),
		.qs(cfg1_prescale_qs)
	);
	// Trace: design.sv:100080:3
	localparam signed [31:0] sv2v_uu_u_cfg1_step_DW = 8;
	// removed localparam type sv2v_uu_u_cfg1_step_d
	localparam [7:0] sv2v_uu_u_cfg1_step_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("RW"),
		.RESVAL(8'h01)
	) u_cfg1_step(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cfg1_step_we),
		.wd(cfg1_step_wd),
		.de(1'b0),
		.d(sv2v_uu_u_cfg1_step_ext_d_0),
		.qe(),
		.q(reg2hw[141-:8]),
		.qs(cfg1_step_qs)
	);
	// Trace: design.sv:100107:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_timer_v_lower1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timer_v_lower1_we),
		.wd(timer_v_lower1_wd),
		.de(hw2reg[35]),
		.d(hw2reg[67-:32]),
		.qe(),
		.q(reg2hw[133-:32]),
		.qs(timer_v_lower1_qs)
	);
	// Trace: design.sv:100134:3
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'h00000000)
	) u_timer_v_upper1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timer_v_upper1_we),
		.wd(timer_v_upper1_wd),
		.de(hw2reg[2]),
		.d(hw2reg[34-:32]),
		.qe(),
		.q(reg2hw[101-:32]),
		.qs(timer_v_upper1_qs)
	);
	// Trace: design.sv:100161:3
	localparam signed [31:0] sv2v_uu_u_compare_lower1_0_DW = 32;
	// removed localparam type sv2v_uu_u_compare_lower1_0_d
	localparam [31:0] sv2v_uu_u_compare_lower1_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'hffffffff)
	) u_compare_lower1_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(compare_lower1_0_we),
		.wd(compare_lower1_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_compare_lower1_0_ext_d_0),
		.qe(reg2hw[37]),
		.q(reg2hw[69-:32]),
		.qs(compare_lower1_0_qs)
	);
	// Trace: design.sv:100188:3
	localparam signed [31:0] sv2v_uu_u_compare_upper1_0_DW = 32;
	// removed localparam type sv2v_uu_u_compare_upper1_0_d
	localparam [31:0] sv2v_uu_u_compare_upper1_0_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(32),
		.SWACCESS("RW"),
		.RESVAL(32'hffffffff)
	) u_compare_upper1_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(compare_upper1_0_we),
		.wd(compare_upper1_0_wd),
		.de(1'b0),
		.d(sv2v_uu_u_compare_upper1_0_ext_d_0),
		.qe(reg2hw[4]),
		.q(reg2hw[36-:32]),
		.qs(compare_upper1_0_qs)
	);
	// Trace: design.sv:100217:3
	localparam signed [31:0] sv2v_uu_u_intr_enable1_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable1_d
	localparam [0:0] sv2v_uu_u_intr_enable1_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable1_we),
		.wd(intr_enable1_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable1_ext_d_0),
		.qe(),
		.q(reg2hw[3]),
		.qs(intr_enable1_qs)
	);
	// Trace: design.sv:100246:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state1_we),
		.wd(intr_state1_wd),
		.de(hw2reg[0]),
		.d(hw2reg[1]),
		.qe(),
		.q(reg2hw[2]),
		.qs(intr_state1_qs)
	);
	// Trace: design.sv:100275:3
	localparam [31:0] sv2v_uu_u_intr_test1_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test1_d
	localparam [0:0] sv2v_uu_u_intr_test1_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test1(
		.re(1'b0),
		.we(intr_test1_we),
		.wd(intr_test1_wd),
		.d(sv2v_uu_u_intr_test1_ext_d_0),
		.qre(),
		.qe(reg2hw[0]),
		.q(reg2hw[1]),
		.qs()
	);
	// Trace: design.sv:100291:3
	reg [16:0] addr_hit;
	// Trace: design.sv:100292:3
	localparam signed [31:0] rv_timer_reg_pkg_BlockAw = 10;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_CFG0_OFFSET = 10'h100;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_CFG1_OFFSET = 10'h200;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_COMPARE_LOWER0_0_OFFSET = 10'h10c;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_COMPARE_LOWER1_0_OFFSET = 10'h20c;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_COMPARE_UPPER0_0_OFFSET = 10'h110;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_COMPARE_UPPER1_0_OFFSET = 10'h210;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_CTRL_OFFSET = 10'h000;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_INTR_ENABLE0_OFFSET = 10'h114;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_INTR_ENABLE1_OFFSET = 10'h214;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_INTR_STATE0_OFFSET = 10'h118;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_INTR_STATE1_OFFSET = 10'h218;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_INTR_TEST0_OFFSET = 10'h11c;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_INTR_TEST1_OFFSET = 10'h21c;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_TIMER_V_LOWER0_OFFSET = 10'h104;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_TIMER_V_LOWER1_OFFSET = 10'h204;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_TIMER_V_UPPER0_OFFSET = 10'h108;
	localparam [9:0] rv_timer_reg_pkg_RV_TIMER_TIMER_V_UPPER1_OFFSET = 10'h208;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:100293:5
		addr_hit = 1'sb0;
		// Trace: design.sv:100294:5
		addr_hit[0] = reg_addr == rv_timer_reg_pkg_RV_TIMER_CTRL_OFFSET;
		// Trace: design.sv:100295:5
		addr_hit[1] = reg_addr == rv_timer_reg_pkg_RV_TIMER_CFG0_OFFSET;
		// Trace: design.sv:100296:5
		addr_hit[2] = reg_addr == rv_timer_reg_pkg_RV_TIMER_TIMER_V_LOWER0_OFFSET;
		// Trace: design.sv:100297:5
		addr_hit[3] = reg_addr == rv_timer_reg_pkg_RV_TIMER_TIMER_V_UPPER0_OFFSET;
		// Trace: design.sv:100298:5
		addr_hit[4] = reg_addr == rv_timer_reg_pkg_RV_TIMER_COMPARE_LOWER0_0_OFFSET;
		// Trace: design.sv:100299:5
		addr_hit[5] = reg_addr == rv_timer_reg_pkg_RV_TIMER_COMPARE_UPPER0_0_OFFSET;
		// Trace: design.sv:100300:5
		addr_hit[6] = reg_addr == rv_timer_reg_pkg_RV_TIMER_INTR_ENABLE0_OFFSET;
		// Trace: design.sv:100301:5
		addr_hit[7] = reg_addr == rv_timer_reg_pkg_RV_TIMER_INTR_STATE0_OFFSET;
		// Trace: design.sv:100302:5
		addr_hit[8] = reg_addr == rv_timer_reg_pkg_RV_TIMER_INTR_TEST0_OFFSET;
		// Trace: design.sv:100303:5
		addr_hit[9] = reg_addr == rv_timer_reg_pkg_RV_TIMER_CFG1_OFFSET;
		// Trace: design.sv:100304:5
		addr_hit[10] = reg_addr == rv_timer_reg_pkg_RV_TIMER_TIMER_V_LOWER1_OFFSET;
		// Trace: design.sv:100305:5
		addr_hit[11] = reg_addr == rv_timer_reg_pkg_RV_TIMER_TIMER_V_UPPER1_OFFSET;
		// Trace: design.sv:100306:5
		addr_hit[12] = reg_addr == rv_timer_reg_pkg_RV_TIMER_COMPARE_LOWER1_0_OFFSET;
		// Trace: design.sv:100307:5
		addr_hit[13] = reg_addr == rv_timer_reg_pkg_RV_TIMER_COMPARE_UPPER1_0_OFFSET;
		// Trace: design.sv:100308:5
		addr_hit[14] = reg_addr == rv_timer_reg_pkg_RV_TIMER_INTR_ENABLE1_OFFSET;
		// Trace: design.sv:100309:5
		addr_hit[15] = reg_addr == rv_timer_reg_pkg_RV_TIMER_INTR_STATE1_OFFSET;
		// Trace: design.sv:100310:5
		addr_hit[16] = reg_addr == rv_timer_reg_pkg_RV_TIMER_INTR_TEST1_OFFSET;
	end
	// Trace: design.sv:100313:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:100316:3
	localparam [67:0] rv_timer_reg_pkg_RV_TIMER_PERMIT = 68'b00010111111111111111111100010001000101111111111111111111000100010001;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:100317:5
		wr_err = reg_we & (((((((((((((((((addr_hit[0] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[64+:4] & ~reg_be)) | (addr_hit[1] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[60+:4] & ~reg_be))) | (addr_hit[2] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[56+:4] & ~reg_be))) | (addr_hit[3] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[52+:4] & ~reg_be))) | (addr_hit[4] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[48+:4] & ~reg_be))) | (addr_hit[5] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[44+:4] & ~reg_be))) | (addr_hit[6] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[40+:4] & ~reg_be))) | (addr_hit[7] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[36+:4] & ~reg_be))) | (addr_hit[8] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[32+:4] & ~reg_be))) | (addr_hit[9] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[28+:4] & ~reg_be))) | (addr_hit[10] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[24+:4] & ~reg_be))) | (addr_hit[11] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[20+:4] & ~reg_be))) | (addr_hit[12] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[16+:4] & ~reg_be))) | (addr_hit[13] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[12+:4] & ~reg_be))) | (addr_hit[14] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[8+:4] & ~reg_be))) | (addr_hit[15] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[4+:4] & ~reg_be))) | (addr_hit[16] & |(rv_timer_reg_pkg_RV_TIMER_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:100337:3
	assign ctrl_active_0_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:100338:3
	assign ctrl_active_0_wd = reg_wdata[0];
	// Trace: design.sv:100340:3
	assign ctrl_active_1_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:100341:3
	assign ctrl_active_1_wd = reg_wdata[1];
	// Trace: design.sv:100343:3
	assign cfg0_prescale_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:100344:3
	assign cfg0_prescale_wd = reg_wdata[11:0];
	// Trace: design.sv:100346:3
	assign cfg0_step_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:100347:3
	assign cfg0_step_wd = reg_wdata[23:16];
	// Trace: design.sv:100349:3
	assign timer_v_lower0_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:100350:3
	assign timer_v_lower0_wd = reg_wdata[31:0];
	// Trace: design.sv:100352:3
	assign timer_v_upper0_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:100353:3
	assign timer_v_upper0_wd = reg_wdata[31:0];
	// Trace: design.sv:100355:3
	assign compare_lower0_0_we = (addr_hit[4] & reg_we) & !reg_error;
	// Trace: design.sv:100356:3
	assign compare_lower0_0_wd = reg_wdata[31:0];
	// Trace: design.sv:100358:3
	assign compare_upper0_0_we = (addr_hit[5] & reg_we) & !reg_error;
	// Trace: design.sv:100359:3
	assign compare_upper0_0_wd = reg_wdata[31:0];
	// Trace: design.sv:100361:3
	assign intr_enable0_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:100362:3
	assign intr_enable0_wd = reg_wdata[0];
	// Trace: design.sv:100364:3
	assign intr_state0_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:100365:3
	assign intr_state0_wd = reg_wdata[0];
	// Trace: design.sv:100367:3
	assign intr_test0_we = (addr_hit[8] & reg_we) & !reg_error;
	// Trace: design.sv:100368:3
	assign intr_test0_wd = reg_wdata[0];
	// Trace: design.sv:100370:3
	assign cfg1_prescale_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:100371:3
	assign cfg1_prescale_wd = reg_wdata[11:0];
	// Trace: design.sv:100373:3
	assign cfg1_step_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:100374:3
	assign cfg1_step_wd = reg_wdata[23:16];
	// Trace: design.sv:100376:3
	assign timer_v_lower1_we = (addr_hit[10] & reg_we) & !reg_error;
	// Trace: design.sv:100377:3
	assign timer_v_lower1_wd = reg_wdata[31:0];
	// Trace: design.sv:100379:3
	assign timer_v_upper1_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:100380:3
	assign timer_v_upper1_wd = reg_wdata[31:0];
	// Trace: design.sv:100382:3
	assign compare_lower1_0_we = (addr_hit[12] & reg_we) & !reg_error;
	// Trace: design.sv:100383:3
	assign compare_lower1_0_wd = reg_wdata[31:0];
	// Trace: design.sv:100385:3
	assign compare_upper1_0_we = (addr_hit[13] & reg_we) & !reg_error;
	// Trace: design.sv:100386:3
	assign compare_upper1_0_wd = reg_wdata[31:0];
	// Trace: design.sv:100388:3
	assign intr_enable1_we = (addr_hit[14] & reg_we) & !reg_error;
	// Trace: design.sv:100389:3
	assign intr_enable1_wd = reg_wdata[0];
	// Trace: design.sv:100391:3
	assign intr_state1_we = (addr_hit[15] & reg_we) & !reg_error;
	// Trace: design.sv:100392:3
	assign intr_state1_wd = reg_wdata[0];
	// Trace: design.sv:100394:3
	assign intr_test1_we = (addr_hit[16] & reg_we) & !reg_error;
	// Trace: design.sv:100395:3
	assign intr_test1_wd = reg_wdata[0];
	// Trace: design.sv:100398:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:100399:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:100400:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]: begin
				// Trace: design.sv:100402:9
				reg_rdata_next[0] = ctrl_active_0_qs;
				// Trace: design.sv:100403:9
				reg_rdata_next[1] = ctrl_active_1_qs;
			end
			addr_hit[1]: begin
				// Trace: design.sv:100407:9
				reg_rdata_next[11:0] = cfg0_prescale_qs;
				// Trace: design.sv:100408:9
				reg_rdata_next[23:16] = cfg0_step_qs;
			end
			addr_hit[2]:
				// Trace: design.sv:100412:9
				reg_rdata_next[31:0] = timer_v_lower0_qs;
			addr_hit[3]:
				// Trace: design.sv:100416:9
				reg_rdata_next[31:0] = timer_v_upper0_qs;
			addr_hit[4]:
				// Trace: design.sv:100420:9
				reg_rdata_next[31:0] = compare_lower0_0_qs;
			addr_hit[5]:
				// Trace: design.sv:100424:9
				reg_rdata_next[31:0] = compare_upper0_0_qs;
			addr_hit[6]:
				// Trace: design.sv:100428:9
				reg_rdata_next[0] = intr_enable0_qs;
			addr_hit[7]:
				// Trace: design.sv:100432:9
				reg_rdata_next[0] = intr_state0_qs;
			addr_hit[8]:
				// Trace: design.sv:100436:9
				reg_rdata_next[0] = 1'sb0;
			addr_hit[9]: begin
				// Trace: design.sv:100440:9
				reg_rdata_next[11:0] = cfg1_prescale_qs;
				// Trace: design.sv:100441:9
				reg_rdata_next[23:16] = cfg1_step_qs;
			end
			addr_hit[10]:
				// Trace: design.sv:100445:9
				reg_rdata_next[31:0] = timer_v_lower1_qs;
			addr_hit[11]:
				// Trace: design.sv:100449:9
				reg_rdata_next[31:0] = timer_v_upper1_qs;
			addr_hit[12]:
				// Trace: design.sv:100453:9
				reg_rdata_next[31:0] = compare_lower1_0_qs;
			addr_hit[13]:
				// Trace: design.sv:100457:9
				reg_rdata_next[31:0] = compare_upper1_0_qs;
			addr_hit[14]:
				// Trace: design.sv:100461:9
				reg_rdata_next[0] = intr_enable1_qs;
			addr_hit[15]:
				// Trace: design.sv:100465:9
				reg_rdata_next[0] = intr_state1_qs;
			addr_hit[16]:
				// Trace: design.sv:100469:9
				reg_rdata_next[0] = 1'sb0;
			default:
				// Trace: design.sv:100473:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:100482:3
	wire unused_wdata;
	// Trace: design.sv:100483:3
	wire unused_be;
	// Trace: design.sv:100484:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:100485:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module timer_core (
	clk_i,
	rst_ni,
	active,
	prescaler,
	step,
	tick,
	mtime_d,
	mtime,
	mtimecmp,
	intr
);
	// Trace: design.sv:100507:13
	parameter signed [31:0] N = 1;
	// Trace: design.sv:100509:3
	input clk_i;
	// Trace: design.sv:100510:3
	input rst_ni;
	// Trace: design.sv:100512:3
	input active;
	// Trace: design.sv:100513:3
	input [11:0] prescaler;
	// Trace: design.sv:100514:3
	input [7:0] step;
	// Trace: design.sv:100516:3
	output wire tick;
	// Trace: design.sv:100517:3
	output wire [63:0] mtime_d;
	// Trace: design.sv:100518:3
	input [63:0] mtime;
	// Trace: design.sv:100519:3
	input [(N * 64) - 1:0] mtimecmp;
	// Trace: design.sv:100521:3
	output wire [N - 1:0] intr;
	// Trace: design.sv:100524:3
	reg [11:0] tick_count;
	// Trace: design.sv:100526:3
	always @(posedge clk_i or negedge rst_ni) begin : generate_tick
		// Trace: design.sv:100527:5
		if (!rst_ni)
			// Trace: design.sv:100528:7
			tick_count <= 12'h000;
		else if (!active)
			// Trace: design.sv:100530:7
			tick_count <= 12'h000;
		else if (tick_count == prescaler)
			// Trace: design.sv:100532:7
			tick_count <= 12'h000;
		else
			// Trace: design.sv:100534:7
			tick_count <= tick_count + 1'b1;
	end
	// Trace: design.sv:100538:3
	assign tick = active & (tick_count >= prescaler);
	// Trace: design.sv:100540:3
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	assign mtime_d = mtime + sv2v_cast_64(step);
	// Trace: design.sv:100544:3
	genvar _gv_t_1;
	generate
		for (_gv_t_1 = 0; _gv_t_1 < N; _gv_t_1 = _gv_t_1 + 1) begin : gen_intr
			localparam t = _gv_t_1;
			// Trace: design.sv:100545:5
			assign intr[t] = active & (mtime >= mtimecmp[((N - 1) - t) * 64+:64]);
		end
	endgenerate
endmodule
module rv_timer (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	intr_timer_expired_0_0_o,
	intr_timer_expired_1_0_o
);
	// Trace: design.sv:100556:3
	input clk_i;
	// Trace: design.sv:100557:3
	input rst_ni;
	// Trace: design.sv:100559:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:100560:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:100562:3
	output wire intr_timer_expired_0_0_o;
	// Trace: design.sv:100563:3
	output wire intr_timer_expired_1_0_o;
	// Trace: design.sv:100566:3
	localparam signed [31:0] N_HARTS = 2;
	// Trace: design.sv:100567:3
	localparam signed [31:0] N_TIMERS = 1;
	// Trace: design.sv:100569:3
	// removed import rv_timer_reg_pkg::*;
	// Trace: design.sv:100571:3
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_cfg0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_cfg1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_compare_lower0_0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_compare_lower1_0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_compare_upper0_0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_compare_upper1_0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_ctrl_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_enable0_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_enable1_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_state0_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_state1_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_test0_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_intr_test1_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_timer_v_lower0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_timer_v_lower1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_timer_v_upper0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_timer_v_upper1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_reg2hw_t
	wire [309:0] reg2hw;
	// Trace: design.sv:100572:3
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_intr_state0_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_intr_state1_mreg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_timer_v_lower0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_timer_v_lower1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_timer_v_upper0_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_timer_v_upper1_reg_t
	// removed localparam type rv_timer_reg_pkg_rv_timer_hw2reg_t
	wire [135:0] hw2reg;
	// Trace: design.sv:100574:3
	wire [1:0] active;
	// Trace: design.sv:100576:3
	wire [11:0] prescaler [0:1];
	// Trace: design.sv:100577:3
	wire [7:0] step [0:1];
	// Trace: design.sv:100579:3
	wire [1:0] tick;
	// Trace: design.sv:100581:3
	wire [63:0] mtime_d [0:1];
	// Trace: design.sv:100582:3
	wire [63:0] mtime [0:1];
	// Trace: design.sv:100583:3
	wire [63:0] mtimecmp [0:1];
	// Trace: design.sv:100584:3
	wire mtimecmp_update [0:1][0:0];
	// Trace: design.sv:100586:3
	wire [(N_HARTS * N_TIMERS) - 1:0] intr_timer_set;
	// Trace: design.sv:100587:3
	wire [(N_HARTS * N_TIMERS) - 1:0] intr_timer_en;
	// Trace: design.sv:100588:3
	wire [(N_HARTS * N_TIMERS) - 1:0] intr_timer_test_q;
	// Trace: design.sv:100589:3
	wire [1:0] intr_timer_test_qe;
	// Trace: design.sv:100590:3
	wire [(N_HARTS * N_TIMERS) - 1:0] intr_timer_state_q;
	// Trace: design.sv:100591:3
	wire [1:0] intr_timer_state_de;
	// Trace: design.sv:100592:3
	wire [(N_HARTS * N_TIMERS) - 1:0] intr_timer_state_d;
	// Trace: design.sv:100594:3
	wire [(N_HARTS * N_TIMERS) - 1:0] intr_out;
	// Trace: design.sv:100602:3
	assign active[0] = reg2hw[308];
	// Trace: design.sv:100603:3
	assign active[1] = reg2hw[309];
	// Trace: design.sv:100605:3
	assign prescaler[0] = reg2hw[307-:12];
	// Trace: design.sv:100606:3
	assign prescaler[1] = reg2hw[153-:12];
	// Trace: design.sv:100608:3
	assign step[0] = reg2hw[295-:8];
	// Trace: design.sv:100609:3
	assign step[1] = reg2hw[141-:8];
	// Trace: design.sv:100611:3
	assign hw2reg[70] = tick[0];
	// Trace: design.sv:100612:3
	assign hw2reg[103] = tick[0];
	// Trace: design.sv:100613:3
	assign hw2reg[2] = tick[1];
	// Trace: design.sv:100614:3
	assign hw2reg[35] = tick[1];
	// Trace: design.sv:100616:3
	assign hw2reg[102-:32] = mtime_d[0][63:32];
	// Trace: design.sv:100617:3
	assign hw2reg[135-:32] = mtime_d[0][31:0];
	// Trace: design.sv:100619:3
	assign hw2reg[34-:32] = mtime_d[1][63:32];
	// Trace: design.sv:100620:3
	assign hw2reg[67-:32] = mtime_d[1][31:0];
	// Trace: design.sv:100622:3
	assign mtime[0] = {reg2hw[255-:32], reg2hw[287-:32]};
	// Trace: design.sv:100623:3
	assign mtime[1] = {reg2hw[101-:32], reg2hw[133-:32]};
	// Trace: design.sv:100625:3
	assign mtimecmp[0][0+:64] = {reg2hw[190-:32], reg2hw[223-:32]};
	// Trace: design.sv:100626:3
	assign mtimecmp[1][0+:64] = {reg2hw[36-:32], reg2hw[69-:32]};
	// Trace: design.sv:100628:3
	assign mtimecmp_update[0][0] = reg2hw[158] | reg2hw[191];
	// Trace: design.sv:100629:3
	assign mtimecmp_update[1][0] = reg2hw[158] | reg2hw[191];
	// Trace: design.sv:100631:3
	assign intr_timer_expired_0_0_o = intr_out[0];
	// Trace: design.sv:100632:3
	assign intr_timer_en[0] = reg2hw[157];
	// Trace: design.sv:100633:3
	assign intr_timer_state_q[0] = reg2hw[156];
	// Trace: design.sv:100634:3
	assign intr_timer_test_q[0] = reg2hw[155];
	// Trace: design.sv:100635:3
	assign intr_timer_test_qe[0] = reg2hw[154];
	// Trace: design.sv:100636:3
	assign intr_timer_expired_1_0_o = intr_out[1];
	// Trace: design.sv:100637:3
	assign intr_timer_en[1] = reg2hw[3];
	// Trace: design.sv:100638:3
	assign intr_timer_state_q[1] = reg2hw[2];
	// Trace: design.sv:100639:3
	assign intr_timer_test_q[1] = reg2hw[1];
	// Trace: design.sv:100640:3
	assign intr_timer_test_qe[1] = reg2hw[0];
	// Trace: design.sv:100642:3
	assign hw2reg[68] = intr_timer_state_de[0] | mtimecmp_update[0][0];
	// Trace: design.sv:100643:3
	assign hw2reg[69] = intr_timer_state_d[0] & ~mtimecmp_update[0][0];
	// Trace: design.sv:100644:3
	assign hw2reg[0] = intr_timer_state_de[1] | mtimecmp_update[1][0];
	// Trace: design.sv:100645:3
	assign hw2reg[1] = intr_timer_state_d[1] & ~mtimecmp_update[1][0];
	// Trace: design.sv:100647:3
	genvar _gv_h_1;
	generate
		for (_gv_h_1 = 0; _gv_h_1 < N_HARTS; _gv_h_1 = _gv_h_1 + 1) begin : gen_harts
			localparam h = _gv_h_1;
			// Trace: design.sv:100648:5
			prim_intr_hw #(.Width(N_TIMERS)) u_intr_hw(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.event_intr_i(intr_timer_set[h]),
				.reg2hw_intr_enable_q_i(intr_timer_en[h * N_TIMERS+:N_TIMERS]),
				.reg2hw_intr_test_q_i(intr_timer_test_q[h * N_TIMERS+:N_TIMERS]),
				.reg2hw_intr_test_qe_i(intr_timer_test_qe[h]),
				.reg2hw_intr_state_q_i(intr_timer_state_q[h * N_TIMERS+:N_TIMERS]),
				.hw2reg_intr_state_de_o(intr_timer_state_de[h]),
				.hw2reg_intr_state_d_o(intr_timer_state_d[h * N_TIMERS+:N_TIMERS]),
				.intr_o(intr_out[h * N_TIMERS+:N_TIMERS])
			);
			// Trace: design.sv:100665:5
			timer_core #(.N(N_TIMERS)) u_core(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.active(active[h]),
				.prescaler(prescaler[h]),
				.step(step[h]),
				.tick(tick[h]),
				.mtime_d(mtime_d[h]),
				.mtime(mtime[h]),
				.mtimecmp(mtimecmp[h]),
				.intr(intr_timer_set[h * N_TIMERS+:N_TIMERS])
			);
		end
	endgenerate
	// Trace: design.sv:100682:3
	rv_timer_reg_top u_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.tl_o(tl_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.intg_err_o(),
		.devmode_i(1'b1)
	);
endmodule
// removed package "uart_reg_pkg"
module uart_reg_top (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	reg2hw,
	hw2reg,
	intg_err_o,
	devmode_i
);
	reg _sv2v_0;
	// Trace: design.sv:101093:3
	input clk_i;
	// Trace: design.sv:101094:3
	input rst_ni;
	// Trace: design.sv:101096:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:101097:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:101099:3
	// removed localparam type uart_reg_pkg_uart_reg2hw_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_fifo_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_enable_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_state_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_test_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_ovrd_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_rdata_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_status_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_timeout_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_wdata_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_t
	output wire [124:0] reg2hw;
	// Trace: design.sv:101100:3
	// removed localparam type uart_reg_pkg_uart_hw2reg_fifo_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_fifo_status_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_intr_state_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_rdata_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_status_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_val_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_t
	input wire [64:0] hw2reg;
	// Trace: design.sv:101103:3
	output wire intg_err_o;
	// Trace: design.sv:101106:3
	input devmode_i;
	// Trace: design.sv:101109:3
	// removed import uart_reg_pkg::*;
	// Trace: design.sv:101111:3
	localparam signed [31:0] AW = 6;
	// Trace: design.sv:101112:3
	localparam signed [31:0] DW = 32;
	// Trace: design.sv:101113:3
	localparam signed [31:0] DBW = 4;
	// Trace: design.sv:101116:3
	wire reg_we;
	// Trace: design.sv:101117:3
	wire reg_re;
	// Trace: design.sv:101118:3
	wire [5:0] reg_addr;
	// Trace: design.sv:101119:3
	wire [31:0] reg_wdata;
	// Trace: design.sv:101120:3
	wire [3:0] reg_be;
	// Trace: design.sv:101121:3
	wire [31:0] reg_rdata;
	// Trace: design.sv:101122:3
	wire reg_error;
	// Trace: design.sv:101124:3
	wire addrmiss;
	reg wr_err;
	// Trace: design.sv:101126:3
	reg [31:0] reg_rdata_next;
	// Trace: design.sv:101128:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_reg_h2d;
	// Trace: design.sv:101129:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_reg_d2h;
	// Trace: design.sv:101131:3
	assign intg_err_o = 1'sb0;
	// Trace: design.sv:101133:3
	assign tl_reg_h2d = tl_i;
	// Trace: design.sv:101134:3
	assign tl_o = tl_reg_d2h;
	// Trace: design.sv:101136:3
	tlul_adapter_reg #(
		.RegAw(AW),
		.RegDw(DW),
		.EnableDataIntgGen(0)
	) u_reg_if(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_reg_h2d),
		.tl_o(tl_reg_d2h),
		.we_o(reg_we),
		.re_o(reg_re),
		.addr_o(reg_addr),
		.wdata_o(reg_wdata),
		.be_o(reg_be),
		.rdata_i(reg_rdata),
		.error_i(reg_error)
	);
	// Trace: design.sv:101156:3
	assign reg_rdata = reg_rdata_next;
	// Trace: design.sv:101157:3
	assign reg_error = (devmode_i & addrmiss) | wr_err;
	// Trace: design.sv:101162:3
	wire intr_state_tx_watermark_qs;
	// Trace: design.sv:101163:3
	wire intr_state_tx_watermark_wd;
	// Trace: design.sv:101164:3
	wire intr_state_tx_watermark_we;
	// Trace: design.sv:101165:3
	wire intr_state_rx_watermark_qs;
	// Trace: design.sv:101166:3
	wire intr_state_rx_watermark_wd;
	// Trace: design.sv:101167:3
	wire intr_state_rx_watermark_we;
	// Trace: design.sv:101168:3
	wire intr_state_tx_empty_qs;
	// Trace: design.sv:101169:3
	wire intr_state_tx_empty_wd;
	// Trace: design.sv:101170:3
	wire intr_state_tx_empty_we;
	// Trace: design.sv:101171:3
	wire intr_state_rx_overflow_qs;
	// Trace: design.sv:101172:3
	wire intr_state_rx_overflow_wd;
	// Trace: design.sv:101173:3
	wire intr_state_rx_overflow_we;
	// Trace: design.sv:101174:3
	wire intr_state_rx_frame_err_qs;
	// Trace: design.sv:101175:3
	wire intr_state_rx_frame_err_wd;
	// Trace: design.sv:101176:3
	wire intr_state_rx_frame_err_we;
	// Trace: design.sv:101177:3
	wire intr_state_rx_break_err_qs;
	// Trace: design.sv:101178:3
	wire intr_state_rx_break_err_wd;
	// Trace: design.sv:101179:3
	wire intr_state_rx_break_err_we;
	// Trace: design.sv:101180:3
	wire intr_state_rx_timeout_qs;
	// Trace: design.sv:101181:3
	wire intr_state_rx_timeout_wd;
	// Trace: design.sv:101182:3
	wire intr_state_rx_timeout_we;
	// Trace: design.sv:101183:3
	wire intr_state_rx_parity_err_qs;
	// Trace: design.sv:101184:3
	wire intr_state_rx_parity_err_wd;
	// Trace: design.sv:101185:3
	wire intr_state_rx_parity_err_we;
	// Trace: design.sv:101186:3
	wire intr_enable_tx_watermark_qs;
	// Trace: design.sv:101187:3
	wire intr_enable_tx_watermark_wd;
	// Trace: design.sv:101188:3
	wire intr_enable_tx_watermark_we;
	// Trace: design.sv:101189:3
	wire intr_enable_rx_watermark_qs;
	// Trace: design.sv:101190:3
	wire intr_enable_rx_watermark_wd;
	// Trace: design.sv:101191:3
	wire intr_enable_rx_watermark_we;
	// Trace: design.sv:101192:3
	wire intr_enable_tx_empty_qs;
	// Trace: design.sv:101193:3
	wire intr_enable_tx_empty_wd;
	// Trace: design.sv:101194:3
	wire intr_enable_tx_empty_we;
	// Trace: design.sv:101195:3
	wire intr_enable_rx_overflow_qs;
	// Trace: design.sv:101196:3
	wire intr_enable_rx_overflow_wd;
	// Trace: design.sv:101197:3
	wire intr_enable_rx_overflow_we;
	// Trace: design.sv:101198:3
	wire intr_enable_rx_frame_err_qs;
	// Trace: design.sv:101199:3
	wire intr_enable_rx_frame_err_wd;
	// Trace: design.sv:101200:3
	wire intr_enable_rx_frame_err_we;
	// Trace: design.sv:101201:3
	wire intr_enable_rx_break_err_qs;
	// Trace: design.sv:101202:3
	wire intr_enable_rx_break_err_wd;
	// Trace: design.sv:101203:3
	wire intr_enable_rx_break_err_we;
	// Trace: design.sv:101204:3
	wire intr_enable_rx_timeout_qs;
	// Trace: design.sv:101205:3
	wire intr_enable_rx_timeout_wd;
	// Trace: design.sv:101206:3
	wire intr_enable_rx_timeout_we;
	// Trace: design.sv:101207:3
	wire intr_enable_rx_parity_err_qs;
	// Trace: design.sv:101208:3
	wire intr_enable_rx_parity_err_wd;
	// Trace: design.sv:101209:3
	wire intr_enable_rx_parity_err_we;
	// Trace: design.sv:101210:3
	wire intr_test_tx_watermark_wd;
	// Trace: design.sv:101211:3
	wire intr_test_tx_watermark_we;
	// Trace: design.sv:101212:3
	wire intr_test_rx_watermark_wd;
	// Trace: design.sv:101213:3
	wire intr_test_rx_watermark_we;
	// Trace: design.sv:101214:3
	wire intr_test_tx_empty_wd;
	// Trace: design.sv:101215:3
	wire intr_test_tx_empty_we;
	// Trace: design.sv:101216:3
	wire intr_test_rx_overflow_wd;
	// Trace: design.sv:101217:3
	wire intr_test_rx_overflow_we;
	// Trace: design.sv:101218:3
	wire intr_test_rx_frame_err_wd;
	// Trace: design.sv:101219:3
	wire intr_test_rx_frame_err_we;
	// Trace: design.sv:101220:3
	wire intr_test_rx_break_err_wd;
	// Trace: design.sv:101221:3
	wire intr_test_rx_break_err_we;
	// Trace: design.sv:101222:3
	wire intr_test_rx_timeout_wd;
	// Trace: design.sv:101223:3
	wire intr_test_rx_timeout_we;
	// Trace: design.sv:101224:3
	wire intr_test_rx_parity_err_wd;
	// Trace: design.sv:101225:3
	wire intr_test_rx_parity_err_we;
	// Trace: design.sv:101226:3
	wire ctrl_tx_qs;
	// Trace: design.sv:101227:3
	wire ctrl_tx_wd;
	// Trace: design.sv:101228:3
	wire ctrl_tx_we;
	// Trace: design.sv:101229:3
	wire ctrl_rx_qs;
	// Trace: design.sv:101230:3
	wire ctrl_rx_wd;
	// Trace: design.sv:101231:3
	wire ctrl_rx_we;
	// Trace: design.sv:101232:3
	wire ctrl_nf_qs;
	// Trace: design.sv:101233:3
	wire ctrl_nf_wd;
	// Trace: design.sv:101234:3
	wire ctrl_nf_we;
	// Trace: design.sv:101235:3
	wire ctrl_slpbk_qs;
	// Trace: design.sv:101236:3
	wire ctrl_slpbk_wd;
	// Trace: design.sv:101237:3
	wire ctrl_slpbk_we;
	// Trace: design.sv:101238:3
	wire ctrl_llpbk_qs;
	// Trace: design.sv:101239:3
	wire ctrl_llpbk_wd;
	// Trace: design.sv:101240:3
	wire ctrl_llpbk_we;
	// Trace: design.sv:101241:3
	wire ctrl_parity_en_qs;
	// Trace: design.sv:101242:3
	wire ctrl_parity_en_wd;
	// Trace: design.sv:101243:3
	wire ctrl_parity_en_we;
	// Trace: design.sv:101244:3
	wire ctrl_parity_odd_qs;
	// Trace: design.sv:101245:3
	wire ctrl_parity_odd_wd;
	// Trace: design.sv:101246:3
	wire ctrl_parity_odd_we;
	// Trace: design.sv:101247:3
	wire [1:0] ctrl_rxblvl_qs;
	// Trace: design.sv:101248:3
	wire [1:0] ctrl_rxblvl_wd;
	// Trace: design.sv:101249:3
	wire ctrl_rxblvl_we;
	// Trace: design.sv:101250:3
	wire [15:0] ctrl_nco_qs;
	// Trace: design.sv:101251:3
	wire [15:0] ctrl_nco_wd;
	// Trace: design.sv:101252:3
	wire ctrl_nco_we;
	// Trace: design.sv:101253:3
	wire status_txfull_qs;
	// Trace: design.sv:101254:3
	wire status_txfull_re;
	// Trace: design.sv:101255:3
	wire status_rxfull_qs;
	// Trace: design.sv:101256:3
	wire status_rxfull_re;
	// Trace: design.sv:101257:3
	wire status_txempty_qs;
	// Trace: design.sv:101258:3
	wire status_txempty_re;
	// Trace: design.sv:101259:3
	wire status_txidle_qs;
	// Trace: design.sv:101260:3
	wire status_txidle_re;
	// Trace: design.sv:101261:3
	wire status_rxidle_qs;
	// Trace: design.sv:101262:3
	wire status_rxidle_re;
	// Trace: design.sv:101263:3
	wire status_rxempty_qs;
	// Trace: design.sv:101264:3
	wire status_rxempty_re;
	// Trace: design.sv:101265:3
	wire [7:0] rdata_qs;
	// Trace: design.sv:101266:3
	wire rdata_re;
	// Trace: design.sv:101267:3
	wire [7:0] wdata_wd;
	// Trace: design.sv:101268:3
	wire wdata_we;
	// Trace: design.sv:101269:3
	wire fifo_ctrl_rxrst_wd;
	// Trace: design.sv:101270:3
	wire fifo_ctrl_rxrst_we;
	// Trace: design.sv:101271:3
	wire fifo_ctrl_txrst_wd;
	// Trace: design.sv:101272:3
	wire fifo_ctrl_txrst_we;
	// Trace: design.sv:101273:3
	wire [2:0] fifo_ctrl_rxilvl_qs;
	// Trace: design.sv:101274:3
	wire [2:0] fifo_ctrl_rxilvl_wd;
	// Trace: design.sv:101275:3
	wire fifo_ctrl_rxilvl_we;
	// Trace: design.sv:101276:3
	wire [1:0] fifo_ctrl_txilvl_qs;
	// Trace: design.sv:101277:3
	wire [1:0] fifo_ctrl_txilvl_wd;
	// Trace: design.sv:101278:3
	wire fifo_ctrl_txilvl_we;
	// Trace: design.sv:101279:3
	wire [5:0] fifo_status_txlvl_qs;
	// Trace: design.sv:101280:3
	wire fifo_status_txlvl_re;
	// Trace: design.sv:101281:3
	wire [5:0] fifo_status_rxlvl_qs;
	// Trace: design.sv:101282:3
	wire fifo_status_rxlvl_re;
	// Trace: design.sv:101283:3
	wire ovrd_txen_qs;
	// Trace: design.sv:101284:3
	wire ovrd_txen_wd;
	// Trace: design.sv:101285:3
	wire ovrd_txen_we;
	// Trace: design.sv:101286:3
	wire ovrd_txval_qs;
	// Trace: design.sv:101287:3
	wire ovrd_txval_wd;
	// Trace: design.sv:101288:3
	wire ovrd_txval_we;
	// Trace: design.sv:101289:3
	wire [15:0] val_qs;
	// Trace: design.sv:101290:3
	wire val_re;
	// Trace: design.sv:101291:3
	wire [23:0] timeout_ctrl_val_qs;
	// Trace: design.sv:101292:3
	wire [23:0] timeout_ctrl_val_wd;
	// Trace: design.sv:101293:3
	wire timeout_ctrl_val_we;
	// Trace: design.sv:101294:3
	wire timeout_ctrl_en_qs;
	// Trace: design.sv:101295:3
	wire timeout_ctrl_en_wd;
	// Trace: design.sv:101296:3
	wire timeout_ctrl_en_we;
	// Trace: design.sv:101302:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_tx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_tx_watermark_we),
		.wd(intr_state_tx_watermark_wd),
		.de(hw2reg[63]),
		.d(hw2reg[64]),
		.qe(),
		.q(reg2hw[124]),
		.qs(intr_state_tx_watermark_qs)
	);
	// Trace: design.sv:101328:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_rx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_rx_watermark_we),
		.wd(intr_state_rx_watermark_wd),
		.de(hw2reg[61]),
		.d(hw2reg[62]),
		.qe(),
		.q(reg2hw[123]),
		.qs(intr_state_rx_watermark_qs)
	);
	// Trace: design.sv:101354:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_tx_empty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_tx_empty_we),
		.wd(intr_state_tx_empty_wd),
		.de(hw2reg[59]),
		.d(hw2reg[60]),
		.qe(),
		.q(reg2hw[122]),
		.qs(intr_state_tx_empty_qs)
	);
	// Trace: design.sv:101380:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_rx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_rx_overflow_we),
		.wd(intr_state_rx_overflow_wd),
		.de(hw2reg[57]),
		.d(hw2reg[58]),
		.qe(),
		.q(reg2hw[121]),
		.qs(intr_state_rx_overflow_qs)
	);
	// Trace: design.sv:101406:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_rx_frame_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_rx_frame_err_we),
		.wd(intr_state_rx_frame_err_wd),
		.de(hw2reg[55]),
		.d(hw2reg[56]),
		.qe(),
		.q(reg2hw[120]),
		.qs(intr_state_rx_frame_err_qs)
	);
	// Trace: design.sv:101432:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_rx_break_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_rx_break_err_we),
		.wd(intr_state_rx_break_err_wd),
		.de(hw2reg[53]),
		.d(hw2reg[54]),
		.qe(),
		.q(reg2hw[119]),
		.qs(intr_state_rx_break_err_qs)
	);
	// Trace: design.sv:101458:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_rx_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_rx_timeout_we),
		.wd(intr_state_rx_timeout_wd),
		.de(hw2reg[51]),
		.d(hw2reg[52]),
		.qe(),
		.q(reg2hw[118]),
		.qs(intr_state_rx_timeout_qs)
	);
	// Trace: design.sv:101484:3
	prim_subreg #(
		.DW(1),
		.SWACCESS("W1C"),
		.RESVAL(1'h0)
	) u_intr_state_rx_parity_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_rx_parity_err_we),
		.wd(intr_state_rx_parity_err_wd),
		.de(hw2reg[49]),
		.d(hw2reg[50]),
		.qe(),
		.q(reg2hw[117]),
		.qs(intr_state_rx_parity_err_qs)
	);
	// Trace: design.sv:101512:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_tx_watermark_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_tx_watermark_d
	localparam [0:0] sv2v_uu_u_intr_enable_tx_watermark_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_tx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_tx_watermark_we),
		.wd(intr_enable_tx_watermark_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_tx_watermark_ext_d_0),
		.qe(),
		.q(reg2hw[116]),
		.qs(intr_enable_tx_watermark_qs)
	);
	// Trace: design.sv:101538:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_rx_watermark_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_rx_watermark_d
	localparam [0:0] sv2v_uu_u_intr_enable_rx_watermark_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_rx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_rx_watermark_we),
		.wd(intr_enable_rx_watermark_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_rx_watermark_ext_d_0),
		.qe(),
		.q(reg2hw[115]),
		.qs(intr_enable_rx_watermark_qs)
	);
	// Trace: design.sv:101564:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_tx_empty_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_tx_empty_d
	localparam [0:0] sv2v_uu_u_intr_enable_tx_empty_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_tx_empty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_tx_empty_we),
		.wd(intr_enable_tx_empty_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_tx_empty_ext_d_0),
		.qe(),
		.q(reg2hw[114]),
		.qs(intr_enable_tx_empty_qs)
	);
	// Trace: design.sv:101590:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_rx_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_rx_overflow_d
	localparam [0:0] sv2v_uu_u_intr_enable_rx_overflow_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_rx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_rx_overflow_we),
		.wd(intr_enable_rx_overflow_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_rx_overflow_ext_d_0),
		.qe(),
		.q(reg2hw[113]),
		.qs(intr_enable_rx_overflow_qs)
	);
	// Trace: design.sv:101616:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_rx_frame_err_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_rx_frame_err_d
	localparam [0:0] sv2v_uu_u_intr_enable_rx_frame_err_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_rx_frame_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_rx_frame_err_we),
		.wd(intr_enable_rx_frame_err_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_rx_frame_err_ext_d_0),
		.qe(),
		.q(reg2hw[112]),
		.qs(intr_enable_rx_frame_err_qs)
	);
	// Trace: design.sv:101642:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_rx_break_err_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_rx_break_err_d
	localparam [0:0] sv2v_uu_u_intr_enable_rx_break_err_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_rx_break_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_rx_break_err_we),
		.wd(intr_enable_rx_break_err_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_rx_break_err_ext_d_0),
		.qe(),
		.q(reg2hw[111]),
		.qs(intr_enable_rx_break_err_qs)
	);
	// Trace: design.sv:101668:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_rx_timeout_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_rx_timeout_d
	localparam [0:0] sv2v_uu_u_intr_enable_rx_timeout_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_rx_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_rx_timeout_we),
		.wd(intr_enable_rx_timeout_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_rx_timeout_ext_d_0),
		.qe(),
		.q(reg2hw[110]),
		.qs(intr_enable_rx_timeout_qs)
	);
	// Trace: design.sv:101694:3
	localparam signed [31:0] sv2v_uu_u_intr_enable_rx_parity_err_DW = 1;
	// removed localparam type sv2v_uu_u_intr_enable_rx_parity_err_d
	localparam [0:0] sv2v_uu_u_intr_enable_rx_parity_err_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_intr_enable_rx_parity_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_rx_parity_err_we),
		.wd(intr_enable_rx_parity_err_wd),
		.de(1'b0),
		.d(sv2v_uu_u_intr_enable_rx_parity_err_ext_d_0),
		.qe(),
		.q(reg2hw[109]),
		.qs(intr_enable_rx_parity_err_qs)
	);
	// Trace: design.sv:101722:3
	localparam [31:0] sv2v_uu_u_intr_test_tx_watermark_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_tx_watermark_d
	localparam [0:0] sv2v_uu_u_intr_test_tx_watermark_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_tx_watermark(
		.re(1'b0),
		.we(intr_test_tx_watermark_we),
		.wd(intr_test_tx_watermark_wd),
		.d(sv2v_uu_u_intr_test_tx_watermark_ext_d_0),
		.qre(),
		.qe(reg2hw[107]),
		.q(reg2hw[108]),
		.qs()
	);
	// Trace: design.sv:101737:3
	localparam [31:0] sv2v_uu_u_intr_test_rx_watermark_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_rx_watermark_d
	localparam [0:0] sv2v_uu_u_intr_test_rx_watermark_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_rx_watermark(
		.re(1'b0),
		.we(intr_test_rx_watermark_we),
		.wd(intr_test_rx_watermark_wd),
		.d(sv2v_uu_u_intr_test_rx_watermark_ext_d_0),
		.qre(),
		.qe(reg2hw[105]),
		.q(reg2hw[106]),
		.qs()
	);
	// Trace: design.sv:101752:3
	localparam [31:0] sv2v_uu_u_intr_test_tx_empty_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_tx_empty_d
	localparam [0:0] sv2v_uu_u_intr_test_tx_empty_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_tx_empty(
		.re(1'b0),
		.we(intr_test_tx_empty_we),
		.wd(intr_test_tx_empty_wd),
		.d(sv2v_uu_u_intr_test_tx_empty_ext_d_0),
		.qre(),
		.qe(reg2hw[103]),
		.q(reg2hw[104]),
		.qs()
	);
	// Trace: design.sv:101767:3
	localparam [31:0] sv2v_uu_u_intr_test_rx_overflow_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_rx_overflow_d
	localparam [0:0] sv2v_uu_u_intr_test_rx_overflow_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_rx_overflow(
		.re(1'b0),
		.we(intr_test_rx_overflow_we),
		.wd(intr_test_rx_overflow_wd),
		.d(sv2v_uu_u_intr_test_rx_overflow_ext_d_0),
		.qre(),
		.qe(reg2hw[101]),
		.q(reg2hw[102]),
		.qs()
	);
	// Trace: design.sv:101782:3
	localparam [31:0] sv2v_uu_u_intr_test_rx_frame_err_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_rx_frame_err_d
	localparam [0:0] sv2v_uu_u_intr_test_rx_frame_err_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_rx_frame_err(
		.re(1'b0),
		.we(intr_test_rx_frame_err_we),
		.wd(intr_test_rx_frame_err_wd),
		.d(sv2v_uu_u_intr_test_rx_frame_err_ext_d_0),
		.qre(),
		.qe(reg2hw[99]),
		.q(reg2hw[100]),
		.qs()
	);
	// Trace: design.sv:101797:3
	localparam [31:0] sv2v_uu_u_intr_test_rx_break_err_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_rx_break_err_d
	localparam [0:0] sv2v_uu_u_intr_test_rx_break_err_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_rx_break_err(
		.re(1'b0),
		.we(intr_test_rx_break_err_we),
		.wd(intr_test_rx_break_err_wd),
		.d(sv2v_uu_u_intr_test_rx_break_err_ext_d_0),
		.qre(),
		.qe(reg2hw[97]),
		.q(reg2hw[98]),
		.qs()
	);
	// Trace: design.sv:101812:3
	localparam [31:0] sv2v_uu_u_intr_test_rx_timeout_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_rx_timeout_d
	localparam [0:0] sv2v_uu_u_intr_test_rx_timeout_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_rx_timeout(
		.re(1'b0),
		.we(intr_test_rx_timeout_we),
		.wd(intr_test_rx_timeout_wd),
		.d(sv2v_uu_u_intr_test_rx_timeout_ext_d_0),
		.qre(),
		.qe(reg2hw[95]),
		.q(reg2hw[96]),
		.qs()
	);
	// Trace: design.sv:101827:3
	localparam [31:0] sv2v_uu_u_intr_test_rx_parity_err_DW = 1;
	// removed localparam type sv2v_uu_u_intr_test_rx_parity_err_d
	localparam [0:0] sv2v_uu_u_intr_test_rx_parity_err_ext_d_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_intr_test_rx_parity_err(
		.re(1'b0),
		.we(intr_test_rx_parity_err_we),
		.wd(intr_test_rx_parity_err_wd),
		.d(sv2v_uu_u_intr_test_rx_parity_err_ext_d_0),
		.qre(),
		.qe(reg2hw[93]),
		.q(reg2hw[94]),
		.qs()
	);
	// Trace: design.sv:101844:3
	localparam signed [31:0] sv2v_uu_u_ctrl_tx_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_tx_d
	localparam [0:0] sv2v_uu_u_ctrl_tx_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_tx(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_tx_we),
		.wd(ctrl_tx_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_tx_ext_d_0),
		.qe(),
		.q(reg2hw[92]),
		.qs(ctrl_tx_qs)
	);
	// Trace: design.sv:101870:3
	localparam signed [31:0] sv2v_uu_u_ctrl_rx_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_rx_d
	localparam [0:0] sv2v_uu_u_ctrl_rx_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_rx(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_rx_we),
		.wd(ctrl_rx_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_rx_ext_d_0),
		.qe(),
		.q(reg2hw[91]),
		.qs(ctrl_rx_qs)
	);
	// Trace: design.sv:101896:3
	localparam signed [31:0] sv2v_uu_u_ctrl_nf_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_nf_d
	localparam [0:0] sv2v_uu_u_ctrl_nf_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_nf(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_nf_we),
		.wd(ctrl_nf_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_nf_ext_d_0),
		.qe(),
		.q(reg2hw[90]),
		.qs(ctrl_nf_qs)
	);
	// Trace: design.sv:101922:3
	localparam signed [31:0] sv2v_uu_u_ctrl_slpbk_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_slpbk_d
	localparam [0:0] sv2v_uu_u_ctrl_slpbk_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_slpbk(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_slpbk_we),
		.wd(ctrl_slpbk_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_slpbk_ext_d_0),
		.qe(),
		.q(reg2hw[89]),
		.qs(ctrl_slpbk_qs)
	);
	// Trace: design.sv:101948:3
	localparam signed [31:0] sv2v_uu_u_ctrl_llpbk_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_llpbk_d
	localparam [0:0] sv2v_uu_u_ctrl_llpbk_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_llpbk(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_llpbk_we),
		.wd(ctrl_llpbk_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_llpbk_ext_d_0),
		.qe(),
		.q(reg2hw[88]),
		.qs(ctrl_llpbk_qs)
	);
	// Trace: design.sv:101974:3
	localparam signed [31:0] sv2v_uu_u_ctrl_parity_en_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_parity_en_d
	localparam [0:0] sv2v_uu_u_ctrl_parity_en_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_parity_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_parity_en_we),
		.wd(ctrl_parity_en_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_parity_en_ext_d_0),
		.qe(),
		.q(reg2hw[87]),
		.qs(ctrl_parity_en_qs)
	);
	// Trace: design.sv:102000:3
	localparam signed [31:0] sv2v_uu_u_ctrl_parity_odd_DW = 1;
	// removed localparam type sv2v_uu_u_ctrl_parity_odd_d
	localparam [0:0] sv2v_uu_u_ctrl_parity_odd_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ctrl_parity_odd(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_parity_odd_we),
		.wd(ctrl_parity_odd_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_parity_odd_ext_d_0),
		.qe(),
		.q(reg2hw[86]),
		.qs(ctrl_parity_odd_qs)
	);
	// Trace: design.sv:102026:3
	localparam signed [31:0] sv2v_uu_u_ctrl_rxblvl_DW = 2;
	// removed localparam type sv2v_uu_u_ctrl_rxblvl_d
	localparam [1:0] sv2v_uu_u_ctrl_rxblvl_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_ctrl_rxblvl(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_rxblvl_we),
		.wd(ctrl_rxblvl_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_rxblvl_ext_d_0),
		.qe(),
		.q(reg2hw[85-:2]),
		.qs(ctrl_rxblvl_qs)
	);
	// Trace: design.sv:102052:3
	localparam signed [31:0] sv2v_uu_u_ctrl_nco_DW = 16;
	// removed localparam type sv2v_uu_u_ctrl_nco_d
	localparam [15:0] sv2v_uu_u_ctrl_nco_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(16),
		.SWACCESS("RW"),
		.RESVAL(16'h0000)
	) u_ctrl_nco(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ctrl_nco_we),
		.wd(ctrl_nco_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ctrl_nco_ext_d_0),
		.qe(),
		.q(reg2hw[83-:16]),
		.qs(ctrl_nco_qs)
	);
	// Trace: design.sv:102080:3
	localparam [31:0] sv2v_uu_u_status_txfull_DW = 1;
	// removed localparam type sv2v_uu_u_status_txfull_wd
	localparam [0:0] sv2v_uu_u_status_txfull_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_txfull(
		.re(status_txfull_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txfull_ext_wd_0),
		.d(hw2reg[48]),
		.qre(reg2hw[66]),
		.qe(),
		.q(reg2hw[67]),
		.qs(status_txfull_qs)
	);
	// Trace: design.sv:102095:3
	localparam [31:0] sv2v_uu_u_status_rxfull_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxfull_wd
	localparam [0:0] sv2v_uu_u_status_rxfull_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_rxfull(
		.re(status_rxfull_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxfull_ext_wd_0),
		.d(hw2reg[47]),
		.qre(reg2hw[64]),
		.qe(),
		.q(reg2hw[65]),
		.qs(status_rxfull_qs)
	);
	// Trace: design.sv:102110:3
	localparam [31:0] sv2v_uu_u_status_txempty_DW = 1;
	// removed localparam type sv2v_uu_u_status_txempty_wd
	localparam [0:0] sv2v_uu_u_status_txempty_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_txempty(
		.re(status_txempty_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txempty_ext_wd_0),
		.d(hw2reg[46]),
		.qre(reg2hw[62]),
		.qe(),
		.q(reg2hw[63]),
		.qs(status_txempty_qs)
	);
	// Trace: design.sv:102125:3
	localparam [31:0] sv2v_uu_u_status_txidle_DW = 1;
	// removed localparam type sv2v_uu_u_status_txidle_wd
	localparam [0:0] sv2v_uu_u_status_txidle_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_txidle(
		.re(status_txidle_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_txidle_ext_wd_0),
		.d(hw2reg[45]),
		.qre(reg2hw[60]),
		.qe(),
		.q(reg2hw[61]),
		.qs(status_txidle_qs)
	);
	// Trace: design.sv:102140:3
	localparam [31:0] sv2v_uu_u_status_rxidle_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxidle_wd
	localparam [0:0] sv2v_uu_u_status_rxidle_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_rxidle(
		.re(status_rxidle_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxidle_ext_wd_0),
		.d(hw2reg[44]),
		.qre(reg2hw[58]),
		.qe(),
		.q(reg2hw[59]),
		.qs(status_rxidle_qs)
	);
	// Trace: design.sv:102155:3
	localparam [31:0] sv2v_uu_u_status_rxempty_DW = 1;
	// removed localparam type sv2v_uu_u_status_rxempty_wd
	localparam [0:0] sv2v_uu_u_status_rxempty_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(1)) u_status_rxempty(
		.re(status_rxempty_re),
		.we(1'b0),
		.wd(sv2v_uu_u_status_rxempty_ext_wd_0),
		.d(hw2reg[43]),
		.qre(reg2hw[56]),
		.qe(),
		.q(reg2hw[57]),
		.qs(status_rxempty_qs)
	);
	// Trace: design.sv:102171:3
	localparam [31:0] sv2v_uu_u_rdata_DW = 8;
	// removed localparam type sv2v_uu_u_rdata_wd
	localparam [7:0] sv2v_uu_u_rdata_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(8)) u_rdata(
		.re(rdata_re),
		.we(1'b0),
		.wd(sv2v_uu_u_rdata_ext_wd_0),
		.d(hw2reg[42-:8]),
		.qre(reg2hw[47]),
		.qe(),
		.q(reg2hw[55-:8]),
		.qs(rdata_qs)
	);
	// Trace: design.sv:102187:3
	localparam signed [31:0] sv2v_uu_u_wdata_DW = 8;
	// removed localparam type sv2v_uu_u_wdata_d
	localparam [7:0] sv2v_uu_u_wdata_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(8),
		.SWACCESS("WO"),
		.RESVAL(8'h00)
	) u_wdata(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wdata_we),
		.wd(wdata_wd),
		.de(1'b0),
		.d(sv2v_uu_u_wdata_ext_d_0),
		.qe(reg2hw[38]),
		.q(reg2hw[46-:8]),
		.qs()
	);
	// Trace: design.sv:102214:3
	localparam signed [31:0] sv2v_uu_u_fifo_ctrl_rxrst_DW = 1;
	// removed localparam type sv2v_uu_u_fifo_ctrl_rxrst_d
	localparam [0:0] sv2v_uu_u_fifo_ctrl_rxrst_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fifo_ctrl_rxrst(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_rxrst_we),
		.wd(fifo_ctrl_rxrst_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fifo_ctrl_rxrst_ext_d_0),
		.qe(reg2hw[36]),
		.q(reg2hw[37]),
		.qs()
	);
	// Trace: design.sv:102239:3
	localparam signed [31:0] sv2v_uu_u_fifo_ctrl_txrst_DW = 1;
	// removed localparam type sv2v_uu_u_fifo_ctrl_txrst_d
	localparam [0:0] sv2v_uu_u_fifo_ctrl_txrst_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("WO"),
		.RESVAL(1'h0)
	) u_fifo_ctrl_txrst(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_txrst_we),
		.wd(fifo_ctrl_txrst_wd),
		.de(1'b0),
		.d(sv2v_uu_u_fifo_ctrl_txrst_ext_d_0),
		.qe(reg2hw[34]),
		.q(reg2hw[35]),
		.qs()
	);
	// Trace: design.sv:102264:3
	prim_subreg #(
		.DW(3),
		.SWACCESS("RW"),
		.RESVAL(3'h0)
	) u_fifo_ctrl_rxilvl(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_rxilvl_we),
		.wd(fifo_ctrl_rxilvl_wd),
		.de(hw2reg[31]),
		.d(hw2reg[34-:3]),
		.qe(reg2hw[30]),
		.q(reg2hw[33-:3]),
		.qs(fifo_ctrl_rxilvl_qs)
	);
	// Trace: design.sv:102290:3
	prim_subreg #(
		.DW(2),
		.SWACCESS("RW"),
		.RESVAL(2'h0)
	) u_fifo_ctrl_txilvl(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(fifo_ctrl_txilvl_we),
		.wd(fifo_ctrl_txilvl_wd),
		.de(hw2reg[28]),
		.d(hw2reg[30-:2]),
		.qe(reg2hw[27]),
		.q(reg2hw[29-:2]),
		.qs(fifo_ctrl_txilvl_qs)
	);
	// Trace: design.sv:102318:3
	localparam [31:0] sv2v_uu_u_fifo_status_txlvl_DW = 6;
	// removed localparam type sv2v_uu_u_fifo_status_txlvl_wd
	localparam [5:0] sv2v_uu_u_fifo_status_txlvl_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(6)) u_fifo_status_txlvl(
		.re(fifo_status_txlvl_re),
		.we(1'b0),
		.wd(sv2v_uu_u_fifo_status_txlvl_ext_wd_0),
		.d(hw2reg[27-:6]),
		.qre(),
		.qe(),
		.q(),
		.qs(fifo_status_txlvl_qs)
	);
	// Trace: design.sv:102333:3
	localparam [31:0] sv2v_uu_u_fifo_status_rxlvl_DW = 6;
	// removed localparam type sv2v_uu_u_fifo_status_rxlvl_wd
	localparam [5:0] sv2v_uu_u_fifo_status_rxlvl_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(6)) u_fifo_status_rxlvl(
		.re(fifo_status_rxlvl_re),
		.we(1'b0),
		.wd(sv2v_uu_u_fifo_status_rxlvl_ext_wd_0),
		.d(hw2reg[21-:6]),
		.qre(),
		.qe(),
		.q(),
		.qs(fifo_status_rxlvl_qs)
	);
	// Trace: design.sv:102350:3
	localparam signed [31:0] sv2v_uu_u_ovrd_txen_DW = 1;
	// removed localparam type sv2v_uu_u_ovrd_txen_d
	localparam [0:0] sv2v_uu_u_ovrd_txen_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ovrd_txen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ovrd_txen_we),
		.wd(ovrd_txen_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ovrd_txen_ext_d_0),
		.qe(),
		.q(reg2hw[26]),
		.qs(ovrd_txen_qs)
	);
	// Trace: design.sv:102376:3
	localparam signed [31:0] sv2v_uu_u_ovrd_txval_DW = 1;
	// removed localparam type sv2v_uu_u_ovrd_txval_d
	localparam [0:0] sv2v_uu_u_ovrd_txval_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_ovrd_txval(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ovrd_txval_we),
		.wd(ovrd_txval_wd),
		.de(1'b0),
		.d(sv2v_uu_u_ovrd_txval_ext_d_0),
		.qe(),
		.q(reg2hw[25]),
		.qs(ovrd_txval_qs)
	);
	// Trace: design.sv:102403:3
	localparam [31:0] sv2v_uu_u_val_DW = 16;
	// removed localparam type sv2v_uu_u_val_wd
	localparam [15:0] sv2v_uu_u_val_ext_wd_0 = 1'sb0;
	prim_subreg_ext #(.DW(16)) u_val(
		.re(val_re),
		.we(1'b0),
		.wd(sv2v_uu_u_val_ext_wd_0),
		.d(hw2reg[15-:16]),
		.qre(),
		.qe(),
		.q(),
		.qs(val_qs)
	);
	// Trace: design.sv:102420:3
	localparam signed [31:0] sv2v_uu_u_timeout_ctrl_val_DW = 24;
	// removed localparam type sv2v_uu_u_timeout_ctrl_val_d
	localparam [23:0] sv2v_uu_u_timeout_ctrl_val_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(24),
		.SWACCESS("RW"),
		.RESVAL(24'h000000)
	) u_timeout_ctrl_val(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timeout_ctrl_val_we),
		.wd(timeout_ctrl_val_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timeout_ctrl_val_ext_d_0),
		.qe(),
		.q(reg2hw[24-:24]),
		.qs(timeout_ctrl_val_qs)
	);
	// Trace: design.sv:102446:3
	localparam signed [31:0] sv2v_uu_u_timeout_ctrl_en_DW = 1;
	// removed localparam type sv2v_uu_u_timeout_ctrl_en_d
	localparam [0:0] sv2v_uu_u_timeout_ctrl_en_ext_d_0 = 1'sb0;
	prim_subreg #(
		.DW(1),
		.SWACCESS("RW"),
		.RESVAL(1'h0)
	) u_timeout_ctrl_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(timeout_ctrl_en_we),
		.wd(timeout_ctrl_en_wd),
		.de(1'b0),
		.d(sv2v_uu_u_timeout_ctrl_en_ext_d_0),
		.qe(),
		.q(reg2hw[0]),
		.qs(timeout_ctrl_en_qs)
	);
	// Trace: design.sv:102473:3
	reg [11:0] addr_hit;
	// Trace: design.sv:102474:3
	localparam signed [31:0] uart_reg_pkg_BlockAw = 6;
	localparam [5:0] uart_reg_pkg_UART_CTRL_OFFSET = 6'h0c;
	localparam [5:0] uart_reg_pkg_UART_FIFO_CTRL_OFFSET = 6'h1c;
	localparam [5:0] uart_reg_pkg_UART_FIFO_STATUS_OFFSET = 6'h20;
	localparam [5:0] uart_reg_pkg_UART_INTR_ENABLE_OFFSET = 6'h04;
	localparam [5:0] uart_reg_pkg_UART_INTR_STATE_OFFSET = 6'h00;
	localparam [5:0] uart_reg_pkg_UART_INTR_TEST_OFFSET = 6'h08;
	localparam [5:0] uart_reg_pkg_UART_OVRD_OFFSET = 6'h24;
	localparam [5:0] uart_reg_pkg_UART_RDATA_OFFSET = 6'h14;
	localparam [5:0] uart_reg_pkg_UART_STATUS_OFFSET = 6'h10;
	localparam [5:0] uart_reg_pkg_UART_TIMEOUT_CTRL_OFFSET = 6'h2c;
	localparam [5:0] uart_reg_pkg_UART_VAL_OFFSET = 6'h28;
	localparam [5:0] uart_reg_pkg_UART_WDATA_OFFSET = 6'h18;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:102475:5
		addr_hit = 1'sb0;
		// Trace: design.sv:102476:5
		addr_hit[0] = reg_addr == uart_reg_pkg_UART_INTR_STATE_OFFSET;
		// Trace: design.sv:102477:5
		addr_hit[1] = reg_addr == uart_reg_pkg_UART_INTR_ENABLE_OFFSET;
		// Trace: design.sv:102478:5
		addr_hit[2] = reg_addr == uart_reg_pkg_UART_INTR_TEST_OFFSET;
		// Trace: design.sv:102479:5
		addr_hit[3] = reg_addr == uart_reg_pkg_UART_CTRL_OFFSET;
		// Trace: design.sv:102480:5
		addr_hit[4] = reg_addr == uart_reg_pkg_UART_STATUS_OFFSET;
		// Trace: design.sv:102481:5
		addr_hit[5] = reg_addr == uart_reg_pkg_UART_RDATA_OFFSET;
		// Trace: design.sv:102482:5
		addr_hit[6] = reg_addr == uart_reg_pkg_UART_WDATA_OFFSET;
		// Trace: design.sv:102483:5
		addr_hit[7] = reg_addr == uart_reg_pkg_UART_FIFO_CTRL_OFFSET;
		// Trace: design.sv:102484:5
		addr_hit[8] = reg_addr == uart_reg_pkg_UART_FIFO_STATUS_OFFSET;
		// Trace: design.sv:102485:5
		addr_hit[9] = reg_addr == uart_reg_pkg_UART_OVRD_OFFSET;
		// Trace: design.sv:102486:5
		addr_hit[10] = reg_addr == uart_reg_pkg_UART_VAL_OFFSET;
		// Trace: design.sv:102487:5
		addr_hit[11] = reg_addr == uart_reg_pkg_UART_TIMEOUT_CTRL_OFFSET;
	end
	// Trace: design.sv:102490:3
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	// Trace: design.sv:102493:3
	localparam [47:0] uart_reg_pkg_UART_PERMIT = 48'b000100010001111100010001000100010111000100111111;
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:102494:5
		wr_err = reg_we & ((((((((((((addr_hit[0] & |(uart_reg_pkg_UART_PERMIT[44+:4] & ~reg_be)) | (addr_hit[1] & |(uart_reg_pkg_UART_PERMIT[40+:4] & ~reg_be))) | (addr_hit[2] & |(uart_reg_pkg_UART_PERMIT[36+:4] & ~reg_be))) | (addr_hit[3] & |(uart_reg_pkg_UART_PERMIT[32+:4] & ~reg_be))) | (addr_hit[4] & |(uart_reg_pkg_UART_PERMIT[28+:4] & ~reg_be))) | (addr_hit[5] & |(uart_reg_pkg_UART_PERMIT[24+:4] & ~reg_be))) | (addr_hit[6] & |(uart_reg_pkg_UART_PERMIT[20+:4] & ~reg_be))) | (addr_hit[7] & |(uart_reg_pkg_UART_PERMIT[16+:4] & ~reg_be))) | (addr_hit[8] & |(uart_reg_pkg_UART_PERMIT[12+:4] & ~reg_be))) | (addr_hit[9] & |(uart_reg_pkg_UART_PERMIT[8+:4] & ~reg_be))) | (addr_hit[10] & |(uart_reg_pkg_UART_PERMIT[4+:4] & ~reg_be))) | (addr_hit[11] & |(uart_reg_pkg_UART_PERMIT[0+:4] & ~reg_be)));
	end
	// Trace: design.sv:102509:3
	assign intr_state_tx_watermark_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:102510:3
	assign intr_state_tx_watermark_wd = reg_wdata[0];
	// Trace: design.sv:102512:3
	assign intr_state_rx_watermark_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:102513:3
	assign intr_state_rx_watermark_wd = reg_wdata[1];
	// Trace: design.sv:102515:3
	assign intr_state_tx_empty_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:102516:3
	assign intr_state_tx_empty_wd = reg_wdata[2];
	// Trace: design.sv:102518:3
	assign intr_state_rx_overflow_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:102519:3
	assign intr_state_rx_overflow_wd = reg_wdata[3];
	// Trace: design.sv:102521:3
	assign intr_state_rx_frame_err_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:102522:3
	assign intr_state_rx_frame_err_wd = reg_wdata[4];
	// Trace: design.sv:102524:3
	assign intr_state_rx_break_err_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:102525:3
	assign intr_state_rx_break_err_wd = reg_wdata[5];
	// Trace: design.sv:102527:3
	assign intr_state_rx_timeout_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:102528:3
	assign intr_state_rx_timeout_wd = reg_wdata[6];
	// Trace: design.sv:102530:3
	assign intr_state_rx_parity_err_we = (addr_hit[0] & reg_we) & !reg_error;
	// Trace: design.sv:102531:3
	assign intr_state_rx_parity_err_wd = reg_wdata[7];
	// Trace: design.sv:102533:3
	assign intr_enable_tx_watermark_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:102534:3
	assign intr_enable_tx_watermark_wd = reg_wdata[0];
	// Trace: design.sv:102536:3
	assign intr_enable_rx_watermark_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:102537:3
	assign intr_enable_rx_watermark_wd = reg_wdata[1];
	// Trace: design.sv:102539:3
	assign intr_enable_tx_empty_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:102540:3
	assign intr_enable_tx_empty_wd = reg_wdata[2];
	// Trace: design.sv:102542:3
	assign intr_enable_rx_overflow_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:102543:3
	assign intr_enable_rx_overflow_wd = reg_wdata[3];
	// Trace: design.sv:102545:3
	assign intr_enable_rx_frame_err_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:102546:3
	assign intr_enable_rx_frame_err_wd = reg_wdata[4];
	// Trace: design.sv:102548:3
	assign intr_enable_rx_break_err_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:102549:3
	assign intr_enable_rx_break_err_wd = reg_wdata[5];
	// Trace: design.sv:102551:3
	assign intr_enable_rx_timeout_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:102552:3
	assign intr_enable_rx_timeout_wd = reg_wdata[6];
	// Trace: design.sv:102554:3
	assign intr_enable_rx_parity_err_we = (addr_hit[1] & reg_we) & !reg_error;
	// Trace: design.sv:102555:3
	assign intr_enable_rx_parity_err_wd = reg_wdata[7];
	// Trace: design.sv:102557:3
	assign intr_test_tx_watermark_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:102558:3
	assign intr_test_tx_watermark_wd = reg_wdata[0];
	// Trace: design.sv:102560:3
	assign intr_test_rx_watermark_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:102561:3
	assign intr_test_rx_watermark_wd = reg_wdata[1];
	// Trace: design.sv:102563:3
	assign intr_test_tx_empty_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:102564:3
	assign intr_test_tx_empty_wd = reg_wdata[2];
	// Trace: design.sv:102566:3
	assign intr_test_rx_overflow_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:102567:3
	assign intr_test_rx_overflow_wd = reg_wdata[3];
	// Trace: design.sv:102569:3
	assign intr_test_rx_frame_err_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:102570:3
	assign intr_test_rx_frame_err_wd = reg_wdata[4];
	// Trace: design.sv:102572:3
	assign intr_test_rx_break_err_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:102573:3
	assign intr_test_rx_break_err_wd = reg_wdata[5];
	// Trace: design.sv:102575:3
	assign intr_test_rx_timeout_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:102576:3
	assign intr_test_rx_timeout_wd = reg_wdata[6];
	// Trace: design.sv:102578:3
	assign intr_test_rx_parity_err_we = (addr_hit[2] & reg_we) & !reg_error;
	// Trace: design.sv:102579:3
	assign intr_test_rx_parity_err_wd = reg_wdata[7];
	// Trace: design.sv:102581:3
	assign ctrl_tx_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102582:3
	assign ctrl_tx_wd = reg_wdata[0];
	// Trace: design.sv:102584:3
	assign ctrl_rx_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102585:3
	assign ctrl_rx_wd = reg_wdata[1];
	// Trace: design.sv:102587:3
	assign ctrl_nf_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102588:3
	assign ctrl_nf_wd = reg_wdata[2];
	// Trace: design.sv:102590:3
	assign ctrl_slpbk_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102591:3
	assign ctrl_slpbk_wd = reg_wdata[4];
	// Trace: design.sv:102593:3
	assign ctrl_llpbk_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102594:3
	assign ctrl_llpbk_wd = reg_wdata[5];
	// Trace: design.sv:102596:3
	assign ctrl_parity_en_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102597:3
	assign ctrl_parity_en_wd = reg_wdata[6];
	// Trace: design.sv:102599:3
	assign ctrl_parity_odd_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102600:3
	assign ctrl_parity_odd_wd = reg_wdata[7];
	// Trace: design.sv:102602:3
	assign ctrl_rxblvl_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102603:3
	assign ctrl_rxblvl_wd = reg_wdata[9:8];
	// Trace: design.sv:102605:3
	assign ctrl_nco_we = (addr_hit[3] & reg_we) & !reg_error;
	// Trace: design.sv:102606:3
	assign ctrl_nco_wd = reg_wdata[31:16];
	// Trace: design.sv:102608:3
	assign status_txfull_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:102610:3
	assign status_rxfull_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:102612:3
	assign status_txempty_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:102614:3
	assign status_txidle_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:102616:3
	assign status_rxidle_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:102618:3
	assign status_rxempty_re = (addr_hit[4] & reg_re) & !reg_error;
	// Trace: design.sv:102620:3
	assign rdata_re = (addr_hit[5] & reg_re) & !reg_error;
	// Trace: design.sv:102622:3
	assign wdata_we = (addr_hit[6] & reg_we) & !reg_error;
	// Trace: design.sv:102623:3
	assign wdata_wd = reg_wdata[7:0];
	// Trace: design.sv:102625:3
	assign fifo_ctrl_rxrst_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:102626:3
	assign fifo_ctrl_rxrst_wd = reg_wdata[0];
	// Trace: design.sv:102628:3
	assign fifo_ctrl_txrst_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:102629:3
	assign fifo_ctrl_txrst_wd = reg_wdata[1];
	// Trace: design.sv:102631:3
	assign fifo_ctrl_rxilvl_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:102632:3
	assign fifo_ctrl_rxilvl_wd = reg_wdata[4:2];
	// Trace: design.sv:102634:3
	assign fifo_ctrl_txilvl_we = (addr_hit[7] & reg_we) & !reg_error;
	// Trace: design.sv:102635:3
	assign fifo_ctrl_txilvl_wd = reg_wdata[6:5];
	// Trace: design.sv:102637:3
	assign fifo_status_txlvl_re = (addr_hit[8] & reg_re) & !reg_error;
	// Trace: design.sv:102639:3
	assign fifo_status_rxlvl_re = (addr_hit[8] & reg_re) & !reg_error;
	// Trace: design.sv:102641:3
	assign ovrd_txen_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:102642:3
	assign ovrd_txen_wd = reg_wdata[0];
	// Trace: design.sv:102644:3
	assign ovrd_txval_we = (addr_hit[9] & reg_we) & !reg_error;
	// Trace: design.sv:102645:3
	assign ovrd_txval_wd = reg_wdata[1];
	// Trace: design.sv:102647:3
	assign val_re = (addr_hit[10] & reg_re) & !reg_error;
	// Trace: design.sv:102649:3
	assign timeout_ctrl_val_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:102650:3
	assign timeout_ctrl_val_wd = reg_wdata[23:0];
	// Trace: design.sv:102652:3
	assign timeout_ctrl_en_we = (addr_hit[11] & reg_we) & !reg_error;
	// Trace: design.sv:102653:3
	assign timeout_ctrl_en_wd = reg_wdata[31];
	// Trace: design.sv:102656:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:102657:5
		reg_rdata_next = 1'sb0;
		// Trace: design.sv:102658:5
		(* full_case, parallel_case *)
		case (1'b1)
			addr_hit[0]: begin
				// Trace: design.sv:102660:9
				reg_rdata_next[0] = intr_state_tx_watermark_qs;
				// Trace: design.sv:102661:9
				reg_rdata_next[1] = intr_state_rx_watermark_qs;
				// Trace: design.sv:102662:9
				reg_rdata_next[2] = intr_state_tx_empty_qs;
				// Trace: design.sv:102663:9
				reg_rdata_next[3] = intr_state_rx_overflow_qs;
				// Trace: design.sv:102664:9
				reg_rdata_next[4] = intr_state_rx_frame_err_qs;
				// Trace: design.sv:102665:9
				reg_rdata_next[5] = intr_state_rx_break_err_qs;
				// Trace: design.sv:102666:9
				reg_rdata_next[6] = intr_state_rx_timeout_qs;
				// Trace: design.sv:102667:9
				reg_rdata_next[7] = intr_state_rx_parity_err_qs;
			end
			addr_hit[1]: begin
				// Trace: design.sv:102671:9
				reg_rdata_next[0] = intr_enable_tx_watermark_qs;
				// Trace: design.sv:102672:9
				reg_rdata_next[1] = intr_enable_rx_watermark_qs;
				// Trace: design.sv:102673:9
				reg_rdata_next[2] = intr_enable_tx_empty_qs;
				// Trace: design.sv:102674:9
				reg_rdata_next[3] = intr_enable_rx_overflow_qs;
				// Trace: design.sv:102675:9
				reg_rdata_next[4] = intr_enable_rx_frame_err_qs;
				// Trace: design.sv:102676:9
				reg_rdata_next[5] = intr_enable_rx_break_err_qs;
				// Trace: design.sv:102677:9
				reg_rdata_next[6] = intr_enable_rx_timeout_qs;
				// Trace: design.sv:102678:9
				reg_rdata_next[7] = intr_enable_rx_parity_err_qs;
			end
			addr_hit[2]: begin
				// Trace: design.sv:102682:9
				reg_rdata_next[0] = 1'sb0;
				// Trace: design.sv:102683:9
				reg_rdata_next[1] = 1'sb0;
				// Trace: design.sv:102684:9
				reg_rdata_next[2] = 1'sb0;
				// Trace: design.sv:102685:9
				reg_rdata_next[3] = 1'sb0;
				// Trace: design.sv:102686:9
				reg_rdata_next[4] = 1'sb0;
				// Trace: design.sv:102687:9
				reg_rdata_next[5] = 1'sb0;
				// Trace: design.sv:102688:9
				reg_rdata_next[6] = 1'sb0;
				// Trace: design.sv:102689:9
				reg_rdata_next[7] = 1'sb0;
			end
			addr_hit[3]: begin
				// Trace: design.sv:102693:9
				reg_rdata_next[0] = ctrl_tx_qs;
				// Trace: design.sv:102694:9
				reg_rdata_next[1] = ctrl_rx_qs;
				// Trace: design.sv:102695:9
				reg_rdata_next[2] = ctrl_nf_qs;
				// Trace: design.sv:102696:9
				reg_rdata_next[4] = ctrl_slpbk_qs;
				// Trace: design.sv:102697:9
				reg_rdata_next[5] = ctrl_llpbk_qs;
				// Trace: design.sv:102698:9
				reg_rdata_next[6] = ctrl_parity_en_qs;
				// Trace: design.sv:102699:9
				reg_rdata_next[7] = ctrl_parity_odd_qs;
				// Trace: design.sv:102700:9
				reg_rdata_next[9:8] = ctrl_rxblvl_qs;
				// Trace: design.sv:102701:9
				reg_rdata_next[31:16] = ctrl_nco_qs;
			end
			addr_hit[4]: begin
				// Trace: design.sv:102705:9
				reg_rdata_next[0] = status_txfull_qs;
				// Trace: design.sv:102706:9
				reg_rdata_next[1] = status_rxfull_qs;
				// Trace: design.sv:102707:9
				reg_rdata_next[2] = status_txempty_qs;
				// Trace: design.sv:102708:9
				reg_rdata_next[3] = status_txidle_qs;
				// Trace: design.sv:102709:9
				reg_rdata_next[4] = status_rxidle_qs;
				// Trace: design.sv:102710:9
				reg_rdata_next[5] = status_rxempty_qs;
			end
			addr_hit[5]:
				// Trace: design.sv:102714:9
				reg_rdata_next[7:0] = rdata_qs;
			addr_hit[6]:
				// Trace: design.sv:102718:9
				reg_rdata_next[7:0] = 1'sb0;
			addr_hit[7]: begin
				// Trace: design.sv:102722:9
				reg_rdata_next[0] = 1'sb0;
				// Trace: design.sv:102723:9
				reg_rdata_next[1] = 1'sb0;
				// Trace: design.sv:102724:9
				reg_rdata_next[4:2] = fifo_ctrl_rxilvl_qs;
				// Trace: design.sv:102725:9
				reg_rdata_next[6:5] = fifo_ctrl_txilvl_qs;
			end
			addr_hit[8]: begin
				// Trace: design.sv:102729:9
				reg_rdata_next[5:0] = fifo_status_txlvl_qs;
				// Trace: design.sv:102730:9
				reg_rdata_next[21:16] = fifo_status_rxlvl_qs;
			end
			addr_hit[9]: begin
				// Trace: design.sv:102734:9
				reg_rdata_next[0] = ovrd_txen_qs;
				// Trace: design.sv:102735:9
				reg_rdata_next[1] = ovrd_txval_qs;
			end
			addr_hit[10]:
				// Trace: design.sv:102739:9
				reg_rdata_next[15:0] = val_qs;
			addr_hit[11]: begin
				// Trace: design.sv:102743:9
				reg_rdata_next[23:0] = timeout_ctrl_val_qs;
				// Trace: design.sv:102744:9
				reg_rdata_next[31] = timeout_ctrl_en_qs;
			end
			default:
				// Trace: design.sv:102748:9
				reg_rdata_next = 1'sb1;
		endcase
	end
	// Trace: design.sv:102757:3
	wire unused_wdata;
	// Trace: design.sv:102758:3
	wire unused_be;
	// Trace: design.sv:102759:3
	assign unused_wdata = ^reg_wdata;
	// Trace: design.sv:102760:3
	assign unused_be = ^reg_be;
	initial _sv2v_0 = 0;
endmodule
module uart_rx (
	clk_i,
	rst_ni,
	rx_enable,
	tick_baud_x16,
	parity_enable,
	parity_odd,
	tick_baud,
	rx_valid,
	rx_data,
	idle,
	frame_err,
	rx_parity_err,
	rx
);
	reg _sv2v_0;
	// Trace: design.sv:102783:3
	input clk_i;
	// Trace: design.sv:102784:3
	input rst_ni;
	// Trace: design.sv:102786:3
	input rx_enable;
	// Trace: design.sv:102787:3
	input tick_baud_x16;
	// Trace: design.sv:102788:3
	input parity_enable;
	// Trace: design.sv:102789:3
	input parity_odd;
	// Trace: design.sv:102791:3
	output wire tick_baud;
	// Trace: design.sv:102792:3
	output wire rx_valid;
	// Trace: design.sv:102793:3
	output wire [7:0] rx_data;
	// Trace: design.sv:102794:3
	output wire idle;
	// Trace: design.sv:102795:3
	output wire frame_err;
	// Trace: design.sv:102796:3
	output wire rx_parity_err;
	// Trace: design.sv:102798:3
	input rx;
	// Trace: design.sv:102801:3
	reg rx_valid_q;
	// Trace: design.sv:102802:3
	reg [10:0] sreg_q;
	reg [10:0] sreg_d;
	// Trace: design.sv:102803:3
	reg [3:0] bit_cnt_q;
	reg [3:0] bit_cnt_d;
	// Trace: design.sv:102804:3
	reg [3:0] baud_div_q;
	reg [3:0] baud_div_d;
	// Trace: design.sv:102805:3
	reg tick_baud_d;
	reg tick_baud_q;
	// Trace: design.sv:102806:3
	reg idle_d;
	reg idle_q;
	// Trace: design.sv:102808:3
	assign tick_baud = tick_baud_q;
	// Trace: design.sv:102809:3
	assign idle = idle_q;
	// Trace: design.sv:102811:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:102812:5
		if (!rst_ni) begin
			// Trace: design.sv:102813:7
			sreg_q <= 11'h000;
			// Trace: design.sv:102814:7
			bit_cnt_q <= 4'h0;
			// Trace: design.sv:102815:7
			baud_div_q <= 4'h0;
			// Trace: design.sv:102816:7
			tick_baud_q <= 1'b0;
			// Trace: design.sv:102817:7
			idle_q <= 1'b1;
		end
		else begin
			// Trace: design.sv:102819:7
			sreg_q <= sreg_d;
			// Trace: design.sv:102820:7
			bit_cnt_q <= bit_cnt_d;
			// Trace: design.sv:102821:7
			baud_div_q <= baud_div_d;
			// Trace: design.sv:102822:7
			tick_baud_q <= tick_baud_d;
			// Trace: design.sv:102823:7
			idle_q <= idle_d;
		end
	// Trace: design.sv:102827:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:102828:5
		if (!rx_enable) begin
			// Trace: design.sv:102829:7
			sreg_d = 11'h000;
			// Trace: design.sv:102830:7
			bit_cnt_d = 4'h0;
			// Trace: design.sv:102831:7
			baud_div_d = 4'h0;
			// Trace: design.sv:102832:7
			tick_baud_d = 1'b0;
			// Trace: design.sv:102833:7
			idle_d = 1'b1;
		end
		else begin
			// Trace: design.sv:102835:7
			tick_baud_d = 1'b0;
			// Trace: design.sv:102836:7
			sreg_d = sreg_q;
			// Trace: design.sv:102837:7
			bit_cnt_d = bit_cnt_q;
			// Trace: design.sv:102838:7
			baud_div_d = baud_div_q;
			// Trace: design.sv:102839:7
			idle_d = idle_q;
			// Trace: design.sv:102840:7
			if (tick_baud_x16)
				// Trace: design.sv:102841:9
				{tick_baud_d, baud_div_d} = {1'b0, baud_div_q} + 5'h01;
			if (idle_q && !rx) begin
				// Trace: design.sv:102846:9
				baud_div_d = 4'd8;
				// Trace: design.sv:102847:9
				tick_baud_d = 1'b0;
				// Trace: design.sv:102848:9
				bit_cnt_d = (parity_enable ? 4'd11 : 4'd10);
				// Trace: design.sv:102849:9
				sreg_d = 11'h000;
				// Trace: design.sv:102850:9
				idle_d = 1'b0;
			end
			else if (!idle_q && tick_baud_q) begin
				begin
					// Trace: design.sv:102852:9
					if ((bit_cnt_q == (parity_enable ? 4'd11 : 4'd10)) && rx) begin
						// Trace: design.sv:102855:11
						idle_d = 1'b1;
						// Trace: design.sv:102856:11
						bit_cnt_d = 4'h0;
					end
					else begin
						// Trace: design.sv:102858:11
						sreg_d = {rx, sreg_q[10:1]};
						// Trace: design.sv:102859:11
						bit_cnt_d = bit_cnt_q - 4'h1;
						// Trace: design.sv:102860:11
						idle_d = bit_cnt_q == 4'h1;
					end
				end
			end
		end
	end
	// Trace: design.sv:102866:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:102867:5
		if (!rst_ni)
			// Trace: design.sv:102867:18
			rx_valid_q <= 1'b0;
		else
			// Trace: design.sv:102868:18
			rx_valid_q <= tick_baud_q & (bit_cnt_q == 4'h1);
	// Trace: design.sv:102872:3
	assign rx_valid = rx_valid_q;
	// Trace: design.sv:102873:3
	assign rx_data = (parity_enable ? sreg_q[8:1] : sreg_q[9:2]);
	// Trace: design.sv:102875:3
	assign frame_err = rx_valid_q & ~sreg_q[10];
	// Trace: design.sv:102876:3
	assign rx_parity_err = (parity_enable & rx_valid_q) & ^{sreg_q[9:1], parity_odd};
	initial _sv2v_0 = 0;
endmodule
module uart_tx (
	clk_i,
	rst_ni,
	tx_enable,
	tick_baud_x16,
	parity_enable,
	wr,
	wr_parity,
	wr_data,
	idle,
	tx
);
	reg _sv2v_0;
	// Trace: design.sv:102888:3
	input clk_i;
	// Trace: design.sv:102889:3
	input rst_ni;
	// Trace: design.sv:102891:3
	input tx_enable;
	// Trace: design.sv:102892:3
	input tick_baud_x16;
	// Trace: design.sv:102893:3
	input wire parity_enable;
	// Trace: design.sv:102895:3
	input wr;
	// Trace: design.sv:102896:3
	input wire wr_parity;
	// Trace: design.sv:102897:3
	input [7:0] wr_data;
	// Trace: design.sv:102898:3
	output wire idle;
	// Trace: design.sv:102900:3
	output wire tx;
	// Trace: design.sv:102904:3
	reg [3:0] baud_div_q;
	// Trace: design.sv:102905:3
	reg tick_baud_q;
	// Trace: design.sv:102907:3
	reg [3:0] bit_cnt_q;
	reg [3:0] bit_cnt_d;
	// Trace: design.sv:102908:3
	reg [10:0] sreg_q;
	reg [10:0] sreg_d;
	// Trace: design.sv:102909:3
	reg tx_q;
	reg tx_d;
	// Trace: design.sv:102911:3
	assign tx = tx_q;
	// Trace: design.sv:102913:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:102914:5
		if (!rst_ni) begin
			// Trace: design.sv:102915:7
			baud_div_q <= 4'h0;
			// Trace: design.sv:102916:7
			tick_baud_q <= 1'b0;
		end
		else if (tick_baud_x16)
			// Trace: design.sv:102918:7
			{tick_baud_q, baud_div_q} <= {1'b0, baud_div_q} + 5'h01;
		else
			// Trace: design.sv:102920:7
			tick_baud_q <= 1'b0;
	// Trace: design.sv:102924:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:102925:5
		if (!rst_ni) begin
			// Trace: design.sv:102926:7
			bit_cnt_q <= 4'h0;
			// Trace: design.sv:102927:7
			sreg_q <= 11'h7ff;
			// Trace: design.sv:102928:7
			tx_q <= 1'b1;
		end
		else begin
			// Trace: design.sv:102930:7
			bit_cnt_q <= bit_cnt_d;
			// Trace: design.sv:102931:7
			sreg_q <= sreg_d;
			// Trace: design.sv:102932:7
			tx_q <= tx_d;
		end
	// Trace: design.sv:102936:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:102937:5
		if (!tx_enable) begin
			// Trace: design.sv:102938:7
			bit_cnt_d = 4'h0;
			// Trace: design.sv:102939:7
			sreg_d = 11'h7ff;
			// Trace: design.sv:102940:7
			tx_d = 1'b1;
		end
		else begin
			// Trace: design.sv:102942:7
			bit_cnt_d = bit_cnt_q;
			// Trace: design.sv:102943:7
			sreg_d = sreg_q;
			// Trace: design.sv:102944:7
			tx_d = tx_q;
			// Trace: design.sv:102945:7
			if (wr) begin
				// Trace: design.sv:102946:9
				sreg_d = {1'b1, (parity_enable ? wr_parity : 1'b1), wr_data, 1'b0};
				// Trace: design.sv:102947:9
				bit_cnt_d = (parity_enable ? 4'd11 : 4'd10);
			end
			else if (tick_baud_q && (bit_cnt_q != 4'h0)) begin
				// Trace: design.sv:102949:9
				sreg_d = {1'b1, sreg_q[10:1]};
				// Trace: design.sv:102950:9
				tx_d = sreg_q[0];
				// Trace: design.sv:102951:9
				bit_cnt_d = bit_cnt_q - 4'h1;
			end
		end
	end
	// Trace: design.sv:102956:3
	assign idle = (tx_enable ? bit_cnt_q == 4'h0 : 1'b1);
	initial _sv2v_0 = 0;
endmodule
module uart_core (
	clk_i,
	rst_ni,
	reg2hw,
	hw2reg,
	rx,
	tx,
	intr_tx_watermark_o,
	intr_rx_watermark_o,
	intr_tx_empty_o,
	intr_rx_overflow_o,
	intr_rx_frame_err_o,
	intr_rx_break_err_o,
	intr_rx_timeout_o,
	intr_rx_parity_err_o
);
	reg _sv2v_0;
	// Trace: design.sv:102967:3
	input clk_i;
	// Trace: design.sv:102968:3
	input rst_ni;
	// Trace: design.sv:102970:3
	// removed localparam type uart_reg_pkg_uart_reg2hw_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_fifo_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_enable_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_state_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_test_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_ovrd_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_rdata_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_status_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_timeout_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_wdata_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_t
	input wire [124:0] reg2hw;
	// Trace: design.sv:102971:3
	// removed localparam type uart_reg_pkg_uart_hw2reg_fifo_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_fifo_status_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_intr_state_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_rdata_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_status_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_val_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_t
	output wire [64:0] hw2reg;
	// Trace: design.sv:102973:3
	input rx;
	// Trace: design.sv:102974:3
	output wire tx;
	// Trace: design.sv:102976:3
	output wire intr_tx_watermark_o;
	// Trace: design.sv:102977:3
	output wire intr_rx_watermark_o;
	// Trace: design.sv:102978:3
	output wire intr_tx_empty_o;
	// Trace: design.sv:102979:3
	output wire intr_rx_overflow_o;
	// Trace: design.sv:102980:3
	output wire intr_rx_frame_err_o;
	// Trace: design.sv:102981:3
	output wire intr_rx_break_err_o;
	// Trace: design.sv:102982:3
	output wire intr_rx_timeout_o;
	// Trace: design.sv:102983:3
	output wire intr_rx_parity_err_o;
	// Trace: design.sv:102986:3
	// removed import uart_reg_pkg::*;
	// Trace: design.sv:102988:3
	localparam signed [31:0] NcoWidth = 16;
	// Trace: design.sv:102990:3
	reg [15:0] rx_val_q;
	// Trace: design.sv:102991:3
	wire [7:0] uart_rdata;
	// Trace: design.sv:102992:3
	wire tick_baud_x16;
	wire rx_tick_baud;
	// Trace: design.sv:102993:3
	wire [5:0] tx_fifo_depth;
	wire [5:0] rx_fifo_depth;
	// Trace: design.sv:102994:3
	reg [5:0] rx_fifo_depth_prev_q;
	// Trace: design.sv:102995:3
	wire [23:0] rx_timeout_count_d;
	reg [23:0] rx_timeout_count_q;
	wire [23:0] uart_rxto_val;
	// Trace: design.sv:102996:3
	wire rx_fifo_depth_changed;
	wire uart_rxto_en;
	// Trace: design.sv:102997:3
	wire tx_enable;
	wire rx_enable;
	// Trace: design.sv:102998:3
	wire sys_loopback;
	wire line_loopback;
	wire rxnf_enable;
	// Trace: design.sv:102999:3
	wire uart_fifo_rxrst;
	wire uart_fifo_txrst;
	// Trace: design.sv:103000:3
	wire [2:0] uart_fifo_rxilvl;
	// Trace: design.sv:103001:3
	wire [1:0] uart_fifo_txilvl;
	// Trace: design.sv:103002:3
	wire ovrd_tx_en;
	wire ovrd_tx_val;
	// Trace: design.sv:103003:3
	wire [7:0] tx_fifo_data;
	// Trace: design.sv:103004:3
	wire tx_fifo_rready;
	wire tx_fifo_rvalid;
	// Trace: design.sv:103005:3
	wire tx_fifo_wready;
	wire tx_uart_idle;
	// Trace: design.sv:103006:3
	wire tx_out;
	// Trace: design.sv:103007:3
	reg tx_out_q;
	// Trace: design.sv:103008:3
	wire [7:0] rx_fifo_data;
	// Trace: design.sv:103009:3
	wire rx_valid;
	wire rx_fifo_wvalid;
	wire rx_fifo_rvalid;
	// Trace: design.sv:103010:3
	wire rx_fifo_wready;
	wire rx_uart_idle;
	// Trace: design.sv:103011:3
	wire rx_sync;
	// Trace: design.sv:103012:3
	wire rx_in;
	// Trace: design.sv:103013:3
	reg break_err;
	// Trace: design.sv:103014:3
	wire [4:0] allzero_cnt_d;
	reg [4:0] allzero_cnt_q;
	// Trace: design.sv:103015:3
	wire allzero_err;
	wire not_allzero_char;
	// Trace: design.sv:103016:3
	wire event_tx_watermark;
	wire event_rx_watermark;
	wire event_tx_empty;
	wire event_rx_overflow;
	// Trace: design.sv:103017:3
	wire event_rx_frame_err;
	wire event_rx_break_err;
	wire event_rx_timeout;
	wire event_rx_parity_err;
	// Trace: design.sv:103018:3
	reg tx_watermark_d;
	reg tx_watermark_prev_q;
	// Trace: design.sv:103019:3
	reg rx_watermark_d;
	reg rx_watermark_prev_q;
	// Trace: design.sv:103020:3
	reg tx_uart_idle_q;
	// Trace: design.sv:103022:3
	assign tx_enable = reg2hw[92];
	// Trace: design.sv:103023:3
	assign rx_enable = reg2hw[91];
	// Trace: design.sv:103024:3
	assign rxnf_enable = reg2hw[90];
	// Trace: design.sv:103025:3
	assign sys_loopback = reg2hw[89];
	// Trace: design.sv:103026:3
	assign line_loopback = reg2hw[88];
	// Trace: design.sv:103028:3
	assign uart_fifo_rxrst = reg2hw[37] & reg2hw[36];
	// Trace: design.sv:103029:3
	assign uart_fifo_txrst = reg2hw[35] & reg2hw[34];
	// Trace: design.sv:103030:3
	assign uart_fifo_rxilvl = reg2hw[33-:3];
	// Trace: design.sv:103031:3
	assign uart_fifo_txilvl = reg2hw[29-:2];
	// Trace: design.sv:103033:3
	assign ovrd_tx_en = reg2hw[26];
	// Trace: design.sv:103034:3
	assign ovrd_tx_val = reg2hw[25];
	// Trace: design.sv:103036:3
	// removed localparam type break_st_e
	// Trace: design.sv:103041:3
	reg break_st_q;
	// Trace: design.sv:103043:3
	assign not_allzero_char = rx_valid & (~event_rx_frame_err | (rx_fifo_data != 8'h00));
	// Trace: design.sv:103044:3
	assign allzero_err = event_rx_frame_err & (rx_fifo_data == 8'h00);
	// Trace: design.sv:103047:3
	assign allzero_cnt_d = ((break_st_q == 1'd1) || not_allzero_char ? 5'h00 : (allzero_err ? allzero_cnt_q + 5'd1 : allzero_cnt_q));
	// Trace: design.sv:103053:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:103054:5
		if (!rst_ni)
			// Trace: design.sv:103054:25
			allzero_cnt_q <= 1'sb0;
		else if (rx_enable)
			// Trace: design.sv:103055:25
			allzero_cnt_q <= allzero_cnt_d;
	// Trace: design.sv:103061:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:103062:5
		(* full_case, parallel_case *)
		case (reg2hw[85-:2])
			2'h0:
				// Trace: design.sv:103063:16
				break_err = allzero_cnt_d >= 5'd2;
			2'h1:
				// Trace: design.sv:103064:16
				break_err = allzero_cnt_d >= 5'd4;
			2'h2:
				// Trace: design.sv:103065:16
				break_err = allzero_cnt_d >= 5'd8;
			default:
				// Trace: design.sv:103066:16
				break_err = allzero_cnt_d >= 5'd16;
		endcase
	end
	// Trace: design.sv:103070:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:103071:5
		if (!rst_ni)
			// Trace: design.sv:103071:18
			break_st_q <= 1'd0;
		else
			// Trace: design.sv:103073:7
			(* full_case, parallel_case *)
			case (break_st_q)
				1'd0:
					// Trace: design.sv:103075:11
					if (event_rx_break_err)
						// Trace: design.sv:103075:35
						break_st_q <= 1'd1;
				1'd1:
					// Trace: design.sv:103079:11
					if (rx_in)
						// Trace: design.sv:103079:22
						break_st_q <= 1'd0;
				default:
					// Trace: design.sv:103083:11
					break_st_q <= 1'd0;
			endcase
	// Trace: design.sv:103089:3
	assign hw2reg[15-:16] = rx_val_q;
	// Trace: design.sv:103091:3
	assign hw2reg[42-:8] = uart_rdata;
	// Trace: design.sv:103093:3
	assign hw2reg[43] = ~rx_fifo_rvalid;
	// Trace: design.sv:103094:3
	assign hw2reg[44] = rx_uart_idle;
	// Trace: design.sv:103095:3
	assign hw2reg[45] = tx_uart_idle & ~tx_fifo_rvalid;
	// Trace: design.sv:103096:3
	assign hw2reg[46] = ~tx_fifo_rvalid;
	// Trace: design.sv:103097:3
	assign hw2reg[47] = ~rx_fifo_wready;
	// Trace: design.sv:103098:3
	assign hw2reg[48] = ~tx_fifo_wready;
	// Trace: design.sv:103100:3
	assign hw2reg[27-:6] = tx_fifo_depth;
	// Trace: design.sv:103101:3
	assign hw2reg[21-:6] = rx_fifo_depth;
	// Trace: design.sv:103104:3
	assign hw2reg[31] = 1'b0;
	// Trace: design.sv:103105:3
	assign hw2reg[34-:3] = 3'h0;
	// Trace: design.sv:103106:3
	assign hw2reg[28] = 1'b0;
	// Trace: design.sv:103107:3
	assign hw2reg[30-:2] = 2'h0;
	// Trace: design.sv:103112:3
	reg [NcoWidth:0] nco_sum_q;
	// Trace: design.sv:103114:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:103115:5
		if (!rst_ni)
			// Trace: design.sv:103116:7
			nco_sum_q <= 17'h00000;
		else if (tx_enable || rx_enable)
			// Trace: design.sv:103118:7
			nco_sum_q <= {1'b0, nco_sum_q[15:0]} + {1'b0, reg2hw[83:68]};
	// Trace: design.sv:103122:3
	assign tick_baud_x16 = nco_sum_q[16];
	// Trace: design.sv:103128:3
	assign tx_fifo_rready = (tx_uart_idle & tx_fifo_rvalid) & tx_enable;
	// Trace: design.sv:103130:3
	prim_fifo_sync #(
		.Width(8),
		.Pass(1'b0),
		.Depth(32)
	) u_uart_txfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(uart_fifo_txrst),
		.wvalid_i(reg2hw[38]),
		.wready_o(tx_fifo_wready),
		.wdata_i(reg2hw[46-:8]),
		.depth_o(tx_fifo_depth),
		.full_o(),
		.rvalid_o(tx_fifo_rvalid),
		.rready_i(tx_fifo_rready),
		.rdata_o(tx_fifo_data)
	);
	// Trace: design.sv:103148:3
	uart_tx uart_tx(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tx_enable(tx_enable),
		.tick_baud_x16(tick_baud_x16),
		.parity_enable(reg2hw[87]),
		.wr(tx_fifo_rready),
		.wr_parity(^tx_fifo_data ^ reg2hw[86]),
		.wr_data(tx_fifo_data),
		.idle(tx_uart_idle),
		.tx(tx_out)
	);
	// Trace: design.sv:103161:3
	assign tx = (line_loopback ? rx : tx_out_q);
	// Trace: design.sv:103162:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:103163:5
		if (!rst_ni)
			// Trace: design.sv:103164:7
			tx_out_q <= 1'b1;
		else if (ovrd_tx_en)
			// Trace: design.sv:103166:7
			tx_out_q <= ovrd_tx_val;
		else if (sys_loopback)
			// Trace: design.sv:103168:7
			tx_out_q <= 1'b1;
		else
			// Trace: design.sv:103170:7
			tx_out_q <= tx_out;
	// Trace: design.sv:103179:3
	prim_flop_2sync #(
		.Width(1),
		.ResetValue(1'b1)
	) sync_rx(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(rx),
		.q_o(rx_sync)
	);
	// Trace: design.sv:103191:3
	reg rx_sync_q1;
	reg rx_sync_q2;
	wire rx_in_mx;
	wire rx_in_maj;
	// Trace: design.sv:103193:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:103194:5
		if (!rst_ni) begin
			// Trace: design.sv:103195:7
			rx_sync_q1 <= 1'b1;
			// Trace: design.sv:103196:7
			rx_sync_q2 <= 1'b1;
		end
		else begin
			// Trace: design.sv:103198:7
			rx_sync_q1 <= rx_sync;
			// Trace: design.sv:103199:7
			rx_sync_q2 <= rx_sync_q1;
		end
	// Trace: design.sv:103203:3
	assign rx_in_maj = ((rx_sync & rx_sync_q1) | (rx_sync & rx_sync_q2)) | (rx_sync_q1 & rx_sync_q2);
	// Trace: design.sv:103206:3
	assign rx_in_mx = (rxnf_enable ? rx_in_maj : rx_sync);
	// Trace: design.sv:103208:3
	assign rx_in = (sys_loopback ? tx_out : (line_loopback ? 1'b1 : rx_in_mx));
	// Trace: design.sv:103212:3
	uart_rx uart_rx(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rx_enable(rx_enable),
		.tick_baud_x16(tick_baud_x16),
		.parity_enable(reg2hw[87]),
		.parity_odd(reg2hw[86]),
		.tick_baud(rx_tick_baud),
		.rx_valid(rx_valid),
		.rx_data(rx_fifo_data),
		.idle(rx_uart_idle),
		.frame_err(event_rx_frame_err),
		.rx(rx_in),
		.rx_parity_err(event_rx_parity_err)
	);
	// Trace: design.sv:103228:3
	assign rx_fifo_wvalid = (rx_valid & ~event_rx_frame_err) & ~event_rx_parity_err;
	// Trace: design.sv:103230:3
	prim_fifo_sync #(
		.Width(8),
		.Pass(1'b0),
		.Depth(32)
	) u_uart_rxfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(uart_fifo_rxrst),
		.wvalid_i(rx_fifo_wvalid),
		.wready_o(rx_fifo_wready),
		.wdata_i(rx_fifo_data),
		.depth_o(rx_fifo_depth),
		.full_o(),
		.rvalid_o(rx_fifo_rvalid),
		.rready_i(reg2hw[47]),
		.rdata_o(uart_rdata)
	);
	// Trace: design.sv:103248:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:103249:5
		if (!rst_ni)
			// Trace: design.sv:103249:29
			rx_val_q <= 16'h0000;
		else if (tick_baud_x16)
			// Trace: design.sv:103250:29
			rx_val_q <= {rx_val_q[14:0], rx_in};
	// Trace: design.sv:103257:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:103258:5
		(* full_case, parallel_case *)
		case (uart_fifo_txilvl)
			2'h0:
				// Trace: design.sv:103259:16
				tx_watermark_d = tx_fifo_depth < 6'd2;
			2'h1:
				// Trace: design.sv:103260:16
				tx_watermark_d = tx_fifo_depth < 6'd4;
			2'h2:
				// Trace: design.sv:103261:16
				tx_watermark_d = tx_fifo_depth < 6'd8;
			default:
				// Trace: design.sv:103262:16
				tx_watermark_d = tx_fifo_depth < 6'd16;
		endcase
	end
	// Trace: design.sv:103266:3
	assign event_tx_watermark = tx_watermark_d & ~tx_watermark_prev_q;
	// Trace: design.sv:103278:3
	assign event_tx_empty = (~tx_fifo_rvalid & ~tx_uart_idle_q) & tx_uart_idle;
	// Trace: design.sv:103280:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:103281:5
		if (!rst_ni) begin
			// Trace: design.sv:103282:7
			tx_watermark_prev_q <= 1'b1;
			// Trace: design.sv:103283:7
			rx_watermark_prev_q <= 1'b0;
			// Trace: design.sv:103284:7
			tx_uart_idle_q <= 1'b1;
		end
		else begin
			// Trace: design.sv:103286:7
			tx_watermark_prev_q <= tx_watermark_d;
			// Trace: design.sv:103287:7
			rx_watermark_prev_q <= rx_watermark_d;
			// Trace: design.sv:103288:7
			tx_uart_idle_q <= tx_uart_idle;
		end
	// Trace: design.sv:103292:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:103293:5
		(* full_case, parallel_case *)
		case (uart_fifo_rxilvl)
			3'h0:
				// Trace: design.sv:103294:16
				rx_watermark_d = rx_fifo_depth >= 6'd1;
			3'h1:
				// Trace: design.sv:103295:16
				rx_watermark_d = rx_fifo_depth >= 6'd4;
			3'h2:
				// Trace: design.sv:103296:16
				rx_watermark_d = rx_fifo_depth >= 6'd8;
			3'h3:
				// Trace: design.sv:103297:16
				rx_watermark_d = rx_fifo_depth >= 6'd16;
			3'h4:
				// Trace: design.sv:103298:16
				rx_watermark_d = rx_fifo_depth >= 6'd30;
			default:
				// Trace: design.sv:103299:16
				rx_watermark_d = 1'b0;
		endcase
	end
	// Trace: design.sv:103303:3
	assign event_rx_watermark = rx_watermark_d & ~rx_watermark_prev_q;
	// Trace: design.sv:103306:3
	assign uart_rxto_en = reg2hw[0];
	// Trace: design.sv:103307:3
	assign uart_rxto_val = reg2hw[24-:24];
	// Trace: design.sv:103309:3
	assign rx_fifo_depth_changed = rx_fifo_depth != rx_fifo_depth_prev_q;
	// Trace: design.sv:103311:3
	assign rx_timeout_count_d = (uart_rxto_en == 1'b0 ? 24'd0 : (event_rx_timeout ? 24'd0 : (rx_fifo_depth_changed ? 24'd0 : (rx_fifo_depth == {6 {1'sb0}} ? 24'd0 : (rx_tick_baud ? rx_timeout_count_q + 24'd1 : rx_timeout_count_q)))));
	// Trace: design.sv:103329:3
	assign event_rx_timeout = (rx_timeout_count_q == uart_rxto_val) & uart_rxto_en;
	// Trace: design.sv:103331:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: design.sv:103332:5
		if (!rst_ni) begin
			// Trace: design.sv:103333:7
			rx_timeout_count_q <= 24'd0;
			// Trace: design.sv:103334:7
			rx_fifo_depth_prev_q <= 6'd0;
		end
		else begin
			// Trace: design.sv:103336:7
			rx_timeout_count_q <= rx_timeout_count_d;
			// Trace: design.sv:103337:7
			rx_fifo_depth_prev_q <= rx_fifo_depth;
		end
	// Trace: design.sv:103341:3
	assign event_rx_overflow = rx_fifo_wvalid & ~rx_fifo_wready;
	// Trace: design.sv:103342:3
	assign event_rx_break_err = break_err & (break_st_q == 1'd0);
	// Trace: design.sv:103346:3
	prim_intr_hw #(.Width(1)) intr_hw_tx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_tx_watermark),
		.reg2hw_intr_enable_q_i(reg2hw[116]),
		.reg2hw_intr_test_q_i(reg2hw[108]),
		.reg2hw_intr_test_qe_i(reg2hw[107]),
		.reg2hw_intr_state_q_i(reg2hw[124]),
		.hw2reg_intr_state_de_o(hw2reg[63]),
		.hw2reg_intr_state_d_o(hw2reg[64]),
		.intr_o(intr_tx_watermark_o)
	);
	// Trace: design.sv:103359:3
	prim_intr_hw #(.Width(1)) intr_hw_rx_watermark(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_rx_watermark),
		.reg2hw_intr_enable_q_i(reg2hw[115]),
		.reg2hw_intr_test_q_i(reg2hw[106]),
		.reg2hw_intr_test_qe_i(reg2hw[105]),
		.reg2hw_intr_state_q_i(reg2hw[123]),
		.hw2reg_intr_state_de_o(hw2reg[61]),
		.hw2reg_intr_state_d_o(hw2reg[62]),
		.intr_o(intr_rx_watermark_o)
	);
	// Trace: design.sv:103372:3
	prim_intr_hw #(.Width(1)) intr_hw_tx_empty(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_tx_empty),
		.reg2hw_intr_enable_q_i(reg2hw[114]),
		.reg2hw_intr_test_q_i(reg2hw[104]),
		.reg2hw_intr_test_qe_i(reg2hw[103]),
		.reg2hw_intr_state_q_i(reg2hw[122]),
		.hw2reg_intr_state_de_o(hw2reg[59]),
		.hw2reg_intr_state_d_o(hw2reg[60]),
		.intr_o(intr_tx_empty_o)
	);
	// Trace: design.sv:103385:3
	prim_intr_hw #(.Width(1)) intr_hw_rx_overflow(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_rx_overflow),
		.reg2hw_intr_enable_q_i(reg2hw[113]),
		.reg2hw_intr_test_q_i(reg2hw[102]),
		.reg2hw_intr_test_qe_i(reg2hw[101]),
		.reg2hw_intr_state_q_i(reg2hw[121]),
		.hw2reg_intr_state_de_o(hw2reg[57]),
		.hw2reg_intr_state_d_o(hw2reg[58]),
		.intr_o(intr_rx_overflow_o)
	);
	// Trace: design.sv:103398:3
	prim_intr_hw #(.Width(1)) intr_hw_rx_frame_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_rx_frame_err),
		.reg2hw_intr_enable_q_i(reg2hw[112]),
		.reg2hw_intr_test_q_i(reg2hw[100]),
		.reg2hw_intr_test_qe_i(reg2hw[99]),
		.reg2hw_intr_state_q_i(reg2hw[120]),
		.hw2reg_intr_state_de_o(hw2reg[55]),
		.hw2reg_intr_state_d_o(hw2reg[56]),
		.intr_o(intr_rx_frame_err_o)
	);
	// Trace: design.sv:103411:3
	prim_intr_hw #(.Width(1)) intr_hw_rx_break_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_rx_break_err),
		.reg2hw_intr_enable_q_i(reg2hw[111]),
		.reg2hw_intr_test_q_i(reg2hw[98]),
		.reg2hw_intr_test_qe_i(reg2hw[97]),
		.reg2hw_intr_state_q_i(reg2hw[119]),
		.hw2reg_intr_state_de_o(hw2reg[53]),
		.hw2reg_intr_state_d_o(hw2reg[54]),
		.intr_o(intr_rx_break_err_o)
	);
	// Trace: design.sv:103424:3
	prim_intr_hw #(.Width(1)) intr_hw_rx_timeout(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_rx_timeout),
		.reg2hw_intr_enable_q_i(reg2hw[110]),
		.reg2hw_intr_test_q_i(reg2hw[96]),
		.reg2hw_intr_test_qe_i(reg2hw[95]),
		.reg2hw_intr_state_q_i(reg2hw[118]),
		.hw2reg_intr_state_de_o(hw2reg[51]),
		.hw2reg_intr_state_d_o(hw2reg[52]),
		.intr_o(intr_rx_timeout_o)
	);
	// Trace: design.sv:103437:3
	prim_intr_hw #(.Width(1)) intr_hw_rx_parity_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.event_intr_i(event_rx_parity_err),
		.reg2hw_intr_enable_q_i(reg2hw[109]),
		.reg2hw_intr_test_q_i(reg2hw[94]),
		.reg2hw_intr_test_qe_i(reg2hw[93]),
		.reg2hw_intr_state_q_i(reg2hw[117]),
		.hw2reg_intr_state_de_o(hw2reg[49]),
		.hw2reg_intr_state_d_o(hw2reg[50]),
		.intr_o(intr_rx_parity_err_o)
	);
	initial _sv2v_0 = 0;
endmodule
module uart (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	cio_rx_i,
	cio_tx_o,
	cio_tx_en_o,
	intr_tx_watermark_o,
	intr_rx_watermark_o,
	intr_tx_empty_o,
	intr_rx_overflow_o,
	intr_rx_frame_err_o,
	intr_rx_break_err_o,
	intr_rx_timeout_o,
	intr_rx_parity_err_o
);
	// Trace: design.sv:103460:3
	input clk_i;
	// Trace: design.sv:103461:3
	input rst_ni;
	// Trace: design.sv:103464:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] tl_i;
	// Trace: design.sv:103465:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	// Trace: design.sv:103468:3
	input cio_rx_i;
	// Trace: design.sv:103469:3
	output wire cio_tx_o;
	// Trace: design.sv:103470:3
	output wire cio_tx_en_o;
	// Trace: design.sv:103473:3
	output wire intr_tx_watermark_o;
	// Trace: design.sv:103474:3
	output wire intr_rx_watermark_o;
	// Trace: design.sv:103475:3
	output wire intr_tx_empty_o;
	// Trace: design.sv:103476:3
	output wire intr_rx_overflow_o;
	// Trace: design.sv:103477:3
	output wire intr_rx_frame_err_o;
	// Trace: design.sv:103478:3
	output wire intr_rx_break_err_o;
	// Trace: design.sv:103479:3
	output wire intr_rx_timeout_o;
	// Trace: design.sv:103480:3
	output wire intr_rx_parity_err_o;
	// Trace: design.sv:103483:3
	// removed import uart_reg_pkg::*;
	// Trace: design.sv:103485:3
	// removed localparam type uart_reg_pkg_uart_reg2hw_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_fifo_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_enable_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_state_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_intr_test_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_ovrd_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_rdata_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_status_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_timeout_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_wdata_reg_t
	// removed localparam type uart_reg_pkg_uart_reg2hw_t
	wire [124:0] reg2hw;
	// Trace: design.sv:103486:3
	// removed localparam type uart_reg_pkg_uart_hw2reg_fifo_ctrl_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_fifo_status_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_intr_state_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_rdata_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_status_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_val_reg_t
	// removed localparam type uart_reg_pkg_uart_hw2reg_t
	wire [64:0] hw2reg;
	// Trace: design.sv:103488:3
	uart_reg_top u_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.tl_o(tl_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.intg_err_o(),
		.devmode_i(1'b1)
	);
	// Trace: design.sv:103499:3
	uart_core uart_core(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.rx(cio_rx_i),
		.tx(cio_tx_o),
		.intr_tx_watermark_o(intr_tx_watermark_o),
		.intr_rx_watermark_o(intr_rx_watermark_o),
		.intr_tx_empty_o(intr_tx_empty_o),
		.intr_rx_overflow_o(intr_rx_overflow_o),
		.intr_rx_frame_err_o(intr_rx_frame_err_o),
		.intr_rx_break_err_o(intr_rx_break_err_o),
		.intr_rx_timeout_o(intr_rx_timeout_o),
		.intr_rx_parity_err_o(intr_rx_parity_err_o)
	);
	// Trace: design.sv:103519:3
	assign cio_tx_en_o = 1'b1;
endmodule
module core_v_mini_mcu (
	rst_ni,
	clk_i,
	boot_select_i,
	execute_from_flash_i,
	jtag_tck_i,
	jtag_tms_i,
	jtag_trst_ni,
	jtag_tdi_i,
	jtag_tdo_o,
	uart_rx_i,
	uart_tx_o,
	exit_valid_o,
	gpio_0_o,
	gpio_0_i,
	gpio_0_oe_o,
	gpio_1_o,
	gpio_1_i,
	gpio_1_oe_o,
	gpio_2_o,
	gpio_2_i,
	gpio_2_oe_o,
	gpio_3_o,
	gpio_3_i,
	gpio_3_oe_o,
	gpio_4_o,
	gpio_4_i,
	gpio_4_oe_o,
	gpio_5_o,
	gpio_5_i,
	gpio_5_oe_o,
	gpio_6_o,
	gpio_6_i,
	gpio_6_oe_o,
	gpio_7_o,
	gpio_7_i,
	gpio_7_oe_o,
	gpio_8_o,
	gpio_8_i,
	gpio_8_oe_o,
	gpio_9_o,
	gpio_9_i,
	gpio_9_oe_o,
	gpio_10_o,
	gpio_10_i,
	gpio_10_oe_o,
	gpio_11_o,
	gpio_11_i,
	gpio_11_oe_o,
	gpio_12_o,
	gpio_12_i,
	gpio_12_oe_o,
	gpio_13_o,
	gpio_13_i,
	gpio_13_oe_o,
	gpio_14_o,
	gpio_14_i,
	gpio_14_oe_o,
	gpio_15_o,
	gpio_15_i,
	gpio_15_oe_o,
	gpio_16_o,
	gpio_16_i,
	gpio_16_oe_o,
	gpio_17_o,
	gpio_17_i,
	gpio_17_oe_o,
	gpio_18_o,
	gpio_18_i,
	gpio_18_oe_o,
	gpio_19_o,
	gpio_19_i,
	gpio_19_oe_o,
	gpio_20_o,
	gpio_20_i,
	gpio_20_oe_o,
	gpio_21_o,
	gpio_21_i,
	gpio_21_oe_o,
	gpio_22_o,
	gpio_22_i,
	gpio_22_oe_o,
	spi_flash_sck_o,
	spi_flash_sck_i,
	spi_flash_sck_oe_o,
	spi_flash_cs_0_o,
	spi_flash_cs_0_i,
	spi_flash_cs_0_oe_o,
	spi_flash_cs_1_o,
	spi_flash_cs_1_i,
	spi_flash_cs_1_oe_o,
	spi_flash_sd_0_o,
	spi_flash_sd_0_i,
	spi_flash_sd_0_oe_o,
	spi_flash_sd_1_o,
	spi_flash_sd_1_i,
	spi_flash_sd_1_oe_o,
	spi_flash_sd_2_o,
	spi_flash_sd_2_i,
	spi_flash_sd_2_oe_o,
	spi_flash_sd_3_o,
	spi_flash_sd_3_i,
	spi_flash_sd_3_oe_o,
	spi_sck_o,
	spi_sck_i,
	spi_sck_oe_o,
	spi_cs_0_o,
	spi_cs_0_i,
	spi_cs_0_oe_o,
	spi_cs_1_o,
	spi_cs_1_i,
	spi_cs_1_oe_o,
	spi_sd_0_o,
	spi_sd_0_i,
	spi_sd_0_oe_o,
	spi_sd_1_o,
	spi_sd_1_i,
	spi_sd_1_oe_o,
	spi_sd_2_o,
	spi_sd_2_i,
	spi_sd_2_oe_o,
	spi_sd_3_o,
	spi_sd_3_i,
	spi_sd_3_oe_o,
	spi2_cs_0_o,
	spi2_cs_0_i,
	spi2_cs_0_oe_o,
	gpio_23_o,
	gpio_23_i,
	gpio_23_oe_o,
	spi2_cs_1_o,
	spi2_cs_1_i,
	spi2_cs_1_oe_o,
	gpio_24_o,
	gpio_24_i,
	gpio_24_oe_o,
	spi2_sck_o,
	spi2_sck_i,
	spi2_sck_oe_o,
	gpio_25_o,
	gpio_25_i,
	gpio_25_oe_o,
	spi2_sd_0_o,
	spi2_sd_0_i,
	spi2_sd_0_oe_o,
	gpio_26_o,
	gpio_26_i,
	gpio_26_oe_o,
	spi2_sd_1_o,
	spi2_sd_1_i,
	spi2_sd_1_oe_o,
	gpio_27_o,
	gpio_27_i,
	gpio_27_oe_o,
	spi2_sd_2_o,
	spi2_sd_2_i,
	spi2_sd_2_oe_o,
	gpio_28_o,
	gpio_28_i,
	gpio_28_oe_o,
	spi2_sd_3_o,
	spi2_sd_3_i,
	spi2_sd_3_oe_o,
	gpio_29_o,
	gpio_29_i,
	gpio_29_oe_o,
	i2c_scl_o,
	i2c_scl_i,
	i2c_scl_oe_o,
	gpio_31_o,
	gpio_31_i,
	gpio_31_oe_o,
	i2c_sda_o,
	i2c_sda_i,
	i2c_sda_oe_o,
	gpio_30_o,
	gpio_30_i,
	gpio_30_oe_o,
	pad_req_o,
	pad_resp_i,
	ext_xbar_master_req_i,
	ext_xbar_master_resp_o,
	ext_xbar_slave_req_o,
	ext_xbar_slave_resp_i,
	ext_peripheral_slave_req_o,
	ext_peripheral_slave_resp_i,
	intr_vector_ext_i,
	cpu_subsystem_powergate_switch_o,
	cpu_subsystem_powergate_switch_ack_i,
	peripheral_subsystem_powergate_switch_o,
	peripheral_subsystem_powergate_switch_ack_i,
	memory_subsystem_banks_powergate_switch_o,
	memory_subsystem_banks_powergate_switch_ack_i,
	external_subsystem_powergate_switch_o,
	external_subsystem_powergate_switch_ack_i,
	external_subsystem_powergate_iso_o,
	external_subsystem_rst_no,
	external_ram_banks_set_retentive_o,
	exit_value_o
);
	// removed import obi_pkg::*;
	// removed import reg_pkg::*;
	// Trace: design.sv:103544:15
	parameter PULP_XPULP = 0;
	// Trace: design.sv:103545:15
	parameter FPU = 0;
	// Trace: design.sv:103546:15
	parameter PULP_ZFINX = 0;
	// Trace: design.sv:103547:15
	parameter EXT_XBAR_NMASTER = 0;
	// Trace: design.sv:103548:15
	parameter X_EXT = 0;
	// Trace: design.sv:103551:5
	input wire rst_ni;
	// Trace: design.sv:103553:9
	input wire clk_i;
	// Trace: design.sv:103556:9
	input wire boot_select_i;
	// Trace: design.sv:103558:9
	input wire execute_from_flash_i;
	// Trace: design.sv:103560:9
	input wire jtag_tck_i;
	// Trace: design.sv:103562:9
	input wire jtag_tms_i;
	// Trace: design.sv:103564:9
	input wire jtag_trst_ni;
	// Trace: design.sv:103566:9
	input wire jtag_tdi_i;
	// Trace: design.sv:103568:9
	output wire jtag_tdo_o;
	// Trace: design.sv:103570:9
	input wire uart_rx_i;
	// Trace: design.sv:103572:9
	output wire uart_tx_o;
	// Trace: design.sv:103574:9
	output wire exit_valid_o;
	// Trace: design.sv:103576:9
	output wire gpio_0_o;
	// Trace: design.sv:103577:5
	input wire gpio_0_i;
	// Trace: design.sv:103578:5
	output wire gpio_0_oe_o;
	// Trace: design.sv:103580:9
	output wire gpio_1_o;
	// Trace: design.sv:103581:5
	input wire gpio_1_i;
	// Trace: design.sv:103582:5
	output wire gpio_1_oe_o;
	// Trace: design.sv:103584:9
	output wire gpio_2_o;
	// Trace: design.sv:103585:5
	input wire gpio_2_i;
	// Trace: design.sv:103586:5
	output wire gpio_2_oe_o;
	// Trace: design.sv:103588:9
	output wire gpio_3_o;
	// Trace: design.sv:103589:5
	input wire gpio_3_i;
	// Trace: design.sv:103590:5
	output wire gpio_3_oe_o;
	// Trace: design.sv:103592:9
	output wire gpio_4_o;
	// Trace: design.sv:103593:5
	input wire gpio_4_i;
	// Trace: design.sv:103594:5
	output wire gpio_4_oe_o;
	// Trace: design.sv:103596:9
	output wire gpio_5_o;
	// Trace: design.sv:103597:5
	input wire gpio_5_i;
	// Trace: design.sv:103598:5
	output wire gpio_5_oe_o;
	// Trace: design.sv:103600:9
	output wire gpio_6_o;
	// Trace: design.sv:103601:5
	input wire gpio_6_i;
	// Trace: design.sv:103602:5
	output wire gpio_6_oe_o;
	// Trace: design.sv:103604:9
	output wire gpio_7_o;
	// Trace: design.sv:103605:5
	input wire gpio_7_i;
	// Trace: design.sv:103606:5
	output wire gpio_7_oe_o;
	// Trace: design.sv:103608:9
	output wire gpio_8_o;
	// Trace: design.sv:103609:5
	input wire gpio_8_i;
	// Trace: design.sv:103610:5
	output wire gpio_8_oe_o;
	// Trace: design.sv:103612:9
	output wire gpio_9_o;
	// Trace: design.sv:103613:5
	input wire gpio_9_i;
	// Trace: design.sv:103614:5
	output wire gpio_9_oe_o;
	// Trace: design.sv:103616:9
	output wire gpio_10_o;
	// Trace: design.sv:103617:5
	input wire gpio_10_i;
	// Trace: design.sv:103618:5
	output wire gpio_10_oe_o;
	// Trace: design.sv:103620:9
	output wire gpio_11_o;
	// Trace: design.sv:103621:5
	input wire gpio_11_i;
	// Trace: design.sv:103622:5
	output wire gpio_11_oe_o;
	// Trace: design.sv:103624:9
	output wire gpio_12_o;
	// Trace: design.sv:103625:5
	input wire gpio_12_i;
	// Trace: design.sv:103626:5
	output wire gpio_12_oe_o;
	// Trace: design.sv:103628:9
	output wire gpio_13_o;
	// Trace: design.sv:103629:5
	input wire gpio_13_i;
	// Trace: design.sv:103630:5
	output wire gpio_13_oe_o;
	// Trace: design.sv:103632:9
	output wire gpio_14_o;
	// Trace: design.sv:103633:5
	input wire gpio_14_i;
	// Trace: design.sv:103634:5
	output wire gpio_14_oe_o;
	// Trace: design.sv:103636:9
	output wire gpio_15_o;
	// Trace: design.sv:103637:5
	input wire gpio_15_i;
	// Trace: design.sv:103638:5
	output wire gpio_15_oe_o;
	// Trace: design.sv:103640:9
	output wire gpio_16_o;
	// Trace: design.sv:103641:5
	input wire gpio_16_i;
	// Trace: design.sv:103642:5
	output wire gpio_16_oe_o;
	// Trace: design.sv:103644:9
	output wire gpio_17_o;
	// Trace: design.sv:103645:5
	input wire gpio_17_i;
	// Trace: design.sv:103646:5
	output wire gpio_17_oe_o;
	// Trace: design.sv:103648:9
	output wire gpio_18_o;
	// Trace: design.sv:103649:5
	input wire gpio_18_i;
	// Trace: design.sv:103650:5
	output wire gpio_18_oe_o;
	// Trace: design.sv:103652:9
	output wire gpio_19_o;
	// Trace: design.sv:103653:5
	input wire gpio_19_i;
	// Trace: design.sv:103654:5
	output wire gpio_19_oe_o;
	// Trace: design.sv:103656:9
	output wire gpio_20_o;
	// Trace: design.sv:103657:5
	input wire gpio_20_i;
	// Trace: design.sv:103658:5
	output wire gpio_20_oe_o;
	// Trace: design.sv:103660:9
	output wire gpio_21_o;
	// Trace: design.sv:103661:5
	input wire gpio_21_i;
	// Trace: design.sv:103662:5
	output wire gpio_21_oe_o;
	// Trace: design.sv:103664:9
	output wire gpio_22_o;
	// Trace: design.sv:103665:5
	input wire gpio_22_i;
	// Trace: design.sv:103666:5
	output wire gpio_22_oe_o;
	// Trace: design.sv:103668:9
	output wire spi_flash_sck_o;
	// Trace: design.sv:103669:5
	input wire spi_flash_sck_i;
	// Trace: design.sv:103670:5
	output wire spi_flash_sck_oe_o;
	// Trace: design.sv:103672:9
	output wire spi_flash_cs_0_o;
	// Trace: design.sv:103673:5
	input wire spi_flash_cs_0_i;
	// Trace: design.sv:103674:5
	output wire spi_flash_cs_0_oe_o;
	// Trace: design.sv:103676:9
	output wire spi_flash_cs_1_o;
	// Trace: design.sv:103677:5
	input wire spi_flash_cs_1_i;
	// Trace: design.sv:103678:5
	output wire spi_flash_cs_1_oe_o;
	// Trace: design.sv:103680:9
	output wire spi_flash_sd_0_o;
	// Trace: design.sv:103681:5
	input wire spi_flash_sd_0_i;
	// Trace: design.sv:103682:5
	output wire spi_flash_sd_0_oe_o;
	// Trace: design.sv:103684:9
	output wire spi_flash_sd_1_o;
	// Trace: design.sv:103685:5
	input wire spi_flash_sd_1_i;
	// Trace: design.sv:103686:5
	output wire spi_flash_sd_1_oe_o;
	// Trace: design.sv:103688:9
	output wire spi_flash_sd_2_o;
	// Trace: design.sv:103689:5
	input wire spi_flash_sd_2_i;
	// Trace: design.sv:103690:5
	output wire spi_flash_sd_2_oe_o;
	// Trace: design.sv:103692:9
	output wire spi_flash_sd_3_o;
	// Trace: design.sv:103693:5
	input wire spi_flash_sd_3_i;
	// Trace: design.sv:103694:5
	output wire spi_flash_sd_3_oe_o;
	// Trace: design.sv:103696:9
	output wire spi_sck_o;
	// Trace: design.sv:103697:5
	input wire spi_sck_i;
	// Trace: design.sv:103698:5
	output wire spi_sck_oe_o;
	// Trace: design.sv:103700:9
	output wire spi_cs_0_o;
	// Trace: design.sv:103701:5
	input wire spi_cs_0_i;
	// Trace: design.sv:103702:5
	output wire spi_cs_0_oe_o;
	// Trace: design.sv:103704:9
	output wire spi_cs_1_o;
	// Trace: design.sv:103705:5
	input wire spi_cs_1_i;
	// Trace: design.sv:103706:5
	output wire spi_cs_1_oe_o;
	// Trace: design.sv:103708:9
	output wire spi_sd_0_o;
	// Trace: design.sv:103709:5
	input wire spi_sd_0_i;
	// Trace: design.sv:103710:5
	output wire spi_sd_0_oe_o;
	// Trace: design.sv:103712:9
	output wire spi_sd_1_o;
	// Trace: design.sv:103713:5
	input wire spi_sd_1_i;
	// Trace: design.sv:103714:5
	output wire spi_sd_1_oe_o;
	// Trace: design.sv:103716:9
	output wire spi_sd_2_o;
	// Trace: design.sv:103717:5
	input wire spi_sd_2_i;
	// Trace: design.sv:103718:5
	output wire spi_sd_2_oe_o;
	// Trace: design.sv:103720:9
	output wire spi_sd_3_o;
	// Trace: design.sv:103721:5
	input wire spi_sd_3_i;
	// Trace: design.sv:103722:5
	output wire spi_sd_3_oe_o;
	// Trace: design.sv:103724:9
	output wire spi2_cs_0_o;
	// Trace: design.sv:103725:5
	input wire spi2_cs_0_i;
	// Trace: design.sv:103726:5
	output wire spi2_cs_0_oe_o;
	// Trace: design.sv:103727:5
	output wire gpio_23_o;
	// Trace: design.sv:103728:5
	input wire gpio_23_i;
	// Trace: design.sv:103729:5
	output wire gpio_23_oe_o;
	// Trace: design.sv:103731:9
	output wire spi2_cs_1_o;
	// Trace: design.sv:103732:5
	input wire spi2_cs_1_i;
	// Trace: design.sv:103733:5
	output wire spi2_cs_1_oe_o;
	// Trace: design.sv:103734:5
	output wire gpio_24_o;
	// Trace: design.sv:103735:5
	input wire gpio_24_i;
	// Trace: design.sv:103736:5
	output wire gpio_24_oe_o;
	// Trace: design.sv:103738:9
	output wire spi2_sck_o;
	// Trace: design.sv:103739:5
	input wire spi2_sck_i;
	// Trace: design.sv:103740:5
	output wire spi2_sck_oe_o;
	// Trace: design.sv:103741:5
	output wire gpio_25_o;
	// Trace: design.sv:103742:5
	input wire gpio_25_i;
	// Trace: design.sv:103743:5
	output wire gpio_25_oe_o;
	// Trace: design.sv:103745:9
	output wire spi2_sd_0_o;
	// Trace: design.sv:103746:5
	input wire spi2_sd_0_i;
	// Trace: design.sv:103747:5
	output wire spi2_sd_0_oe_o;
	// Trace: design.sv:103748:5
	output wire gpio_26_o;
	// Trace: design.sv:103749:5
	input wire gpio_26_i;
	// Trace: design.sv:103750:5
	output wire gpio_26_oe_o;
	// Trace: design.sv:103752:9
	output wire spi2_sd_1_o;
	// Trace: design.sv:103753:5
	input wire spi2_sd_1_i;
	// Trace: design.sv:103754:5
	output wire spi2_sd_1_oe_o;
	// Trace: design.sv:103755:5
	output wire gpio_27_o;
	// Trace: design.sv:103756:5
	input wire gpio_27_i;
	// Trace: design.sv:103757:5
	output wire gpio_27_oe_o;
	// Trace: design.sv:103759:9
	output wire spi2_sd_2_o;
	// Trace: design.sv:103760:5
	input wire spi2_sd_2_i;
	// Trace: design.sv:103761:5
	output wire spi2_sd_2_oe_o;
	// Trace: design.sv:103762:5
	output wire gpio_28_o;
	// Trace: design.sv:103763:5
	input wire gpio_28_i;
	// Trace: design.sv:103764:5
	output wire gpio_28_oe_o;
	// Trace: design.sv:103766:9
	output wire spi2_sd_3_o;
	// Trace: design.sv:103767:5
	input wire spi2_sd_3_i;
	// Trace: design.sv:103768:5
	output wire spi2_sd_3_oe_o;
	// Trace: design.sv:103769:5
	output wire gpio_29_o;
	// Trace: design.sv:103770:5
	input wire gpio_29_i;
	// Trace: design.sv:103771:5
	output wire gpio_29_oe_o;
	// Trace: design.sv:103773:9
	output wire i2c_scl_o;
	// Trace: design.sv:103774:5
	input wire i2c_scl_i;
	// Trace: design.sv:103775:5
	output wire i2c_scl_oe_o;
	// Trace: design.sv:103776:5
	output wire gpio_31_o;
	// Trace: design.sv:103777:5
	input wire gpio_31_i;
	// Trace: design.sv:103778:5
	output wire gpio_31_oe_o;
	// Trace: design.sv:103780:9
	output wire i2c_sda_o;
	// Trace: design.sv:103781:5
	input wire i2c_sda_i;
	// Trace: design.sv:103782:5
	output wire i2c_sda_oe_o;
	// Trace: design.sv:103783:5
	output wire gpio_30_o;
	// Trace: design.sv:103784:5
	input wire gpio_30_i;
	// Trace: design.sv:103785:5
	output wire gpio_30_oe_o;
	// Trace: design.sv:103796:5
	// removed localparam type reg_pkg_reg_req_t
	output wire [69:0] pad_req_o;
	// Trace: design.sv:103797:5
	// removed localparam type reg_pkg_reg_rsp_t
	input wire [33:0] pad_resp_i;
	// Trace: design.sv:103799:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [(EXT_XBAR_NMASTER * 70) - 1:0] ext_xbar_master_req_i;
	// Trace: design.sv:103800:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [(EXT_XBAR_NMASTER * 34) - 1:0] ext_xbar_master_resp_o;
	// Trace: design.sv:103802:5
	output wire [69:0] ext_xbar_slave_req_o;
	// Trace: design.sv:103803:5
	input wire [33:0] ext_xbar_slave_resp_i;
	// Trace: design.sv:103805:5
	output wire [69:0] ext_peripheral_slave_req_o;
	// Trace: design.sv:103806:5
	input wire [33:0] ext_peripheral_slave_resp_i;
	// Trace: design.sv:103808:5
	localparam core_v_mini_mcu_pkg_PLIC_NINT = 64;
	localparam core_v_mini_mcu_pkg_PLIC_USED_NINT = 50;
	localparam core_v_mini_mcu_pkg_NEXT_INT = 14;
	input wire [13:0] intr_vector_ext_i;
	// Trace: design.sv:103810:5
	output wire cpu_subsystem_powergate_switch_o;
	// Trace: design.sv:103811:5
	input wire cpu_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:103812:5
	output wire peripheral_subsystem_powergate_switch_o;
	// Trace: design.sv:103813:5
	input wire peripheral_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:103814:5
	localparam [31:0] core_v_mini_mcu_pkg_NUM_BANKS = 2;
	output wire [1:0] memory_subsystem_banks_powergate_switch_o;
	// Trace: design.sv:103815:5
	input wire [1:0] memory_subsystem_banks_powergate_switch_ack_i;
	// Trace: design.sv:103816:5
	localparam [31:0] core_v_mini_mcu_pkg_EXTERNAL_DOMAINS = 0;
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_switch_o;
	// Trace: design.sv:103817:5
	input wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:103818:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_iso_o;
	// Trace: design.sv:103819:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_rst_no;
	// Trace: design.sv:103820:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_ram_banks_set_retentive_o;
	// Trace: design.sv:103822:5
	output wire [31:0] exit_value_o;
	// Trace: design.sv:103825:3
	// removed import core_v_mini_mcu_pkg::*;
	// Trace: design.sv:103826:3
	// removed import cv32e40p_apu_core_pkg::*;
	// Trace: design.sv:103828:3
	localparam [31:0] core_v_mini_mcu_pkg_MEM_SIZE = 32'h00010000;
	localparam NUM_BYTES = core_v_mini_mcu_pkg_MEM_SIZE;
	// Trace: design.sv:103829:3
	localparam [31:0] core_v_mini_mcu_pkg_DEBUG_START_ADDRESS = 32'h10000000;
	localparam DM_HALTADDRESS = core_v_mini_mcu_pkg_DEBUG_START_ADDRESS + 32'h00000800;
	// Trace: design.sv:103831:3
	localparam JTAG_IDCODE = 32'h10001c05;
	// Trace: design.sv:103832:3
	localparam [31:0] core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS = 32'h20000000;
	localparam [31:0] core_v_mini_mcu_pkg_BOOTROM_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00010000;
	localparam BOOT_ADDR = core_v_mini_mcu_pkg_BOOTROM_START_ADDRESS;
	// Trace: design.sv:103833:3
	localparam NUM_MHPMCOUNTERS = 1;
	// Trace: design.sv:103843:3
	wire [69:0] core_instr_req;
	// Trace: design.sv:103844:3
	wire [33:0] core_instr_resp;
	// Trace: design.sv:103845:3
	wire [69:0] core_data_req;
	// Trace: design.sv:103846:3
	wire [33:0] core_data_resp;
	// Trace: design.sv:103847:3
	wire [69:0] debug_master_req;
	// Trace: design.sv:103848:3
	wire [33:0] debug_master_resp;
	// Trace: design.sv:103849:3
	wire [69:0] dma_master0_ch0_req;
	// Trace: design.sv:103850:3
	wire [33:0] dma_master0_ch0_resp;
	// Trace: design.sv:103851:3
	wire [69:0] dma_master1_ch0_req;
	// Trace: design.sv:103852:3
	wire [33:0] dma_master1_ch0_resp;
	// Trace: design.sv:103855:3
	wire [139:0] ram_slave_req;
	// Trace: design.sv:103856:3
	wire [67:0] ram_slave_resp;
	// Trace: design.sv:103859:3
	wire [69:0] debug_slave_req;
	// Trace: design.sv:103860:3
	wire [33:0] debug_slave_resp;
	// Trace: design.sv:103863:3
	wire [69:0] ao_peripheral_slave_req;
	// Trace: design.sv:103864:3
	wire [33:0] ao_peripheral_slave_resp;
	// Trace: design.sv:103865:3
	wire [69:0] peripheral_slave_req;
	// Trace: design.sv:103866:3
	wire [33:0] peripheral_slave_resp;
	// Trace: design.sv:103869:3
	wire debug_core_req;
	// Trace: design.sv:103872:3
	wire core_sleep;
	// Trace: design.sv:103875:3
	wire irq_ack;
	// Trace: design.sv:103876:3
	wire [4:0] irq_id_out;
	// Trace: design.sv:103877:3
	wire irq_software;
	// Trace: design.sv:103878:3
	wire irq_external;
	// Trace: design.sv:103879:3
	wire [14:0] irq_fast;
	// Trace: design.sv:103882:3
	wire [69:0] flash_mem_slave_req;
	// Trace: design.sv:103883:3
	wire [33:0] flash_mem_slave_resp;
	// Trace: design.sv:103886:3
	wire [3:0] rv_timer_intr;
	// Trace: design.sv:103889:3
	wire [31:0] intr;
	// Trace: design.sv:103890:3
	wire [14:0] fast_intr;
	// Trace: design.sv:103893:3
	wire cpu_subsystem_powergate_iso;
	// Trace: design.sv:103894:3
	wire cpu_subsystem_rst_n;
	// Trace: design.sv:103895:3
	wire peripheral_subsystem_powergate_iso;
	// Trace: design.sv:103896:3
	wire peripheral_subsystem_rst_n;
	// Trace: design.sv:103897:3
	wire [1:0] memory_subsystem_banks_powergate_iso;
	// Trace: design.sv:103898:3
	wire [1:0] memory_subsystem_banks_set_retentive;
	// Trace: design.sv:103901:4
	wire peripheral_subsystem_clkgate_en;
	// Trace: design.sv:103902:4
	wire [1:0] memory_subsystem_clkgate_en;
	// Trace: design.sv:103905:3
	wire dma_intr;
	// Trace: design.sv:103908:3
	wire spi_flash_intr;
	wire spi_intr;
	// Trace: design.sv:103911:3
	wire [31:8] gpio_in;
	// Trace: design.sv:103912:3
	wire [31:8] gpio_out;
	// Trace: design.sv:103913:3
	wire [31:8] gpio_oe;
	// Trace: design.sv:103916:3
	wire [7:0] gpio_ao_in;
	// Trace: design.sv:103917:3
	wire [7:0] gpio_ao_out;
	// Trace: design.sv:103918:3
	wire [7:0] gpio_ao_oe;
	// Trace: design.sv:103919:3
	wire [7:0] gpio_ao_intr;
	// Trace: design.sv:103922:3
	wire uart_intr_tx_watermark;
	// Trace: design.sv:103923:3
	wire uart_intr_rx_watermark;
	// Trace: design.sv:103924:3
	wire uart_intr_tx_empty;
	// Trace: design.sv:103925:3
	wire uart_intr_rx_overflow;
	// Trace: design.sv:103926:3
	wire uart_intr_rx_frame_err;
	// Trace: design.sv:103927:3
	wire uart_intr_rx_break_err;
	// Trace: design.sv:103928:3
	wire uart_intr_rx_timeout;
	// Trace: design.sv:103929:3
	wire uart_intr_rx_parity_err;
	// Trace: design.sv:103931:3
	assign intr = {1'b0, irq_fast, 4'b0000, irq_external, 3'b000, rv_timer_intr[0], 3'b000, irq_software, 3'b000};
	// Trace: design.sv:103935:3
	assign fast_intr = {1'b0, gpio_ao_intr, spi_flash_intr, spi_intr, dma_intr, rv_timer_intr[3], rv_timer_intr[2], rv_timer_intr[1]};
	// Trace: design.sv:103946:3
	cpu_subsystem #(
		.BOOT_ADDR(BOOT_ADDR),
		.PULP_XPULP(PULP_XPULP),
		.FPU(FPU),
		.PULP_ZFINX(PULP_ZFINX),
		.NUM_MHPMCOUNTERS(NUM_MHPMCOUNTERS),
		.DM_HALTADDRESS(DM_HALTADDRESS),
		.X_EXT(X_EXT)
	) cpu_subsystem_i(
		.clk_i(clk_i),
		.rst_ni(cpu_subsystem_rst_n),
		.core_instr_req_o(core_instr_req),
		.core_instr_resp_i(core_instr_resp),
		.core_data_req_o(core_data_req),
		.core_data_resp_i(core_data_resp),
		.irq_i(intr),
		.irq_ack_o(irq_ack),
		.irq_id_o(irq_id_out),
		.debug_req_i(debug_core_req),
		.core_sleep_o(core_sleep)
	);
	// Trace: design.sv:103977:3
	debug_subsystem #(.JTAG_IDCODE(JTAG_IDCODE)) debug_subsystem_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.jtag_tck_i(jtag_tck_i),
		.jtag_tms_i(jtag_tms_i),
		.jtag_trst_ni(jtag_trst_ni),
		.jtag_tdi_i(jtag_tdi_i),
		.jtag_tdo_o(jtag_tdo_o),
		.debug_core_req_o(debug_core_req),
		.debug_slave_req_i(debug_slave_req),
		.debug_slave_resp_o(debug_slave_resp),
		.debug_master_req_o(debug_master_req),
		.debug_master_resp_i(debug_master_resp)
	);
	// Trace: design.sv:103994:3
	system_bus #(
		.NUM_BANKS(core_v_mini_mcu_pkg_NUM_BANKS),
		.EXT_XBAR_NMASTER(EXT_XBAR_NMASTER)
	) system_bus_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.core_instr_req_i(core_instr_req),
		.core_instr_resp_o(core_instr_resp),
		.core_data_req_i(core_data_req),
		.core_data_resp_o(core_data_resp),
		.debug_master_req_i(debug_master_req),
		.debug_master_resp_o(debug_master_resp),
		.dma_master0_ch0_req_i(dma_master0_ch0_req),
		.dma_master0_ch0_resp_o(dma_master0_ch0_resp),
		.dma_master1_ch0_req_i(dma_master1_ch0_req),
		.dma_master1_ch0_resp_o(dma_master1_ch0_resp),
		.ext_xbar_master_req_i(ext_xbar_master_req_i),
		.ext_xbar_master_resp_o(ext_xbar_master_resp_o),
		.ram_req_o(ram_slave_req),
		.ram_resp_i(ram_slave_resp),
		.debug_slave_req_o(debug_slave_req),
		.debug_slave_resp_i(debug_slave_resp),
		.ao_peripheral_slave_req_o(ao_peripheral_slave_req),
		.ao_peripheral_slave_resp_i(ao_peripheral_slave_resp),
		.peripheral_slave_req_o(peripheral_slave_req),
		.peripheral_slave_resp_i(peripheral_slave_resp),
		.flash_mem_slave_req_o(flash_mem_slave_req),
		.flash_mem_slave_resp_i(flash_mem_slave_resp),
		.ext_xbar_slave_req_o(ext_xbar_slave_req_o),
		.ext_xbar_slave_resp_i(ext_xbar_slave_resp_i)
	);
	// Trace: design.sv:104026:3
	memory_subsystem #(.NUM_BANKS(core_v_mini_mcu_pkg_NUM_BANKS)) memory_subsystem_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clk_gate_en_i(memory_subsystem_clkgate_en),
		.ram_req_i(ram_slave_req),
		.ram_resp_o(ram_slave_resp),
		.set_retentive_i(memory_subsystem_banks_set_retentive)
	);
	// Trace: design.sv:104037:3
	ao_peripheral_subsystem ao_peripheral_subsystem_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.slave_req_i(ao_peripheral_slave_req),
		.slave_resp_o(ao_peripheral_slave_resp),
		.boot_select_i(boot_select_i),
		.execute_from_flash_i(execute_from_flash_i),
		.exit_valid_o(exit_valid_o),
		.exit_value_o(exit_value_o),
		.spimemio_req_i(flash_mem_slave_req),
		.spimemio_resp_o(flash_mem_slave_resp),
		.spi_flash_sck_o(spi_flash_sck_o),
		.spi_flash_sck_en_o(spi_flash_sck_oe_o),
		.spi_flash_csb_o({spi_flash_cs_1_o, spi_flash_cs_0_o}),
		.spi_flash_csb_en_o({spi_flash_cs_1_oe_o, spi_flash_cs_0_oe_o}),
		.spi_flash_sd_o({spi_flash_sd_3_o, spi_flash_sd_2_o, spi_flash_sd_1_o, spi_flash_sd_0_o}),
		.spi_flash_sd_en_o({spi_flash_sd_3_oe_o, spi_flash_sd_2_oe_o, spi_flash_sd_1_oe_o, spi_flash_sd_0_oe_o}),
		.spi_flash_sd_i({spi_flash_sd_3_i, spi_flash_sd_2_i, spi_flash_sd_1_i, spi_flash_sd_0_i}),
		.spi_sck_o(spi_sck_o),
		.spi_sck_en_o(spi_sck_oe_o),
		.spi_csb_o({spi_cs_1_o, spi_cs_0_o}),
		.spi_csb_en_o({spi_cs_1_oe_o, spi_cs_0_oe_o}),
		.spi_sd_o({spi_sd_3_o, spi_sd_2_o, spi_sd_1_o, spi_sd_0_o}),
		.spi_sd_en_o({spi_sd_3_oe_o, spi_sd_2_oe_o, spi_sd_1_oe_o, spi_sd_0_oe_o}),
		.spi_sd_i({spi_sd_3_i, spi_sd_2_i, spi_sd_1_i, spi_sd_0_i}),
		.intr_i(intr),
		.intr_vector_ext_i(intr_vector_ext_i),
		.core_sleep_i(core_sleep),
		.cpu_subsystem_powergate_switch_o(cpu_subsystem_powergate_switch_o),
		.cpu_subsystem_powergate_switch_ack_i(cpu_subsystem_powergate_switch_ack_i),
		.cpu_subsystem_powergate_iso_o(cpu_subsystem_powergate_iso),
		.cpu_subsystem_rst_no(cpu_subsystem_rst_n),
		.peripheral_subsystem_powergate_switch_o(peripheral_subsystem_powergate_switch_o),
		.peripheral_subsystem_powergate_switch_ack_i(peripheral_subsystem_powergate_switch_ack_i),
		.peripheral_subsystem_powergate_iso_o(peripheral_subsystem_powergate_iso),
		.peripheral_subsystem_rst_no(peripheral_subsystem_rst_n),
		.memory_subsystem_banks_powergate_switch_o(memory_subsystem_banks_powergate_switch_o),
		.memory_subsystem_banks_powergate_switch_ack_i(memory_subsystem_banks_powergate_switch_ack_i),
		.memory_subsystem_banks_powergate_iso_o(memory_subsystem_banks_powergate_iso),
		.memory_subsystem_banks_set_retentive_o(memory_subsystem_banks_set_retentive),
		.external_subsystem_powergate_switch_o(external_subsystem_powergate_switch_o),
		.external_subsystem_powergate_switch_ack_i(external_subsystem_powergate_switch_ack_i),
		.external_subsystem_powergate_iso_o(external_subsystem_powergate_iso_o),
		.external_subsystem_rst_no(external_subsystem_rst_no),
		.external_ram_banks_set_retentive_o(external_ram_banks_set_retentive_o),
		.peripheral_subsystem_clkgate_en_o(peripheral_subsystem_clkgate_en),
		.memory_subsystem_clkgate_en_o(memory_subsystem_clkgate_en),
		.rv_timer_0_intr_o(rv_timer_intr[0]),
		.rv_timer_1_intr_o(rv_timer_intr[1]),
		.dma_master0_ch0_req_o(dma_master0_ch0_req),
		.dma_master0_ch0_resp_i(dma_master0_ch0_resp),
		.dma_master1_ch0_req_o(dma_master1_ch0_req),
		.dma_master1_ch0_resp_i(dma_master1_ch0_resp),
		.dma_intr_o(dma_intr),
		.spi_intr_event_o(spi_intr),
		.spi_flash_intr_event_o(spi_flash_intr),
		.pad_req_o(pad_req_o),
		.pad_resp_i(pad_resp_i),
		.fast_intr_i(fast_intr),
		.fast_intr_o(irq_fast),
		.cio_gpio_i(gpio_ao_in),
		.cio_gpio_o(gpio_ao_out),
		.cio_gpio_en_o(gpio_ao_oe),
		.intr_gpio_o(gpio_ao_intr),
		.uart_rx_i(uart_rx_i),
		.uart_tx_o(uart_tx_o),
		.uart_intr_tx_watermark_o(uart_intr_tx_watermark),
		.uart_intr_rx_watermark_o(uart_intr_rx_watermark),
		.uart_intr_tx_empty_o(uart_intr_tx_empty),
		.uart_intr_rx_overflow_o(uart_intr_rx_overflow),
		.uart_intr_rx_frame_err_o(uart_intr_rx_frame_err),
		.uart_intr_rx_break_err_o(uart_intr_rx_break_err),
		.uart_intr_rx_timeout_o(uart_intr_rx_timeout),
		.uart_intr_rx_parity_err_o(uart_intr_rx_parity_err),
		.ext_peripheral_slave_req_o(ext_peripheral_slave_req_o),
		.ext_peripheral_slave_resp_i(ext_peripheral_slave_resp_i)
	);
	// Trace: design.sv:104115:3
	peripheral_subsystem #(.NEXT_INT(core_v_mini_mcu_pkg_NEXT_INT)) peripheral_subsystem_i(
		.clk_i(clk_i),
		.rst_ni(peripheral_subsystem_rst_n),
		.clk_gate_en_i(peripheral_subsystem_clkgate_en),
		.slave_req_i(peripheral_slave_req),
		.slave_resp_o(peripheral_slave_resp),
		.intr_vector_ext_i(intr_vector_ext_i),
		.irq_plic_o(irq_external),
		.msip_o(irq_software),
		.uart_intr_tx_watermark_i(uart_intr_tx_watermark),
		.uart_intr_rx_watermark_i(uart_intr_rx_watermark),
		.uart_intr_tx_empty_i(uart_intr_tx_empty),
		.uart_intr_rx_overflow_i(uart_intr_rx_overflow),
		.uart_intr_rx_frame_err_i(uart_intr_rx_frame_err),
		.uart_intr_rx_break_err_i(uart_intr_rx_break_err),
		.uart_intr_rx_timeout_i(uart_intr_rx_timeout),
		.uart_intr_rx_parity_err_i(uart_intr_rx_parity_err),
		.cio_gpio_i(gpio_in),
		.cio_gpio_o(gpio_out),
		.cio_gpio_en_o(gpio_oe),
		.cio_scl_i(i2c_scl_i),
		.cio_scl_o(i2c_scl_o),
		.cio_scl_en_o(i2c_scl_oe_o),
		.cio_sda_i(i2c_sda_i),
		.cio_sda_o(i2c_sda_o),
		.cio_sda_en_o(i2c_sda_oe_o),
		.spi2_sck_o(spi2_sck_o),
		.spi2_sck_en_o(spi2_sck_oe_o),
		.spi2_csb_o({spi2_cs_1_o, spi2_cs_0_o}),
		.spi2_csb_en_o({spi2_cs_1_oe_o, spi2_cs_0_oe_o}),
		.spi2_sd_o({spi2_sd_3_o, spi2_sd_2_o, spi2_sd_1_o, spi2_sd_0_o}),
		.spi2_sd_en_o({spi2_sd_3_oe_o, spi2_sd_2_oe_o, spi2_sd_1_oe_o, spi2_sd_0_oe_o}),
		.spi2_sd_i({spi2_sd_3_i, spi2_sd_2_i, spi2_sd_1_i, spi2_sd_0_i}),
		.rv_timer_2_intr_o(rv_timer_intr[2]),
		.rv_timer_3_intr_o(rv_timer_intr[3])
	);
	// Trace: design.sv:104154:3
	assign gpio_ao_in[0] = gpio_0_i;
	// Trace: design.sv:104155:3
	assign gpio_0_o = gpio_ao_out[0];
	// Trace: design.sv:104156:3
	assign gpio_0_oe_o = gpio_ao_oe[0];
	// Trace: design.sv:104157:3
	assign gpio_ao_in[1] = gpio_1_i;
	// Trace: design.sv:104158:3
	assign gpio_1_o = gpio_ao_out[1];
	// Trace: design.sv:104159:3
	assign gpio_1_oe_o = gpio_ao_oe[1];
	// Trace: design.sv:104160:3
	assign gpio_ao_in[2] = gpio_2_i;
	// Trace: design.sv:104161:3
	assign gpio_2_o = gpio_ao_out[2];
	// Trace: design.sv:104162:3
	assign gpio_2_oe_o = gpio_ao_oe[2];
	// Trace: design.sv:104163:3
	assign gpio_ao_in[3] = gpio_3_i;
	// Trace: design.sv:104164:3
	assign gpio_3_o = gpio_ao_out[3];
	// Trace: design.sv:104165:3
	assign gpio_3_oe_o = gpio_ao_oe[3];
	// Trace: design.sv:104166:3
	assign gpio_ao_in[4] = gpio_4_i;
	// Trace: design.sv:104167:3
	assign gpio_4_o = gpio_ao_out[4];
	// Trace: design.sv:104168:3
	assign gpio_4_oe_o = gpio_ao_oe[4];
	// Trace: design.sv:104169:3
	assign gpio_ao_in[5] = gpio_5_i;
	// Trace: design.sv:104170:3
	assign gpio_5_o = gpio_ao_out[5];
	// Trace: design.sv:104171:3
	assign gpio_5_oe_o = gpio_ao_oe[5];
	// Trace: design.sv:104172:3
	assign gpio_ao_in[6] = gpio_6_i;
	// Trace: design.sv:104173:3
	assign gpio_6_o = gpio_ao_out[6];
	// Trace: design.sv:104174:3
	assign gpio_6_oe_o = gpio_ao_oe[6];
	// Trace: design.sv:104175:3
	assign gpio_ao_in[7] = gpio_7_i;
	// Trace: design.sv:104176:3
	assign gpio_7_o = gpio_ao_out[7];
	// Trace: design.sv:104177:3
	assign gpio_7_oe_o = gpio_ao_oe[7];
	// Trace: design.sv:104178:3
	assign gpio_in[8] = gpio_8_i;
	// Trace: design.sv:104179:3
	assign gpio_8_o = gpio_out[8];
	// Trace: design.sv:104180:3
	assign gpio_8_oe_o = gpio_oe[8];
	// Trace: design.sv:104181:3
	assign gpio_in[9] = gpio_9_i;
	// Trace: design.sv:104182:3
	assign gpio_9_o = gpio_out[9];
	// Trace: design.sv:104183:3
	assign gpio_9_oe_o = gpio_oe[9];
	// Trace: design.sv:104184:3
	assign gpio_in[10] = gpio_10_i;
	// Trace: design.sv:104185:3
	assign gpio_10_o = gpio_out[10];
	// Trace: design.sv:104186:3
	assign gpio_10_oe_o = gpio_oe[10];
	// Trace: design.sv:104187:3
	assign gpio_in[11] = gpio_11_i;
	// Trace: design.sv:104188:3
	assign gpio_11_o = gpio_out[11];
	// Trace: design.sv:104189:3
	assign gpio_11_oe_o = gpio_oe[11];
	// Trace: design.sv:104190:3
	assign gpio_in[12] = gpio_12_i;
	// Trace: design.sv:104191:3
	assign gpio_12_o = gpio_out[12];
	// Trace: design.sv:104192:3
	assign gpio_12_oe_o = gpio_oe[12];
	// Trace: design.sv:104193:3
	assign gpio_in[13] = gpio_13_i;
	// Trace: design.sv:104194:3
	assign gpio_13_o = gpio_out[13];
	// Trace: design.sv:104195:3
	assign gpio_13_oe_o = gpio_oe[13];
	// Trace: design.sv:104196:3
	assign gpio_in[14] = gpio_14_i;
	// Trace: design.sv:104197:3
	assign gpio_14_o = gpio_out[14];
	// Trace: design.sv:104198:3
	assign gpio_14_oe_o = gpio_oe[14];
	// Trace: design.sv:104199:3
	assign gpio_in[15] = gpio_15_i;
	// Trace: design.sv:104200:3
	assign gpio_15_o = gpio_out[15];
	// Trace: design.sv:104201:3
	assign gpio_15_oe_o = gpio_oe[15];
	// Trace: design.sv:104202:3
	assign gpio_in[16] = gpio_16_i;
	// Trace: design.sv:104203:3
	assign gpio_16_o = gpio_out[16];
	// Trace: design.sv:104204:3
	assign gpio_16_oe_o = gpio_oe[16];
	// Trace: design.sv:104205:3
	assign gpio_in[17] = gpio_17_i;
	// Trace: design.sv:104206:3
	assign gpio_17_o = gpio_out[17];
	// Trace: design.sv:104207:3
	assign gpio_17_oe_o = gpio_oe[17];
	// Trace: design.sv:104208:3
	assign gpio_in[18] = gpio_18_i;
	// Trace: design.sv:104209:3
	assign gpio_18_o = gpio_out[18];
	// Trace: design.sv:104210:3
	assign gpio_18_oe_o = gpio_oe[18];
	// Trace: design.sv:104211:3
	assign gpio_in[19] = gpio_19_i;
	// Trace: design.sv:104212:3
	assign gpio_19_o = gpio_out[19];
	// Trace: design.sv:104213:3
	assign gpio_19_oe_o = gpio_oe[19];
	// Trace: design.sv:104214:3
	assign gpio_in[20] = gpio_20_i;
	// Trace: design.sv:104215:3
	assign gpio_20_o = gpio_out[20];
	// Trace: design.sv:104216:3
	assign gpio_20_oe_o = gpio_oe[20];
	// Trace: design.sv:104217:3
	assign gpio_in[21] = gpio_21_i;
	// Trace: design.sv:104218:3
	assign gpio_21_o = gpio_out[21];
	// Trace: design.sv:104219:3
	assign gpio_21_oe_o = gpio_oe[21];
	// Trace: design.sv:104220:3
	assign gpio_in[22] = gpio_22_i;
	// Trace: design.sv:104221:3
	assign gpio_22_o = gpio_out[22];
	// Trace: design.sv:104222:3
	assign gpio_22_oe_o = gpio_oe[22];
	// Trace: design.sv:104223:3
	assign gpio_in[23] = gpio_23_i;
	// Trace: design.sv:104224:3
	assign gpio_23_o = gpio_out[23];
	// Trace: design.sv:104225:3
	assign gpio_23_oe_o = gpio_oe[23];
	// Trace: design.sv:104226:3
	assign gpio_in[24] = gpio_24_i;
	// Trace: design.sv:104227:3
	assign gpio_24_o = gpio_out[24];
	// Trace: design.sv:104228:3
	assign gpio_24_oe_o = gpio_oe[24];
	// Trace: design.sv:104229:3
	assign gpio_in[25] = gpio_25_i;
	// Trace: design.sv:104230:3
	assign gpio_25_o = gpio_out[25];
	// Trace: design.sv:104231:3
	assign gpio_25_oe_o = gpio_oe[25];
	// Trace: design.sv:104232:3
	assign gpio_in[26] = gpio_26_i;
	// Trace: design.sv:104233:3
	assign gpio_26_o = gpio_out[26];
	// Trace: design.sv:104234:3
	assign gpio_26_oe_o = gpio_oe[26];
	// Trace: design.sv:104235:3
	assign gpio_in[27] = gpio_27_i;
	// Trace: design.sv:104236:3
	assign gpio_27_o = gpio_out[27];
	// Trace: design.sv:104237:3
	assign gpio_27_oe_o = gpio_oe[27];
	// Trace: design.sv:104238:3
	assign gpio_in[28] = gpio_28_i;
	// Trace: design.sv:104239:3
	assign gpio_28_o = gpio_out[28];
	// Trace: design.sv:104240:3
	assign gpio_28_oe_o = gpio_oe[28];
	// Trace: design.sv:104241:3
	assign gpio_in[29] = gpio_29_i;
	// Trace: design.sv:104242:3
	assign gpio_29_o = gpio_out[29];
	// Trace: design.sv:104243:3
	assign gpio_29_oe_o = gpio_oe[29];
	// Trace: design.sv:104244:3
	assign gpio_in[30] = gpio_30_i;
	// Trace: design.sv:104245:3
	assign gpio_30_o = gpio_out[30];
	// Trace: design.sv:104246:3
	assign gpio_30_oe_o = gpio_oe[30];
	// Trace: design.sv:104247:3
	assign gpio_in[31] = gpio_31_i;
	// Trace: design.sv:104248:3
	assign gpio_31_o = gpio_out[31];
	// Trace: design.sv:104249:3
	assign gpio_31_oe_o = gpio_oe[31];
endmodule
module cpu_subsystem (
	clk_i,
	rst_ni,
	core_instr_req_o,
	core_instr_resp_i,
	core_data_req_o,
	core_data_resp_i,
	irq_i,
	irq_ack_o,
	irq_id_o,
	debug_req_i,
	core_sleep_o
);
	// removed import obi_pkg::*;
	// removed import core_v_mini_mcu_pkg::*;
	// Trace: design.sv:104260:15
	parameter BOOT_ADDR = 'h180;
	// Trace: design.sv:104261:15
	parameter PULP_XPULP = 0;
	// Trace: design.sv:104262:15
	parameter FPU = 0;
	// Trace: design.sv:104263:15
	parameter PULP_ZFINX = 0;
	// Trace: design.sv:104264:15
	parameter NUM_MHPMCOUNTERS = 1;
	// Trace: design.sv:104265:15
	parameter DM_HALTADDRESS = 1'sb0;
	// Trace: design.sv:104266:15
	parameter X_EXT = 0;
	// Trace: design.sv:104267:15
	// removed localparam type core_v_mini_mcu_pkg_cpu_type_e
	localparam [1:0] core_v_mini_mcu_pkg_CpuType = 2'd1;
	parameter [1:0] CPU_TYPE = core_v_mini_mcu_pkg_CpuType;
	// Trace: design.sv:104270:5
	input wire clk_i;
	// Trace: design.sv:104271:5
	input wire rst_ni;
	// Trace: design.sv:104274:5
	// removed localparam type obi_pkg_obi_req_t
	output wire [69:0] core_instr_req_o;
	// Trace: design.sv:104275:5
	// removed localparam type obi_pkg_obi_resp_t
	input wire [33:0] core_instr_resp_i;
	// Trace: design.sv:104278:5
	output wire [69:0] core_data_req_o;
	// Trace: design.sv:104279:5
	input wire [33:0] core_data_resp_i;
	// Trace: design.sv:104291:5
	input wire [31:0] irq_i;
	// Trace: design.sv:104292:5
	output wire irq_ack_o;
	// Trace: design.sv:104293:5
	output wire [4:0] irq_id_o;
	// Trace: design.sv:104296:5
	input wire debug_req_i;
	// Trace: design.sv:104299:5
	output wire core_sleep_o;
	// Trace: design.sv:104304:3
	wire fetch_enable;
	// Trace: design.sv:104306:3
	assign fetch_enable = 1'b1;
	// Trace: design.sv:104308:3
	assign core_instr_req_o[31-:32] = 1'sb0;
	// Trace: design.sv:104309:3
	assign core_instr_req_o[68] = 1'sb0;
	// Trace: design.sv:104310:3
	assign core_instr_req_o[67-:4] = 4'b1111;
	// Trace: design.sv:104312:3
	generate
		if (CPU_TYPE == 2'd1) begin : gen_cv32e20
			// Trace: design.sv:104314:5
			wire [4:0] rf_raddr_a;
			wire [4:0] rf_raddr_b;
			wire [4:0] rf_waddr_wb;
			// Trace: design.sv:104315:5
			wire [31:0] rf_rdata_a;
			wire [31:0] rf_rdata_b;
			wire [31:0] rf_wdata_wb;
			// Trace: design.sv:104316:5
			wire rf_we_wb;
			// Trace: design.sv:104318:5
			// removed import ibex_pkg::*;
			// Trace: design.sv:104320:5
			ibex_core #(
				.DmHaltAddr(DM_HALTADDRESS),
				.DmExceptionAddr(32'h00000000),
				.DbgTriggerEn(1'b1),
				.ResetAll(1'b1)
			) cv32e20_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.hart_id_i(32'h00000000),
				.boot_addr_i(BOOT_ADDR),
				.instr_addr_o(core_instr_req_o[63-:32]),
				.instr_req_o(core_instr_req_o[69]),
				.instr_rdata_i(core_instr_resp_i[31-:32]),
				.instr_gnt_i(core_instr_resp_i[33]),
				.instr_rvalid_i(core_instr_resp_i[32]),
				.instr_err_i(1'b0),
				.data_addr_o(core_data_req_o[63-:32]),
				.data_wdata_o(core_data_req_o[31-:32]),
				.data_we_o(core_data_req_o[68]),
				.data_req_o(core_data_req_o[69]),
				.data_be_o(core_data_req_o[67-:4]),
				.data_rdata_i(core_data_resp_i[31-:32]),
				.data_gnt_i(core_data_resp_i[33]),
				.data_rvalid_i(core_data_resp_i[32]),
				.data_err_i(1'b0),
				.dummy_instr_id_o(),
				.rf_raddr_a_o(rf_raddr_a),
				.rf_raddr_b_o(rf_raddr_b),
				.rf_waddr_wb_o(rf_waddr_wb),
				.rf_we_wb_o(rf_we_wb),
				.rf_wdata_wb_ecc_o(rf_wdata_wb),
				.rf_rdata_a_ecc_i(rf_rdata_a),
				.rf_rdata_b_ecc_i(rf_rdata_b),
				.ic_tag_req_o(),
				.ic_tag_write_o(),
				.ic_tag_addr_o(),
				.ic_tag_wdata_o(),
				.ic_tag_rdata_i(),
				.ic_data_req_o(),
				.ic_data_write_o(),
				.ic_data_addr_o(),
				.ic_data_wdata_o(),
				.ic_data_rdata_i(),
				.ic_scr_key_valid_i(),
				.irq_software_i(irq_i[3]),
				.irq_timer_i(irq_i[7]),
				.irq_external_i(irq_i[11]),
				.irq_fast_i(irq_i[30:16]),
				.irq_nm_i(irq_i[31]),
				.irq_pending_o(),
				.debug_req_i(debug_req_i),
				.crash_dump_o(),
				.double_fault_seen_o(),
				.fetch_enable_i(fetch_enable),
				.alert_minor_o(),
				.alert_major_o(),
				.icache_inval_o(),
				.core_sleep_o(core_sleep_o)
			);
			// Trace: design.sv:104388:5
			localparam sv2v_uu_cv32e20_register_file_i_ADDR_WIDTH = 6;
			// removed localparam type sv2v_uu_cv32e20_register_file_i_raddr_c_i
			localparam [5:0] sv2v_uu_cv32e20_register_file_i_ext_raddr_c_i_0 = 1'sb0;
			// removed localparam type sv2v_uu_cv32e20_register_file_i_waddr_b_i
			localparam [5:0] sv2v_uu_cv32e20_register_file_i_ext_waddr_b_i_0 = 1'sb0;
			localparam sv2v_uu_cv32e20_register_file_i_DATA_WIDTH = 32;
			// removed localparam type sv2v_uu_cv32e20_register_file_i_wdata_b_i
			localparam [31:0] sv2v_uu_cv32e20_register_file_i_ext_wdata_b_i_0 = 1'sb0;
			// removed localparam type sv2v_uu_cv32e20_register_file_i_we_b_i
			localparam [0:0] sv2v_uu_cv32e20_register_file_i_ext_we_b_i_0 = 1'sb0;
			cv32e40p_register_file #(.ADDR_WIDTH(6)) cv32e20_register_file_i(
				.clk(clk_i),
				.rst_n(rst_ni),
				.scan_cg_en_i(1'b0),
				.raddr_a_i({1'b0, rf_raddr_a}),
				.rdata_a_o(rf_rdata_a),
				.raddr_b_i({1'b0, rf_raddr_b}),
				.rdata_b_o(rf_rdata_b),
				.raddr_c_i(sv2v_uu_cv32e20_register_file_i_ext_raddr_c_i_0),
				.rdata_c_o(),
				.waddr_a_i({1'b0, rf_waddr_wb}),
				.wdata_a_i(rf_wdata_wb),
				.we_a_i(rf_we_wb),
				.waddr_b_i(sv2v_uu_cv32e20_register_file_i_ext_waddr_b_i_0),
				.wdata_b_i(sv2v_uu_cv32e20_register_file_i_ext_wdata_b_i_0),
				.we_b_i(sv2v_uu_cv32e20_register_file_i_ext_we_b_i_0)
			);
			// Trace: design.sv:104422:5
			assign irq_ack_o = 1'sb0;
			// Trace: design.sv:104423:5
			assign irq_id_o = 1'sb0;
		end
		else if (CPU_TYPE == 2'd2) begin : gen_cv32e40x
			// Trace: design.sv:104428:5
			wire xif_compressed_if;
			wire xif_issue_if;
			wire xif_commit_if;
			wire xif_mem_if;
			wire xif_mem_result_if;
			wire xif_result_if;
			cv32e40x_core #(
				.NUM_MHPMCOUNTERS(NUM_MHPMCOUNTERS),
				.X_EXT(X_EXT)
			) cv32e40x_core_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.scan_cg_en_i(1'b0),
				.boot_addr_i(BOOT_ADDR),
				.dm_exception_addr_i(32'h00000000),
				.dm_halt_addr_i(DM_HALTADDRESS),
				.mhartid_i(32'h00000000),
				.mimpid_patch_i(4'h0),
				.mtvec_addr_i(32'h00000000),
				.instr_req_o(core_instr_req_o[69]),
				.instr_gnt_i(core_instr_resp_i[33]),
				.instr_rvalid_i(core_instr_resp_i[32]),
				.instr_addr_o(core_instr_req_o[63-:32]),
				.instr_memtype_o(),
				.instr_prot_o(),
				.instr_dbg_o(),
				.instr_rdata_i(core_instr_resp_i[31-:32]),
				.instr_err_i(1'b0),
				.data_req_o(core_data_req_o[69]),
				.data_gnt_i(core_data_resp_i[33]),
				.data_rvalid_i(core_data_resp_i[32]),
				.data_addr_o(core_data_req_o[63-:32]),
				.data_be_o(core_data_req_o[67-:4]),
				.data_we_o(core_data_req_o[68]),
				.data_wdata_o(core_data_req_o[31-:32]),
				.data_memtype_o(),
				.data_prot_o(),
				.data_dbg_o(),
				.data_atop_o(),
				.data_rdata_i(core_data_resp_i[31-:32]),
				.data_err_i(1'b0),
				.data_exokay_i(1'b1),
				.mcycle_o(),
				.xif_compressed_if(xif_compressed_if),
				.xif_issue_if(xif_issue_if),
				.xif_commit_if(xif_commit_if),
				.xif_mem_if(xif_mem_if),
				.xif_mem_result_if(xif_mem_result_if),
				.xif_result_if(xif_result_if),
				.irq_i(irq_i),
				.wu_wfe_i(1'b0),
				.clic_irq_i(),
				.clic_irq_id_i(),
				.clic_irq_level_i(),
				.clic_irq_priv_i(),
				.clic_irq_shv_i(),
				.fencei_flush_req_o(),
				.fencei_flush_ack_i(1'b0),
				.debug_req_i(debug_req_i),
				.debug_havereset_o(),
				.debug_running_o(),
				.debug_halted_o(),
				.fetch_enable_i(fetch_enable),
				.core_sleep_o(core_sleep_o)
			);
			// Trace: design.sv:104511:5
			assign irq_ack_o = 1'sb0;
			// Trace: design.sv:104512:5
			assign irq_id_o = 1'sb0;
		end
		else begin : gen_cv32e40p
			// Trace: design.sv:104517:5
			cv32e40p_tb_wrapper #(
				.PULP_XPULP(PULP_XPULP),
				.PULP_CLUSTER(0),
				.FPU(FPU),
				.PULP_ZFINX(PULP_ZFINX),
				.NUM_MHPMCOUNTERS(NUM_MHPMCOUNTERS)
			) cv32e40p_tb_wrapper_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.pulp_clock_en_i(1'b1),
				.scan_cg_en_i(1'b0),
				.boot_addr_i(BOOT_ADDR),
				.mtvec_addr_i(32'h00000000),
				.dm_halt_addr_i(DM_HALTADDRESS),
				.hart_id_i(32'h00000000),
				.dm_exception_addr_i(32'h00000000),
				.instr_addr_o(core_instr_req_o[63-:32]),
				.instr_req_o(core_instr_req_o[69]),
				.instr_rdata_i(core_instr_resp_i[31-:32]),
				.instr_gnt_i(core_instr_resp_i[33]),
				.instr_rvalid_i(core_instr_resp_i[32]),
				.data_addr_o(core_data_req_o[63-:32]),
				.data_wdata_o(core_data_req_o[31-:32]),
				.data_we_o(core_data_req_o[68]),
				.data_req_o(core_data_req_o[69]),
				.data_be_o(core_data_req_o[67-:4]),
				.data_rdata_i(core_data_resp_i[31-:32]),
				.data_gnt_i(core_data_resp_i[33]),
				.data_rvalid_i(core_data_resp_i[32]),
				.irq_i(irq_i),
				.irq_ack_o(irq_ack_o),
				.irq_id_o(irq_id_o),
				.debug_req_i(debug_req_i),
				.debug_havereset_o(),
				.debug_running_o(),
				.debug_halted_o(),
				.fetch_enable_i(fetch_enable),
				.core_sleep_o(core_sleep_o)
			);
		end
	endgenerate
endmodule
module memory_subsystem (
	clk_i,
	rst_ni,
	clk_gate_en_i,
	ram_req_i,
	ram_resp_o,
	set_retentive_i
);
	// removed import obi_pkg::*;
	// Trace: design.sv:104577:15
	parameter NUM_BANKS = 2;
	// Trace: design.sv:104579:5
	input wire clk_i;
	// Trace: design.sv:104580:5
	input wire rst_ni;
	// Trace: design.sv:104583:5
	input wire [NUM_BANKS - 1:0] clk_gate_en_i;
	// Trace: design.sv:104585:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [(NUM_BANKS * 70) - 1:0] ram_req_i;
	// Trace: design.sv:104586:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [(NUM_BANKS * 34) - 1:0] ram_resp_o;
	// Trace: design.sv:104588:5
	localparam [31:0] core_v_mini_mcu_pkg_NUM_BANKS = 2;
	input wire [1:0] set_retentive_i;
	// Trace: design.sv:104591:3
	localparam signed [31:0] NumWords = 8192;
	// Trace: design.sv:104592:3
	localparam signed [31:0] AddrWidth = 15;
	// Trace: design.sv:104594:3
	reg [NUM_BANKS - 1:0] ram_valid_q;
	// Trace: design.sv:104596:3
	wire [NUM_BANKS - 1:0] clk_cg;
	// Trace: design.sv:104597:3
	genvar _gv_i_93;
	generate
		for (_gv_i_93 = 0; _gv_i_93 < NUM_BANKS; _gv_i_93 = _gv_i_93 + 1) begin : gen_sram
			localparam i = _gv_i_93;
			// Trace: design.sv:104599:5
			tc_clk_gating clk_gating_cell_i(
				.clk_i(clk_i),
				.en_i(~clk_gate_en_i[i]),
				.test_en_i(1'b0),
				.clk_o(clk_cg[i])
			);
			// Trace: design.sv:104606:5
			always @(posedge clk_cg[i] or negedge rst_ni)
				// Trace: design.sv:104607:7
				if (!rst_ni)
					// Trace: design.sv:104608:9
					ram_valid_q[i] <= 1'sb0;
				else
					// Trace: design.sv:104610:9
					ram_valid_q[i] <= ram_resp_o[(i * 34) + 33];
			// Trace: design.sv:104614:5
			assign ram_resp_o[(i * 34) + 33] = ram_req_i[(i * 70) + 69];
			// Trace: design.sv:104615:5
			assign ram_resp_o[(i * 34) + 32] = ram_valid_q[i];
			// Trace: design.sv:104618:5
			sram_wrapper #(
				.NumWords(NumWords),
				.DataWidth(32'd32)
			) ram_i(
				.clk_i(clk_cg[i]),
				.rst_ni(rst_ni),
				.req_i(ram_req_i[(i * 70) + 69]),
				.we_i(ram_req_i[(i * 70) + 68]),
				.addr_i(ram_req_i[(i * 70) + 46-:13]),
				.wdata_i(ram_req_i[(i * 70) + 31-:32]),
				.be_i(ram_req_i[(i * 70) + 67-:4]),
				.set_retentive_i(set_retentive_i[i]),
				.rdata_o(ram_resp_o[(i * 34) + 31-:32])
			);
		end
	endgenerate
endmodule
module system_bus (
	clk_i,
	rst_ni,
	core_instr_req_i,
	core_instr_resp_o,
	core_data_req_i,
	core_data_resp_o,
	debug_master_req_i,
	debug_master_resp_o,
	dma_master0_ch0_req_i,
	dma_master0_ch0_resp_o,
	dma_master1_ch0_req_i,
	dma_master1_ch0_resp_o,
	ext_xbar_master_req_i,
	ext_xbar_master_resp_o,
	ram_req_o,
	ram_resp_i,
	debug_slave_req_o,
	debug_slave_resp_i,
	ao_peripheral_slave_req_o,
	ao_peripheral_slave_resp_i,
	peripheral_slave_req_o,
	peripheral_slave_resp_i,
	flash_mem_slave_req_o,
	flash_mem_slave_resp_i,
	ext_xbar_slave_req_o,
	ext_xbar_slave_resp_i
);
	// removed import obi_pkg::*;
	// removed import addr_map_rule_pkg::*;
	// Trace: design.sv:104656:15
	parameter NUM_BANKS = 2;
	// Trace: design.sv:104657:15
	parameter EXT_XBAR_NMASTER = 0;
	// Trace: design.sv:104659:5
	input wire clk_i;
	// Trace: design.sv:104660:5
	input wire rst_ni;
	// Trace: design.sv:104663:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [69:0] core_instr_req_i;
	// Trace: design.sv:104664:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [33:0] core_instr_resp_o;
	// Trace: design.sv:104666:5
	input wire [69:0] core_data_req_i;
	// Trace: design.sv:104667:5
	output wire [33:0] core_data_resp_o;
	// Trace: design.sv:104669:5
	input wire [69:0] debug_master_req_i;
	// Trace: design.sv:104670:5
	output wire [33:0] debug_master_resp_o;
	// Trace: design.sv:104672:5
	input wire [69:0] dma_master0_ch0_req_i;
	// Trace: design.sv:104673:5
	output wire [33:0] dma_master0_ch0_resp_o;
	// Trace: design.sv:104675:5
	input wire [69:0] dma_master1_ch0_req_i;
	// Trace: design.sv:104676:5
	output wire [33:0] dma_master1_ch0_resp_o;
	// Trace: design.sv:104678:5
	input wire [(EXT_XBAR_NMASTER * 70) - 1:0] ext_xbar_master_req_i;
	// Trace: design.sv:104679:5
	output wire [(EXT_XBAR_NMASTER * 34) - 1:0] ext_xbar_master_resp_o;
	// Trace: design.sv:104682:5
	output wire [(NUM_BANKS * 70) - 1:0] ram_req_o;
	// Trace: design.sv:104683:5
	input wire [(NUM_BANKS * 34) - 1:0] ram_resp_i;
	// Trace: design.sv:104685:5
	output wire [69:0] debug_slave_req_o;
	// Trace: design.sv:104686:5
	input wire [33:0] debug_slave_resp_i;
	// Trace: design.sv:104688:5
	output wire [69:0] ao_peripheral_slave_req_o;
	// Trace: design.sv:104689:5
	input wire [33:0] ao_peripheral_slave_resp_i;
	// Trace: design.sv:104691:5
	output wire [69:0] peripheral_slave_req_o;
	// Trace: design.sv:104692:5
	input wire [33:0] peripheral_slave_resp_i;
	// Trace: design.sv:104694:5
	output wire [69:0] flash_mem_slave_req_o;
	// Trace: design.sv:104695:5
	input wire [33:0] flash_mem_slave_resp_i;
	// Trace: design.sv:104697:5
	output wire [69:0] ext_xbar_slave_req_o;
	// Trace: design.sv:104698:5
	input wire [33:0] ext_xbar_slave_resp_i;
	// Trace: design.sv:104701:3
	// removed import core_v_mini_mcu_pkg::*;
	// Trace: design.sv:104703:3
	localparam core_v_mini_mcu_pkg_SYSTEM_XBAR_NMASTER = 5;
	wire [((core_v_mini_mcu_pkg_SYSTEM_XBAR_NMASTER + EXT_XBAR_NMASTER) * 70) - 1:0] master_req;
	// Trace: design.sv:104704:3
	wire [((core_v_mini_mcu_pkg_SYSTEM_XBAR_NMASTER + EXT_XBAR_NMASTER) * 34) - 1:0] master_resp;
	// Trace: design.sv:104705:3
	localparam core_v_mini_mcu_pkg_SYSTEM_XBAR_NSLAVE = 8;
	wire [559:0] slave_req;
	// Trace: design.sv:104706:3
	wire [271:0] slave_resp;
	// Trace: design.sv:104707:3
	wire [69:0] error_slave_req;
	// Trace: design.sv:104708:3
	wire [33:0] error_slave_resp;
	// Trace: design.sv:104710:3
	assign error_slave_resp = 1'sb0;
	// Trace: design.sv:104713:3
	localparam [31:0] core_v_mini_mcu_pkg_CORE_INSTR_IDX = 0;
	assign master_req[0+:70] = core_instr_req_i;
	// Trace: design.sv:104714:3
	localparam [31:0] core_v_mini_mcu_pkg_CORE_DATA_IDX = 1;
	assign master_req[70+:70] = core_data_req_i;
	// Trace: design.sv:104715:3
	localparam [31:0] core_v_mini_mcu_pkg_DEBUG_MASTER_IDX = 2;
	assign master_req[140+:70] = debug_master_req_i;
	// Trace: design.sv:104716:3
	localparam [31:0] core_v_mini_mcu_pkg_DMA_MASTER0_CH0_IDX = 3;
	assign master_req[210+:70] = dma_master0_ch0_req_i;
	// Trace: design.sv:104717:3
	localparam [31:0] core_v_mini_mcu_pkg_DMA_MASTER1_CH0_IDX = 4;
	assign master_req[280+:70] = dma_master1_ch0_req_i;
	// Trace: design.sv:104719:3
	genvar _gv_i_94;
	generate
		for (_gv_i_94 = 0; _gv_i_94 < EXT_XBAR_NMASTER; _gv_i_94 = _gv_i_94 + 1) begin : gen_ext_master_req_map
			localparam i = _gv_i_94;
			// Trace: design.sv:104720:5
			assign master_req[(core_v_mini_mcu_pkg_SYSTEM_XBAR_NMASTER + i) * 70+:70] = ext_xbar_master_req_i[i * 70+:70];
		end
	endgenerate
	// Trace: design.sv:104724:3
	assign core_instr_resp_o = master_resp[0+:34];
	// Trace: design.sv:104725:3
	assign core_data_resp_o = master_resp[34+:34];
	// Trace: design.sv:104726:3
	assign debug_master_resp_o = master_resp[68+:34];
	// Trace: design.sv:104727:3
	assign dma_master0_ch0_resp_o = master_resp[102+:34];
	// Trace: design.sv:104728:3
	assign dma_master1_ch0_resp_o = master_resp[136+:34];
	// Trace: design.sv:104730:3
	genvar _gv_i_95;
	generate
		for (_gv_i_95 = 0; _gv_i_95 < EXT_XBAR_NMASTER; _gv_i_95 = _gv_i_95 + 1) begin : gen_ext_master_resp_map
			localparam i = _gv_i_95;
			// Trace: design.sv:104731:5
			assign ext_xbar_master_resp_o[i * 34+:34] = master_resp[(core_v_mini_mcu_pkg_SYSTEM_XBAR_NMASTER + i) * 34+:34];
		end
	endgenerate
	// Trace: design.sv:104735:3
	localparam [31:0] core_v_mini_mcu_pkg_ERROR_IDX = 32'd0;
	assign error_slave_req = slave_req[0+:70];
	// Trace: design.sv:104736:3
	localparam [31:0] core_v_mini_mcu_pkg_RAM0_IDX = 32'd1;
	assign ram_req_o[0+:70] = slave_req[70+:70];
	// Trace: design.sv:104737:3
	localparam [31:0] core_v_mini_mcu_pkg_RAM1_IDX = 32'd2;
	assign ram_req_o[70+:70] = slave_req[140+:70];
	// Trace: design.sv:104738:3
	localparam [31:0] core_v_mini_mcu_pkg_DEBUG_IDX = 32'd3;
	assign debug_slave_req_o = slave_req[210+:70];
	// Trace: design.sv:104739:3
	localparam [31:0] core_v_mini_mcu_pkg_AO_PERIPHERAL_IDX = 32'd4;
	assign ao_peripheral_slave_req_o = slave_req[280+:70];
	// Trace: design.sv:104740:3
	localparam [31:0] core_v_mini_mcu_pkg_PERIPHERAL_IDX = 32'd5;
	assign peripheral_slave_req_o = slave_req[350+:70];
	// Trace: design.sv:104741:3
	localparam [31:0] core_v_mini_mcu_pkg_FLASH_MEM_IDX = 32'd7;
	assign flash_mem_slave_req_o = slave_req[490+:70];
	// Trace: design.sv:104742:3
	localparam [31:0] core_v_mini_mcu_pkg_EXT_SLAVE_IDX = 32'd6;
	assign ext_xbar_slave_req_o = slave_req[420+:70];
	// Trace: design.sv:104745:3
	assign slave_resp[0+:34] = error_slave_resp;
	// Trace: design.sv:104746:3
	assign slave_resp[34+:34] = ram_resp_i[0+:34];
	// Trace: design.sv:104747:3
	assign slave_resp[68+:34] = ram_resp_i[34+:34];
	// Trace: design.sv:104748:3
	assign slave_resp[102+:34] = debug_slave_resp_i;
	// Trace: design.sv:104749:3
	assign slave_resp[136+:34] = ao_peripheral_slave_resp_i;
	// Trace: design.sv:104750:3
	assign slave_resp[170+:34] = peripheral_slave_resp_i;
	// Trace: design.sv:104751:3
	assign slave_resp[238+:34] = flash_mem_slave_resp_i;
	// Trace: design.sv:104752:3
	assign slave_resp[204+:34] = ext_xbar_slave_resp_i;
	// Trace: design.sv:104771:3
	system_xbar #(
		.XBAR_NMASTER(core_v_mini_mcu_pkg_SYSTEM_XBAR_NMASTER + EXT_XBAR_NMASTER),
		.XBAR_NSLAVE(core_v_mini_mcu_pkg_SYSTEM_XBAR_NSLAVE)
	) system_xbar_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.master_req_i(master_req),
		.master_resp_o(master_resp),
		.slave_req_o(slave_req),
		.slave_resp_i(slave_resp)
	);
endmodule
module system_xbar (
	clk_i,
	rst_ni,
	master_req_i,
	master_resp_o,
	slave_req_o,
	slave_resp_i
);
	// removed import obi_pkg::*;
	// removed import addr_map_rule_pkg::*;
	// removed import core_v_mini_mcu_pkg::*;
	// Trace: design.sv:104793:15
	// removed localparam type core_v_mini_mcu_pkg_bus_type_e
	localparam [0:0] core_v_mini_mcu_pkg_BusType = 1'd1;
	parameter [0:0] BUS_TYPE = core_v_mini_mcu_pkg_BusType;
	// Trace: design.sv:104794:15
	parameter XBAR_NMASTER = 3;
	// Trace: design.sv:104795:15
	parameter XBAR_NSLAVE = 6;
	// Trace: design.sv:104797:5
	input wire clk_i;
	// Trace: design.sv:104798:5
	input wire rst_ni;
	// Trace: design.sv:104800:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [(XBAR_NMASTER * 70) - 1:0] master_req_i;
	// Trace: design.sv:104801:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [(XBAR_NMASTER * 34) - 1:0] master_resp_o;
	// Trace: design.sv:104803:5
	output wire [(XBAR_NSLAVE * 70) - 1:0] slave_req_o;
	// Trace: design.sv:104804:5
	input wire [(XBAR_NSLAVE * 34) - 1:0] slave_resp_i;
	// Trace: design.sv:104808:3
	localparam [31:0] LOG_XBAR_NMASTER = (XBAR_NMASTER > 1 ? $clog2(XBAR_NMASTER) : 32'd1);
	// Trace: design.sv:104809:3
	localparam [31:0] LOG_XBAR_NSLAVE = (XBAR_NSLAVE > 1 ? $clog2(XBAR_NSLAVE) : 32'd1);
	// Trace: design.sv:104813:3
	localparam [31:0] REQ_AGG_DATA_WIDTH = 69;
	// Trace: design.sv:104814:3
	localparam [31:0] RESP_AGG_DATA_WIDTH = 32;
	// Trace: design.sv:104817:3
	wire [(XBAR_NMASTER * LOG_XBAR_NSLAVE) - 1:0] port_sel;
	// Trace: design.sv:104819:3
	wire [LOG_XBAR_NSLAVE - 1:0] port_sel_onetom;
	// Trace: design.sv:104820:3
	wire [0:0] neck_req_req;
	// Trace: design.sv:104821:3
	wire [0:0] neck_resp_gnt;
	// Trace: design.sv:104822:3
	wire [0:0] neck_resp_rvalid;
	// Trace: design.sv:104823:3
	wire [31:0] neck_resp_rdata;
	// Trace: design.sv:104824:3
	wire [69:0] neck_req;
	// Trace: design.sv:104825:3
	wire [68:0] neck_req_out_data;
	// Trace: design.sv:104828:3
	wire [XBAR_NMASTER - 1:0] master_req_req;
	// Trace: design.sv:104829:3
	wire [XBAR_NMASTER - 1:0] master_resp_gnt;
	// Trace: design.sv:104830:3
	wire [XBAR_NMASTER - 1:0] master_resp_rvalid;
	// Trace: design.sv:104831:3
	wire [(XBAR_NMASTER * 32) - 1:0] master_resp_rdata;
	// Trace: design.sv:104833:3
	wire [XBAR_NSLAVE - 1:0] slave_req_req;
	// Trace: design.sv:104834:3
	wire [XBAR_NSLAVE - 1:0] slave_resp_gnt;
	// Trace: design.sv:104835:3
	wire [XBAR_NSLAVE - 1:0] slave_resp_rvalid;
	// Trace: design.sv:104836:3
	wire [(XBAR_NSLAVE * 32) - 1:0] slave_resp_rdata;
	// Trace: design.sv:104839:3
	wire [(XBAR_NMASTER * REQ_AGG_DATA_WIDTH) - 1:0] master_req_out_data;
	// Trace: design.sv:104840:3
	wire [(XBAR_NSLAVE * REQ_AGG_DATA_WIDTH) - 1:0] slave_req_out_data;
	// Trace: design.sv:104842:3
	// removed localparam type addr_map_rule_pkg_addr_map_rule_t
	localparam [31:0] core_v_mini_mcu_pkg_ERROR_IDX = 32'd0;
	localparam [31:0] core_v_mini_mcu_pkg_AO_PERIPHERAL_SIZE = 32'h00100000;
	localparam [31:0] core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS = 32'h20000000;
	localparam [31:0] core_v_mini_mcu_pkg_AO_PERIPHERAL_END_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + core_v_mini_mcu_pkg_AO_PERIPHERAL_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_AO_PERIPHERAL_IDX = 32'd4;
	localparam [31:0] core_v_mini_mcu_pkg_DEBUG_SIZE = 32'h00100000;
	localparam [31:0] core_v_mini_mcu_pkg_DEBUG_START_ADDRESS = 32'h10000000;
	localparam [31:0] core_v_mini_mcu_pkg_DEBUG_END_ADDRESS = core_v_mini_mcu_pkg_DEBUG_START_ADDRESS + core_v_mini_mcu_pkg_DEBUG_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_DEBUG_IDX = 32'd3;
	localparam [31:0] core_v_mini_mcu_pkg_ERROR_SIZE = 32'h00000001;
	localparam [31:0] core_v_mini_mcu_pkg_ERROR_START_ADDRESS = 32'hbadacce5;
	localparam [31:0] core_v_mini_mcu_pkg_ERROR_END_ADDRESS = core_v_mini_mcu_pkg_ERROR_START_ADDRESS + core_v_mini_mcu_pkg_ERROR_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_EXT_SLAVE_SIZE = 32'h01000000;
	localparam [31:0] core_v_mini_mcu_pkg_EXT_SLAVE_START_ADDRESS = 32'hf0000000;
	localparam [31:0] core_v_mini_mcu_pkg_EXT_SLAVE_END_ADDRESS = core_v_mini_mcu_pkg_EXT_SLAVE_START_ADDRESS + core_v_mini_mcu_pkg_EXT_SLAVE_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_EXT_SLAVE_IDX = 32'd6;
	localparam [31:0] core_v_mini_mcu_pkg_FLASH_MEM_SIZE = 32'h01000000;
	localparam [31:0] core_v_mini_mcu_pkg_FLASH_MEM_START_ADDRESS = 32'h40000000;
	localparam [31:0] core_v_mini_mcu_pkg_FLASH_MEM_END_ADDRESS = core_v_mini_mcu_pkg_FLASH_MEM_START_ADDRESS + core_v_mini_mcu_pkg_FLASH_MEM_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_FLASH_MEM_IDX = 32'd7;
	localparam [31:0] core_v_mini_mcu_pkg_PERIPHERAL_SIZE = 32'h00100000;
	localparam [31:0] core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS = 32'h30000000;
	localparam [31:0] core_v_mini_mcu_pkg_PERIPHERAL_END_ADDRESS = core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS + core_v_mini_mcu_pkg_PERIPHERAL_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_PERIPHERAL_IDX = 32'd5;
	localparam [31:0] core_v_mini_mcu_pkg_RAM0_SIZE = 32'h00008000;
	localparam [31:0] core_v_mini_mcu_pkg_RAM0_START_ADDRESS = 32'h00000000;
	localparam [31:0] core_v_mini_mcu_pkg_RAM0_END_ADDRESS = core_v_mini_mcu_pkg_RAM0_START_ADDRESS + core_v_mini_mcu_pkg_RAM0_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_RAM0_IDX = 32'd1;
	localparam [31:0] core_v_mini_mcu_pkg_RAM1_SIZE = 32'h00008000;
	localparam [31:0] core_v_mini_mcu_pkg_RAM1_START_ADDRESS = 32'h00008000;
	localparam [31:0] core_v_mini_mcu_pkg_RAM1_END_ADDRESS = core_v_mini_mcu_pkg_RAM1_START_ADDRESS + core_v_mini_mcu_pkg_RAM1_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_RAM1_IDX = 32'd2;
	localparam core_v_mini_mcu_pkg_SYSTEM_XBAR_NSLAVE = 8;
	localparam [767:0] core_v_mini_mcu_pkg_XBAR_ADDR_RULES = {core_v_mini_mcu_pkg_ERROR_IDX, core_v_mini_mcu_pkg_ERROR_START_ADDRESS, core_v_mini_mcu_pkg_ERROR_END_ADDRESS, core_v_mini_mcu_pkg_RAM0_IDX, core_v_mini_mcu_pkg_RAM0_START_ADDRESS, core_v_mini_mcu_pkg_RAM0_END_ADDRESS, core_v_mini_mcu_pkg_RAM1_IDX, core_v_mini_mcu_pkg_RAM1_START_ADDRESS, core_v_mini_mcu_pkg_RAM1_END_ADDRESS, core_v_mini_mcu_pkg_DEBUG_IDX, core_v_mini_mcu_pkg_DEBUG_START_ADDRESS, core_v_mini_mcu_pkg_DEBUG_END_ADDRESS, core_v_mini_mcu_pkg_AO_PERIPHERAL_IDX, core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS, core_v_mini_mcu_pkg_AO_PERIPHERAL_END_ADDRESS, core_v_mini_mcu_pkg_PERIPHERAL_IDX, core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS, core_v_mini_mcu_pkg_PERIPHERAL_END_ADDRESS, core_v_mini_mcu_pkg_EXT_SLAVE_IDX, core_v_mini_mcu_pkg_EXT_SLAVE_START_ADDRESS, core_v_mini_mcu_pkg_EXT_SLAVE_END_ADDRESS, core_v_mini_mcu_pkg_FLASH_MEM_IDX, core_v_mini_mcu_pkg_FLASH_MEM_START_ADDRESS, core_v_mini_mcu_pkg_FLASH_MEM_END_ADDRESS};
	generate
		if (BUS_TYPE == 1'd0) begin : gen_addr_decoders_NtoM
			genvar _gv_i_96;
			for (_gv_i_96 = 0; _gv_i_96 < XBAR_NMASTER; _gv_i_96 = _gv_i_96 + 1) begin : gen_addr_decoders
				localparam i = _gv_i_96;
				// Trace: design.sv:104844:7
				addr_decode_6EF7A #(
					.NoIndices(XBAR_NSLAVE),
					.NoRules(XBAR_NSLAVE)
				) addr_decode_i(
					.addr_i(master_req_i[(i * 70) + 63-:32]),
					.addr_map_i(core_v_mini_mcu_pkg_XBAR_ADDR_RULES),
					.idx_o(port_sel[i * LOG_XBAR_NSLAVE+:LOG_XBAR_NSLAVE]),
					.dec_valid_o(),
					.dec_error_o(),
					.en_default_idx_i(1'b1),
					.default_idx_i(core_v_mini_mcu_pkg_ERROR_IDX[LOG_XBAR_NSLAVE - 1:0])
				);
			end
		end
	endgenerate
	// Trace: design.sv:104863:3
	genvar _gv_i_97;
	generate
		for (_gv_i_97 = 0; _gv_i_97 < XBAR_NMASTER; _gv_i_97 = _gv_i_97 + 1) begin : gen_unroll_master
			localparam i = _gv_i_97;
			// Trace: design.sv:104864:5
			assign master_req_req[i] = master_req_i[(i * 70) + 69];
			// Trace: design.sv:104865:5
			assign master_req_out_data[i * REQ_AGG_DATA_WIDTH+:REQ_AGG_DATA_WIDTH] = {master_req_i[(i * 70) + 68], master_req_i[(i * 70) + 67-:4], master_req_i[(i * 70) + 63-:32], master_req_i[(i * 70) + 31-:32]};
			// Trace: design.sv:104868:5
			assign master_resp_o[(i * 34) + 33] = master_resp_gnt[i];
			// Trace: design.sv:104869:5
			assign master_resp_o[(i * 34) + 31-:32] = master_resp_rdata[i * 32+:32];
			// Trace: design.sv:104870:5
			assign master_resp_o[(i * 34) + 32] = master_resp_rvalid[i];
		end
	endgenerate
	// Trace: design.sv:104872:3
	genvar _gv_i_98;
	generate
		for (_gv_i_98 = 0; _gv_i_98 < XBAR_NSLAVE; _gv_i_98 = _gv_i_98 + 1) begin : gen_unroll_slave
			localparam i = _gv_i_98;
			// Trace: design.sv:104873:5
			assign slave_req_o[(i * 70) + 69] = slave_req_req[i];
			// Trace: design.sv:104874:5
			assign {slave_req_o[(i * 70) + 68], slave_req_o[(i * 70) + 67-:4], slave_req_o[(i * 70) + 63-:32], slave_req_o[(i * 70) + 31-:32]} = slave_req_out_data[i * REQ_AGG_DATA_WIDTH+:REQ_AGG_DATA_WIDTH];
			// Trace: design.sv:104875:5
			assign slave_resp_rdata[i * 32+:32] = slave_resp_i[(i * 34) + 31-:32];
			// Trace: design.sv:104876:5
			assign slave_resp_gnt[i] = slave_resp_i[(i * 34) + 33];
			// Trace: design.sv:104877:5
			assign slave_resp_rvalid[i] = slave_resp_i[(i * 34) + 32];
		end
	endgenerate
	// Trace: design.sv:104881:3
	generate
		if (BUS_TYPE == 1'd0) begin : gen_xbar_NtoM
			// Trace: design.sv:104884:5
			localparam [31:0] sv2v_uu_i_xbar_NumIn = XBAR_NMASTER;
			localparam [31:0] sv2v_uu_i_xbar_LogNumIn = (sv2v_uu_i_xbar_NumIn > 1 ? $clog2(sv2v_uu_i_xbar_NumIn) : 1);
			localparam [31:0] sv2v_uu_i_xbar_NumOut = XBAR_NSLAVE;
			// removed localparam type sv2v_uu_i_xbar_rr_i
			localparam [(sv2v_uu_i_xbar_NumOut * sv2v_uu_i_xbar_LogNumIn) - 1:0] sv2v_uu_i_xbar_ext_rr_i_0 = 1'sb0;
			xbar_varlat #(
				.AggregateGnt(1),
				.NumIn(XBAR_NMASTER),
				.NumOut(XBAR_NSLAVE),
				.ReqDataWidth(REQ_AGG_DATA_WIDTH),
				.RespDataWidth(RESP_AGG_DATA_WIDTH)
			) i_xbar(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(master_req_req),
				.add_i(port_sel),
				.wdata_i(master_req_out_data),
				.gnt_o(master_resp_gnt),
				.rdata_o(master_resp_rdata),
				.rr_i(sv2v_uu_i_xbar_ext_rr_i_0),
				.vld_o(master_resp_rvalid),
				.gnt_i(slave_resp_gnt),
				.req_o(slave_req_req),
				.vld_i(slave_resp_rvalid),
				.wdata_o(slave_req_out_data),
				.rdata_i(slave_resp_rdata)
			);
		end
		else begin : gen_xbar_1toM
			// Trace: design.sv:104910:5
			localparam [31:0] sv2v_uu_i_xbar_master_NumOut = 1;
			localparam [31:0] sv2v_uu_i_xbar_master_LogNumOut = 1;
			localparam [31:0] sv2v_uu_i_xbar_master_NumIn = XBAR_NMASTER;
			// removed localparam type sv2v_uu_i_xbar_master_add_i
			localparam [(sv2v_uu_i_xbar_master_NumIn * sv2v_uu_i_xbar_master_LogNumOut) - 1:0] sv2v_uu_i_xbar_master_ext_add_i_0 = 1'sb0;
			localparam [31:0] sv2v_uu_i_xbar_master_LogNumIn = (sv2v_uu_i_xbar_master_NumIn > 1 ? $clog2(sv2v_uu_i_xbar_master_NumIn) : 1);
			// removed localparam type sv2v_uu_i_xbar_master_rr_i
			localparam [(sv2v_uu_i_xbar_master_NumOut * sv2v_uu_i_xbar_master_LogNumIn) - 1:0] sv2v_uu_i_xbar_master_ext_rr_i_0 = 1'sb0;
			xbar_varlat #(
				.NumIn(XBAR_NMASTER),
				.NumOut(1),
				.ReqDataWidth(REQ_AGG_DATA_WIDTH),
				.RespDataWidth(RESP_AGG_DATA_WIDTH)
			) i_xbar_master(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(master_req_req),
				.add_i(sv2v_uu_i_xbar_master_ext_add_i_0),
				.wdata_i(master_req_out_data),
				.gnt_o(master_resp_gnt),
				.rdata_o(master_resp_rdata),
				.rr_i(sv2v_uu_i_xbar_master_ext_rr_i_0),
				.vld_o(master_resp_rvalid),
				.gnt_i(neck_resp_gnt),
				.req_o(neck_req_req),
				.vld_i(neck_resp_rvalid),
				.wdata_o(neck_req_out_data),
				.rdata_i(neck_resp_rdata)
			);
			// Trace: design.sv:104932:5
			assign {neck_req[68], neck_req[67-:4], neck_req[63-:32], neck_req[31-:32]} = neck_req_out_data[0+:REQ_AGG_DATA_WIDTH];
			// Trace: design.sv:104934:5
			addr_decode_6EF7A #(
				.NoIndices(XBAR_NSLAVE),
				.NoRules(XBAR_NSLAVE)
			) addr_decode_i(
				.addr_i(neck_req[63-:32]),
				.addr_map_i(core_v_mini_mcu_pkg_XBAR_ADDR_RULES),
				.idx_o(port_sel_onetom[0+:LOG_XBAR_NSLAVE]),
				.dec_valid_o(),
				.dec_error_o(),
				.en_default_idx_i(1'b1),
				.default_idx_i(core_v_mini_mcu_pkg_ERROR_IDX[LOG_XBAR_NSLAVE - 1:0])
			);
			// Trace: design.sv:104951:5
			localparam [31:0] sv2v_uu_i_xbar_slave_NumIn = 1;
			localparam [31:0] sv2v_uu_i_xbar_slave_LogNumIn = 1;
			localparam [31:0] sv2v_uu_i_xbar_slave_NumOut = XBAR_NSLAVE;
			// removed localparam type sv2v_uu_i_xbar_slave_rr_i
			localparam [(sv2v_uu_i_xbar_slave_NumOut * sv2v_uu_i_xbar_slave_LogNumIn) - 1:0] sv2v_uu_i_xbar_slave_ext_rr_i_0 = 1'sb0;
			xbar_varlat #(
				.AggregateGnt(0),
				.NumIn(1),
				.NumOut(XBAR_NSLAVE),
				.ReqDataWidth(REQ_AGG_DATA_WIDTH),
				.RespDataWidth(RESP_AGG_DATA_WIDTH)
			) i_xbar_slave(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(neck_req_req),
				.add_i(port_sel_onetom[0+:LOG_XBAR_NSLAVE]),
				.wdata_i(neck_req_out_data),
				.gnt_o(neck_resp_gnt),
				.rdata_o(neck_resp_rdata),
				.rr_i(sv2v_uu_i_xbar_slave_ext_rr_i_0),
				.vld_o(neck_resp_rvalid),
				.gnt_i(slave_resp_gnt),
				.req_o(slave_req_req),
				.vld_i(slave_resp_rvalid),
				.wdata_o(slave_req_out_data),
				.rdata_i(slave_resp_rdata)
			);
		end
	endgenerate
endmodule
module spi_subsystem (
	clk_i,
	rst_ni,
	use_spimemio_i,
	spimemio_req_i,
	spimemio_resp_o,
	yo_reg_req_i,
	yo_reg_rsp_o,
	ot_reg_req_i,
	ot_reg_rsp_o,
	spi_flash_sck_o,
	spi_flash_sck_en_o,
	spi_flash_csb_o,
	spi_flash_csb_en_o,
	spi_flash_sd_o,
	spi_flash_sd_en_o,
	spi_flash_sd_i,
	spi_flash_intr_error_o,
	spi_flash_intr_event_o,
	spi_flash_rx_valid_o,
	spi_flash_tx_ready_o
);
	reg _sv2v_0;
	// removed import obi_pkg::*;
	// removed import reg_pkg::*;
	// Trace: design.sv:104992:5
	input wire clk_i;
	// Trace: design.sv:104993:5
	input wire rst_ni;
	// Trace: design.sv:104995:5
	input wire use_spimemio_i;
	// Trace: design.sv:104998:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [69:0] spimemio_req_i;
	// Trace: design.sv:104999:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [33:0] spimemio_resp_o;
	// Trace: design.sv:105001:5
	// removed localparam type reg_pkg_reg_req_t
	input wire [69:0] yo_reg_req_i;
	// Trace: design.sv:105002:5
	// removed localparam type reg_pkg_reg_rsp_t
	output wire [33:0] yo_reg_rsp_o;
	// Trace: design.sv:105005:5
	input wire [69:0] ot_reg_req_i;
	// Trace: design.sv:105006:5
	output wire [33:0] ot_reg_rsp_o;
	// Trace: design.sv:105009:5
	output reg spi_flash_sck_o;
	// Trace: design.sv:105010:5
	output reg spi_flash_sck_en_o;
	// Trace: design.sv:105011:5
	localparam signed [31:0] spi_host_reg_pkg_NumCS = 2;
	output reg [1:0] spi_flash_csb_o;
	// Trace: design.sv:105012:5
	output reg [1:0] spi_flash_csb_en_o;
	// Trace: design.sv:105013:5
	output reg [3:0] spi_flash_sd_o;
	// Trace: design.sv:105014:5
	output reg [3:0] spi_flash_sd_en_o;
	// Trace: design.sv:105015:5
	input wire [3:0] spi_flash_sd_i;
	// Trace: design.sv:105018:5
	output reg spi_flash_intr_error_o;
	// Trace: design.sv:105019:5
	output reg spi_flash_intr_event_o;
	// Trace: design.sv:105022:5
	output reg spi_flash_rx_valid_o;
	// Trace: design.sv:105023:5
	output reg spi_flash_tx_ready_o;
	// Trace: design.sv:105027:3
	wire ot_spi_sck;
	// Trace: design.sv:105028:3
	wire ot_spi_sck_en;
	// Trace: design.sv:105029:3
	wire [1:0] ot_spi_csb;
	// Trace: design.sv:105030:3
	wire [1:0] ot_spi_csb_en;
	// Trace: design.sv:105031:3
	wire [3:0] ot_spi_sd_out;
	// Trace: design.sv:105032:3
	wire [3:0] ot_spi_sd_en;
	// Trace: design.sv:105033:3
	reg [3:0] ot_spi_sd_in;
	// Trace: design.sv:105034:3
	wire ot_spi_intr_error;
	// Trace: design.sv:105035:3
	wire ot_spi_intr_event;
	// Trace: design.sv:105036:3
	wire ot_spi_rx_valid;
	// Trace: design.sv:105037:3
	wire ot_spi_tx_ready;
	// Trace: design.sv:105040:3
	wire yo_spi_sck;
	// Trace: design.sv:105041:3
	wire yo_spi_sck_en;
	// Trace: design.sv:105042:3
	wire [1:0] yo_spi_csb;
	// Trace: design.sv:105043:3
	wire [1:0] yo_spi_csb_en;
	// Trace: design.sv:105044:3
	wire [3:0] yo_spi_sd_out;
	// Trace: design.sv:105045:3
	wire [3:0] yo_spi_sd_en;
	// Trace: design.sv:105046:3
	reg [3:0] yo_spi_sd_in;
	// Trace: design.sv:105049:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:105050:5
		if (!use_spimemio_i) begin
			// Trace: design.sv:105051:7
			spi_flash_sck_o = ot_spi_sck;
			// Trace: design.sv:105052:7
			spi_flash_sck_en_o = ot_spi_sck_en;
			// Trace: design.sv:105053:7
			spi_flash_csb_o = ot_spi_csb;
			// Trace: design.sv:105054:7
			spi_flash_csb_en_o = ot_spi_csb_en;
			// Trace: design.sv:105055:7
			spi_flash_sd_o = ot_spi_sd_out;
			// Trace: design.sv:105056:7
			spi_flash_sd_en_o = ot_spi_sd_en;
			// Trace: design.sv:105057:7
			ot_spi_sd_in = spi_flash_sd_i;
			// Trace: design.sv:105058:7
			yo_spi_sd_in = 1'sb0;
			// Trace: design.sv:105059:7
			spi_flash_intr_error_o = ot_spi_intr_error;
			// Trace: design.sv:105060:7
			spi_flash_intr_event_o = ot_spi_intr_event;
			// Trace: design.sv:105061:7
			spi_flash_rx_valid_o = ot_spi_rx_valid;
			// Trace: design.sv:105062:7
			spi_flash_tx_ready_o = ot_spi_tx_ready;
		end
		else begin
			// Trace: design.sv:105064:7
			spi_flash_sck_o = yo_spi_sck;
			// Trace: design.sv:105065:7
			spi_flash_sck_en_o = yo_spi_sck_en;
			// Trace: design.sv:105066:7
			spi_flash_csb_o = yo_spi_csb;
			// Trace: design.sv:105067:7
			spi_flash_csb_en_o = yo_spi_csb_en;
			// Trace: design.sv:105068:7
			spi_flash_sd_o = yo_spi_sd_out;
			// Trace: design.sv:105069:7
			spi_flash_sd_en_o = yo_spi_sd_en;
			// Trace: design.sv:105070:7
			ot_spi_sd_in = 1'sb0;
			// Trace: design.sv:105071:7
			yo_spi_sd_in = spi_flash_sd_i;
			// Trace: design.sv:105072:7
			spi_flash_intr_error_o = 1'b0;
			// Trace: design.sv:105073:7
			spi_flash_intr_event_o = 1'b0;
			// Trace: design.sv:105074:7
			spi_flash_rx_valid_o = 1'b0;
			// Trace: design.sv:105075:7
			spi_flash_tx_ready_o = 1'b0;
		end
	end
	// Trace: design.sv:105080:3
	assign yo_spi_sck_en = 1'b1;
	// Trace: design.sv:105081:3
	assign yo_spi_csb_en = 2'b01;
	// Trace: design.sv:105082:3
	assign yo_spi_csb[1] = 1'b1;
	// Trace: design.sv:105084:3
	obi_spimemio obi_spimemio_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flash_csb_o(yo_spi_csb[0]),
		.flash_clk_o(yo_spi_sck),
		.flash_io0_oe_o(yo_spi_sd_en[0]),
		.flash_io1_oe_o(yo_spi_sd_en[1]),
		.flash_io2_oe_o(yo_spi_sd_en[2]),
		.flash_io3_oe_o(yo_spi_sd_en[3]),
		.flash_io0_do_o(yo_spi_sd_out[0]),
		.flash_io1_do_o(yo_spi_sd_out[1]),
		.flash_io2_do_o(yo_spi_sd_out[2]),
		.flash_io3_do_o(yo_spi_sd_out[3]),
		.flash_io0_di_i(yo_spi_sd_in[0]),
		.flash_io1_di_i(yo_spi_sd_in[1]),
		.flash_io2_di_i(yo_spi_sd_in[2]),
		.flash_io3_di_i(yo_spi_sd_in[3]),
		.reg_req_i(yo_reg_req_i),
		.reg_rsp_o(yo_reg_rsp_o),
		.spimemio_req_i(spimemio_req_i),
		.spimemio_resp_o(spimemio_resp_o)
	);
	// Trace: design.sv:105108:3
	// removed localparam type spi_device_pkg_passthrough_req_t
	localparam [13:0] spi_device_pkg_PASSTHROUGH_REQ_DEFAULT = 14'h0200;
	spi_host_CA356 ot_spi_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(ot_reg_req_i),
		.reg_rsp_o(ot_reg_rsp_o),
		.alert_rx_i(),
		.alert_tx_o(),
		.passthrough_i(spi_device_pkg_PASSTHROUGH_REQ_DEFAULT),
		.passthrough_o(),
		.cio_sck_o(ot_spi_sck),
		.cio_sck_en_o(ot_spi_sck_en),
		.cio_csb_o(ot_spi_csb),
		.cio_csb_en_o(ot_spi_csb_en),
		.cio_sd_o(ot_spi_sd_out),
		.cio_sd_en_o(ot_spi_sd_en),
		.cio_sd_i(ot_spi_sd_in),
		.rx_valid_o(ot_spi_rx_valid),
		.tx_ready_o(ot_spi_tx_ready),
		.intr_error_o(ot_spi_intr_error),
		.intr_spi_event_o(ot_spi_intr_event)
	);
	initial _sv2v_0 = 0;
endmodule
module debug_subsystem (
	clk_i,
	rst_ni,
	jtag_tck_i,
	jtag_tms_i,
	jtag_trst_ni,
	jtag_tdi_i,
	jtag_tdo_o,
	debug_core_req_o,
	debug_slave_req_i,
	debug_slave_resp_o,
	debug_master_req_o,
	debug_master_resp_i
);
	// removed import obi_pkg::*;
	// Trace: design.sv:105152:15
	parameter JTAG_IDCODE = 32'h10001c05;
	// Trace: design.sv:105154:5
	input wire clk_i;
	// Trace: design.sv:105155:5
	input wire rst_ni;
	// Trace: design.sv:105157:5
	input wire jtag_tck_i;
	// Trace: design.sv:105158:5
	input wire jtag_tms_i;
	// Trace: design.sv:105159:5
	input wire jtag_trst_ni;
	// Trace: design.sv:105160:5
	input wire jtag_tdi_i;
	// Trace: design.sv:105161:5
	output wire jtag_tdo_o;
	// Trace: design.sv:105163:5
	output wire debug_core_req_o;
	// Trace: design.sv:105165:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [69:0] debug_slave_req_i;
	// Trace: design.sv:105166:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [33:0] debug_slave_resp_o;
	// Trace: design.sv:105167:5
	output wire [69:0] debug_master_req_o;
	// Trace: design.sv:105168:5
	input wire [33:0] debug_master_resp_i;
	// Trace: design.sv:105172:3
	// removed import dm::*;
	// Trace: design.sv:105174:3
	localparam [11:0] dm_DataAddr = 12'h380;
	localparam [3:0] dm_DataCount = 4'h2;
	// removed localparam type dm_hartinfo_t
	localparam [31:0] hartinfo = {16'h0021, dm_DataCount, dm_DataAddr};
	// Trace: design.sv:105183:3
	// removed localparam type dm_dtm_op_e
	// removed localparam type dm_dmi_req_t
	wire [40:0] dmi_req;
	// Trace: design.sv:105184:3
	wire dmi_req_valid;
	// Trace: design.sv:105185:3
	wire dmi_req_ready;
	// Trace: design.sv:105186:3
	// removed localparam type dm_dmi_resp_t
	wire [33:0] dmi_resp;
	// Trace: design.sv:105187:3
	wire dmi_resp_ready;
	// Trace: design.sv:105188:3
	wire dmi_resp_valid;
	// Trace: design.sv:105191:3
	dmi_jtag #(.IdcodeValue(JTAG_IDCODE)) dmi_jtag_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.testmode_i(1'b0),
		.dmi_req_o(dmi_req),
		.dmi_req_valid_o(dmi_req_valid),
		.dmi_req_ready_i(dmi_req_ready),
		.dmi_resp_i(dmi_resp),
		.dmi_resp_ready_o(dmi_resp_ready),
		.dmi_resp_valid_i(dmi_resp_valid),
		.dmi_rst_no(),
		.tck_i(jtag_tck_i),
		.tms_i(jtag_tms_i),
		.trst_ni(jtag_trst_ni),
		.td_i(jtag_tdi_i),
		.td_o(jtag_tdo_o),
		.tdo_oe_o()
	);
	// Trace: design.sv:105212:3
	localparam [31:0] sv2v_uu_dm_obi_top_i_IdWidth = 1;
	// removed localparam type sv2v_uu_dm_obi_top_i_slave_aid_i
	localparam [0:0] sv2v_uu_dm_obi_top_i_ext_slave_aid_i_0 = 1'sb0;
	dm_obi_top dm_obi_top_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.testmode_i(1'b0),
		.ndmreset_o(),
		.dmactive_o(),
		.debug_req_o(debug_core_req_o),
		.unavailable_i(~1'b1),
		.hartinfo_i(hartinfo),
		.slave_req_i(debug_slave_req_i[69]),
		.slave_gnt_o(debug_slave_resp_o[33]),
		.slave_we_i(debug_slave_req_i[68]),
		.slave_addr_i(debug_slave_req_i[63-:32]),
		.slave_be_i(debug_slave_req_i[67-:4]),
		.slave_wdata_i(debug_slave_req_i[31-:32]),
		.slave_aid_i(sv2v_uu_dm_obi_top_i_ext_slave_aid_i_0),
		.slave_rdata_o(debug_slave_resp_o[31-:32]),
		.slave_rvalid_o(debug_slave_resp_o[32]),
		.slave_rid_o(),
		.master_req_o(debug_master_req_o[69]),
		.master_addr_o(debug_master_req_o[63-:32]),
		.master_we_o(debug_master_req_o[68]),
		.master_wdata_o(debug_master_req_o[31-:32]),
		.master_be_o(debug_master_req_o[67-:4]),
		.master_gnt_i(debug_master_resp_i[33]),
		.master_rvalid_i(debug_master_resp_i[32]),
		.master_err_i(1'b0),
		.master_other_err_i(1'b0),
		.master_rdata_i(debug_master_resp_i[31-:32]),
		.dmi_rst_ni(rst_ni),
		.dmi_req_valid_i(dmi_req_valid),
		.dmi_req_ready_o(dmi_req_ready),
		.dmi_req_i(dmi_req),
		.dmi_resp_valid_o(dmi_resp_valid),
		.dmi_resp_ready_i(dmi_resp_ready),
		.dmi_resp_o(dmi_resp)
	);
endmodule
module peripheral_subsystem (
	clk_i,
	rst_ni,
	clk_gate_en_i,
	slave_req_i,
	slave_resp_o,
	intr_vector_ext_i,
	irq_plic_o,
	msip_o,
	uart_intr_tx_watermark_i,
	uart_intr_rx_watermark_i,
	uart_intr_tx_empty_i,
	uart_intr_rx_overflow_i,
	uart_intr_rx_frame_err_i,
	uart_intr_rx_break_err_i,
	uart_intr_rx_timeout_i,
	uart_intr_rx_parity_err_i,
	cio_gpio_i,
	cio_gpio_o,
	cio_gpio_en_o,
	cio_scl_i,
	cio_scl_o,
	cio_scl_en_o,
	cio_sda_i,
	cio_sda_o,
	cio_sda_en_o,
	spi2_sck_o,
	spi2_sck_en_o,
	spi2_csb_o,
	spi2_csb_en_o,
	spi2_sd_o,
	spi2_sd_en_o,
	spi2_sd_i,
	rv_timer_2_intr_o,
	rv_timer_3_intr_o
);
	// removed import obi_pkg::*;
	// removed import reg_pkg::*;
	// Trace: design.sv:105262:15
	parameter NEXT_INT = 0;
	// Trace: design.sv:105264:5
	input wire clk_i;
	// Trace: design.sv:105265:5
	input wire rst_ni;
	// Trace: design.sv:105268:5
	input wire clk_gate_en_i;
	// Trace: design.sv:105270:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [69:0] slave_req_i;
	// Trace: design.sv:105271:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [33:0] slave_resp_o;
	// Trace: design.sv:105274:5
	input wire [NEXT_INT - 1:0] intr_vector_ext_i;
	// Trace: design.sv:105275:5
	output wire irq_plic_o;
	// Trace: design.sv:105276:5
	output wire msip_o;
	// Trace: design.sv:105279:5
	input wire uart_intr_tx_watermark_i;
	// Trace: design.sv:105280:5
	input wire uart_intr_rx_watermark_i;
	// Trace: design.sv:105281:5
	input wire uart_intr_tx_empty_i;
	// Trace: design.sv:105282:5
	input wire uart_intr_rx_overflow_i;
	// Trace: design.sv:105283:5
	input wire uart_intr_rx_frame_err_i;
	// Trace: design.sv:105284:5
	input wire uart_intr_rx_break_err_i;
	// Trace: design.sv:105285:5
	input wire uart_intr_rx_timeout_i;
	// Trace: design.sv:105286:5
	input wire uart_intr_rx_parity_err_i;
	// Trace: design.sv:105289:5
	input wire [31:8] cio_gpio_i;
	// Trace: design.sv:105290:5
	output wire [31:8] cio_gpio_o;
	// Trace: design.sv:105291:5
	output wire [31:8] cio_gpio_en_o;
	// Trace: design.sv:105294:5
	input wire cio_scl_i;
	// Trace: design.sv:105295:5
	output wire cio_scl_o;
	// Trace: design.sv:105296:5
	output wire cio_scl_en_o;
	// Trace: design.sv:105297:5
	input wire cio_sda_i;
	// Trace: design.sv:105298:5
	output wire cio_sda_o;
	// Trace: design.sv:105299:5
	output wire cio_sda_en_o;
	// Trace: design.sv:105302:5
	output wire spi2_sck_o;
	// Trace: design.sv:105303:5
	output wire spi2_sck_en_o;
	// Trace: design.sv:105304:5
	localparam signed [31:0] spi_host_reg_pkg_NumCS = 2;
	output wire [1:0] spi2_csb_o;
	// Trace: design.sv:105305:5
	output wire [1:0] spi2_csb_en_o;
	// Trace: design.sv:105306:5
	output wire [3:0] spi2_sd_o;
	// Trace: design.sv:105307:5
	output wire [3:0] spi2_sd_en_o;
	// Trace: design.sv:105308:5
	input wire [3:0] spi2_sd_i;
	// Trace: design.sv:105311:5
	output wire rv_timer_2_intr_o;
	// Trace: design.sv:105312:5
	output wire rv_timer_3_intr_o;
	// Trace: design.sv:105315:3
	// removed import core_v_mini_mcu_pkg::*;
	// Trace: design.sv:105316:3
	// removed import tlul_pkg::*;
	// Trace: design.sv:105317:3
	// removed import rv_plic_reg_pkg::*;
	// Trace: design.sv:105319:3
	// removed localparam type reg_pkg_reg_req_t
	wire [69:0] peripheral_req;
	// Trace: design.sv:105320:3
	// removed localparam type reg_pkg_reg_rsp_t
	wire [33:0] peripheral_rsp;
	// Trace: design.sv:105322:3
	localparam core_v_mini_mcu_pkg_PERIPHERALS = 5;
	wire [349:0] peripheral_slv_req;
	// Trace: design.sv:105323:3
	wire [169:0] peripheral_slv_rsp;
	// Trace: design.sv:105325:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] plic_tl_h2d;
	// Trace: design.sv:105326:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] plic_tl_d2h;
	// Trace: design.sv:105328:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] i2c_tl_h2d;
	// Trace: design.sv:105329:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] i2c_tl_d2h;
	// Trace: design.sv:105331:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] rv_timer_tl_h2d;
	// Trace: design.sv:105332:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] rv_timer_tl_d2h;
	// Trace: design.sv:105334:3
	localparam signed [31:0] rv_plic_reg_pkg_NumTarget = 1;
	wire [0:0] irq_plic;
	// Trace: design.sv:105335:3
	localparam signed [31:0] rv_plic_reg_pkg_NumSrc = 64;
	wire [63:0] intr_vector;
	// Trace: design.sv:105336:3
	wire [5:0] irq_id;
	// Trace: design.sv:105337:3
	wire [5:0] unused_irq_id;
	// Trace: design.sv:105339:3
	wire [31:8] gpio_intr;
	// Trace: design.sv:105340:3
	wire [7:0] cio_gpio_unused;
	// Trace: design.sv:105341:3
	wire [7:0] cio_gpio_en_unused;
	// Trace: design.sv:105342:3
	wire [7:0] gpio_int_unused;
	// Trace: design.sv:105344:3
	wire i2c_intr_fmt_watermark;
	// Trace: design.sv:105345:3
	wire i2c_intr_rx_watermark;
	// Trace: design.sv:105346:3
	wire i2c_intr_fmt_overflow;
	// Trace: design.sv:105347:3
	wire i2c_intr_rx_overflow;
	// Trace: design.sv:105348:3
	wire i2c_intr_nak;
	// Trace: design.sv:105349:3
	wire i2c_intr_scl_interference;
	// Trace: design.sv:105350:3
	wire i2c_intr_sda_interference;
	// Trace: design.sv:105351:3
	wire i2c_intr_stretch_timeout;
	// Trace: design.sv:105352:3
	wire i2c_intr_sda_unstable;
	// Trace: design.sv:105353:3
	wire i2c_intr_trans_complete;
	// Trace: design.sv:105354:3
	wire i2c_intr_tx_empty;
	// Trace: design.sv:105355:3
	wire i2c_intr_tx_nonempty;
	// Trace: design.sv:105356:3
	wire i2c_intr_tx_overflow;
	// Trace: design.sv:105357:3
	wire i2c_intr_acq_overflow;
	// Trace: design.sv:105358:3
	wire i2c_intr_ack_stop;
	// Trace: design.sv:105359:3
	wire i2c_intr_host_timeout;
	// Trace: design.sv:105360:3
	wire spi2_intr_event;
	// Trace: design.sv:105363:3
	assign unused_irq_id = irq_id;
	// Trace: design.sv:105366:3
	assign intr_vector[0] = 1'b0;
	// Trace: design.sv:105367:3
	assign intr_vector[1] = uart_intr_tx_watermark_i;
	// Trace: design.sv:105368:3
	assign intr_vector[2] = uart_intr_rx_watermark_i;
	// Trace: design.sv:105369:3
	assign intr_vector[3] = uart_intr_tx_empty_i;
	// Trace: design.sv:105370:3
	assign intr_vector[4] = uart_intr_rx_overflow_i;
	// Trace: design.sv:105371:3
	assign intr_vector[5] = uart_intr_rx_frame_err_i;
	// Trace: design.sv:105372:3
	assign intr_vector[6] = uart_intr_rx_break_err_i;
	// Trace: design.sv:105373:3
	assign intr_vector[7] = uart_intr_rx_timeout_i;
	// Trace: design.sv:105374:3
	assign intr_vector[8] = uart_intr_rx_parity_err_i;
	// Trace: design.sv:105375:3
	assign intr_vector[32:9] = gpio_intr;
	// Trace: design.sv:105376:3
	assign intr_vector[33] = i2c_intr_fmt_watermark;
	// Trace: design.sv:105377:3
	assign intr_vector[34] = i2c_intr_rx_watermark;
	// Trace: design.sv:105378:3
	assign intr_vector[35] = i2c_intr_fmt_overflow;
	// Trace: design.sv:105379:3
	assign intr_vector[36] = i2c_intr_rx_overflow;
	// Trace: design.sv:105380:3
	assign intr_vector[37] = i2c_intr_nak;
	// Trace: design.sv:105381:3
	assign intr_vector[38] = i2c_intr_scl_interference;
	// Trace: design.sv:105382:3
	assign intr_vector[39] = i2c_intr_sda_interference;
	// Trace: design.sv:105383:3
	assign intr_vector[40] = i2c_intr_stretch_timeout;
	// Trace: design.sv:105384:3
	assign intr_vector[41] = i2c_intr_sda_unstable;
	// Trace: design.sv:105385:3
	assign intr_vector[42] = i2c_intr_trans_complete;
	// Trace: design.sv:105386:3
	assign intr_vector[43] = i2c_intr_tx_empty;
	// Trace: design.sv:105387:3
	assign intr_vector[44] = i2c_intr_tx_nonempty;
	// Trace: design.sv:105388:3
	assign intr_vector[45] = i2c_intr_tx_overflow;
	// Trace: design.sv:105389:3
	assign intr_vector[46] = i2c_intr_acq_overflow;
	// Trace: design.sv:105390:3
	assign intr_vector[47] = i2c_intr_ack_stop;
	// Trace: design.sv:105391:3
	assign intr_vector[48] = i2c_intr_host_timeout;
	// Trace: design.sv:105392:3
	assign intr_vector[49] = spi2_intr_event;
	// Trace: design.sv:105395:3
	genvar _gv_i_99;
	localparam core_v_mini_mcu_pkg_PLIC_USED_NINT = 50;
	generate
		for (_gv_i_99 = 0; _gv_i_99 < NEXT_INT; _gv_i_99 = _gv_i_99 + 1) begin : genblk1
			localparam i = _gv_i_99;
			// Trace: design.sv:105396:5
			assign intr_vector[i + core_v_mini_mcu_pkg_PLIC_USED_NINT] = intr_vector_ext_i[i];
		end
	endgenerate
	// Trace: design.sv:105400:3
	localparam [31:0] core_v_mini_mcu_pkg_PERIPHERALS_PORT_SEL_WIDTH = 3;
	wire [2:0] peripheral_select;
	// Trace: design.sv:105403:3
	wire clk_cg;
	// Trace: design.sv:105404:3
	tc_clk_gating clk_gating_cell(
		.clk_i(clk_i),
		.en_i(~clk_gate_en_i),
		.test_en_i(1'b0),
		.clk_o(clk_cg)
	);
	// Trace: design.sv:105411:3
	localparam [31:0] sv2v_uu_periph_to_reg_i_IW = 1;
	// removed localparam type sv2v_uu_periph_to_reg_i_id_i
	localparam [0:0] sv2v_uu_periph_to_reg_i_ext_id_i_0 = 1'sb0;
	periph_to_reg_35129 #(.IW(1)) periph_to_reg_i(
		.clk_i(clk_cg),
		.rst_ni(rst_ni),
		.req_i(slave_req_i[69]),
		.add_i(slave_req_i[63-:32]),
		.wen_i(~slave_req_i[68]),
		.wdata_i(slave_req_i[31-:32]),
		.be_i(slave_req_i[67-:4]),
		.id_i(sv2v_uu_periph_to_reg_i_ext_id_i_0),
		.gnt_o(slave_resp_o[33]),
		.r_rdata_o(slave_resp_o[31-:32]),
		.r_opc_o(),
		.r_id_o(),
		.r_valid_o(slave_resp_o[32]),
		.reg_req_o(peripheral_req),
		.reg_rsp_i(peripheral_rsp)
	);
	// Trace: design.sv:105433:3
	// removed localparam type addr_map_rule_pkg_addr_map_rule_t
	localparam [31:0] core_v_mini_mcu_pkg_GPIO_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS = 32'h30000000;
	localparam [31:0] core_v_mini_mcu_pkg_GPIO_START_ADDRESS = core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS + 32'h00020000;
	localparam [31:0] core_v_mini_mcu_pkg_GPIO_END_ADDRESS = core_v_mini_mcu_pkg_GPIO_START_ADDRESS + core_v_mini_mcu_pkg_GPIO_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_GPIO_IDX = 32'd1;
	localparam [31:0] core_v_mini_mcu_pkg_I2C_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_I2C_START_ADDRESS = core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS + 32'h00030000;
	localparam [31:0] core_v_mini_mcu_pkg_I2C_END_ADDRESS = core_v_mini_mcu_pkg_I2C_START_ADDRESS + core_v_mini_mcu_pkg_I2C_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_I2C_IDX = 32'd2;
	localparam [31:0] core_v_mini_mcu_pkg_RV_PLIC_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_RV_PLIC_START_ADDRESS = core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS + 32'h00000000;
	localparam [31:0] core_v_mini_mcu_pkg_RV_PLIC_END_ADDRESS = core_v_mini_mcu_pkg_RV_PLIC_START_ADDRESS + core_v_mini_mcu_pkg_RV_PLIC_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_RV_PLIC_IDX = 32'd0;
	localparam [31:0] core_v_mini_mcu_pkg_RV_TIMER_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_RV_TIMER_START_ADDRESS = core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS + 32'h00040000;
	localparam [31:0] core_v_mini_mcu_pkg_RV_TIMER_END_ADDRESS = core_v_mini_mcu_pkg_RV_TIMER_START_ADDRESS + core_v_mini_mcu_pkg_RV_TIMER_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_RV_TIMER_IDX = 32'd3;
	localparam [31:0] core_v_mini_mcu_pkg_SPI2_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_SPI2_START_ADDRESS = core_v_mini_mcu_pkg_PERIPHERAL_START_ADDRESS + 32'h00050000;
	localparam [31:0] core_v_mini_mcu_pkg_SPI2_END_ADDRESS = core_v_mini_mcu_pkg_SPI2_START_ADDRESS + core_v_mini_mcu_pkg_SPI2_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_SPI2_IDX = 32'd4;
	localparam [479:0] core_v_mini_mcu_pkg_PERIPHERALS_ADDR_RULES = {core_v_mini_mcu_pkg_RV_PLIC_IDX, core_v_mini_mcu_pkg_RV_PLIC_START_ADDRESS, core_v_mini_mcu_pkg_RV_PLIC_END_ADDRESS, core_v_mini_mcu_pkg_GPIO_IDX, core_v_mini_mcu_pkg_GPIO_START_ADDRESS, core_v_mini_mcu_pkg_GPIO_END_ADDRESS, core_v_mini_mcu_pkg_I2C_IDX, core_v_mini_mcu_pkg_I2C_START_ADDRESS, core_v_mini_mcu_pkg_I2C_END_ADDRESS, core_v_mini_mcu_pkg_RV_TIMER_IDX, core_v_mini_mcu_pkg_RV_TIMER_START_ADDRESS, core_v_mini_mcu_pkg_RV_TIMER_END_ADDRESS, core_v_mini_mcu_pkg_SPI2_IDX, core_v_mini_mcu_pkg_SPI2_START_ADDRESS, core_v_mini_mcu_pkg_SPI2_END_ADDRESS};
	localparam [31:0] sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_NoIndices = core_v_mini_mcu_pkg_PERIPHERALS;
	function automatic [31:0] sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_cf_math_pkg_idx_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:58:9
		sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	localparam [31:0] sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_IdxWidth = sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_cf_math_pkg_idx_width(sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_NoIndices);
	// removed localparam type sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_idx_t
	// removed localparam type sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_default_idx_i
	localparam [sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_IdxWidth - 1:0] sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_ext_default_idx_i_0 = 1'sb0;
	addr_decode_6EF7A #(
		.NoIndices(core_v_mini_mcu_pkg_PERIPHERALS),
		.NoRules(core_v_mini_mcu_pkg_PERIPHERALS)
	) i_addr_decode_soc_regbus_periph_xbar(
		.addr_i(peripheral_req[63-:32]),
		.addr_map_i(core_v_mini_mcu_pkg_PERIPHERALS_ADDR_RULES),
		.idx_o(peripheral_select),
		.dec_valid_o(),
		.dec_error_o(),
		.en_default_idx_i(1'b0),
		.default_idx_i(sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_ext_default_idx_i_0)
	);
	// Trace: design.sv:105448:3
	reg_demux_64ED6 #(.NoPorts(core_v_mini_mcu_pkg_PERIPHERALS)) reg_demux_i(
		.clk_i(clk_cg),
		.rst_ni(rst_ni),
		.in_select_i(peripheral_select),
		.in_req_i(peripheral_req),
		.in_rsp_o(peripheral_rsp),
		.out_req_o(peripheral_slv_req),
		.out_rsp_i(peripheral_slv_rsp)
	);
	// Trace: design.sv:105462:3
	function automatic [6:0] sv2v_cast_4967F;
		input reg [6:0] inp;
		sv2v_cast_4967F = inp;
	endfunction
	function automatic [6:0] sv2v_cast_66F0D;
		input reg [6:0] inp;
		sv2v_cast_66F0D = inp;
	endfunction
	localparam [20:0] tlul_pkg_TL_A_USER_DEFAULT = {7'b0000010, sv2v_cast_4967F(1'sb0), sv2v_cast_66F0D(1'sb0)};
	reg_to_tlul_223C2_EF763 #(
		.tl_a_user_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_a_user_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_d2h_t_tlul_pkg_D2HRspIntgWidth(tlul_pkg_D2HRspIntgWidth),
		.tl_d2h_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_d2h_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_d2h_t_top_pkg_TL_DIW(top_pkg_TL_DIW),
		.tl_d2h_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_d2h_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.tl_h2d_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_h2d_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_h2d_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_h2d_t_top_pkg_TL_AW(top_pkg_TL_AW),
		.tl_h2d_t_top_pkg_TL_DBW(top_pkg_TL_DBW),
		.tl_h2d_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_h2d_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.TL_A_USER_DEFAULT(tlul_pkg_TL_A_USER_DEFAULT),
		.PutFullData(3'h0),
		.Get(3'h4)
	) reg_to_tlul_plic_i(
		.tl_o(plic_tl_h2d),
		.tl_i(plic_tl_d2h),
		.reg_req_i(peripheral_slv_req[0+:70]),
		.reg_rsp_o(peripheral_slv_rsp[0+:34])
	);
	// Trace: design.sv:105479:3
	rv_plic rv_plic_i(
		.clk_i(clk_cg),
		.rst_ni(rst_ni),
		.tl_i(plic_tl_h2d),
		.tl_o(plic_tl_d2h),
		.intr_src_i(intr_vector),
		.irq_o(irq_plic_o),
		.irq_id_o(irq_id),
		.msip_o(msip_o)
	);
	// Trace: design.sv:105491:3
	gpio_B7E66 gpio_i(
		.clk_i(clk_cg),
		.rst_ni(rst_ni),
		.reg_req_i(peripheral_slv_req[70+:70]),
		.reg_rsp_o(peripheral_slv_rsp[34+:34]),
		.gpio_in({cio_gpio_i, 8'b00000000}),
		.gpio_out({cio_gpio_o, cio_gpio_unused}),
		.gpio_tx_en_o({cio_gpio_en_o, cio_gpio_en_unused}),
		.gpio_in_sync_o(),
		.pin_level_interrupts_o({gpio_intr, gpio_int_unused}),
		.global_interrupt_o()
	);
	// Trace: design.sv:105507:3
	reg_to_tlul_223C2_EF763 #(
		.tl_a_user_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_a_user_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_d2h_t_tlul_pkg_D2HRspIntgWidth(tlul_pkg_D2HRspIntgWidth),
		.tl_d2h_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_d2h_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_d2h_t_top_pkg_TL_DIW(top_pkg_TL_DIW),
		.tl_d2h_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_d2h_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.tl_h2d_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_h2d_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_h2d_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_h2d_t_top_pkg_TL_AW(top_pkg_TL_AW),
		.tl_h2d_t_top_pkg_TL_DBW(top_pkg_TL_DBW),
		.tl_h2d_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_h2d_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.TL_A_USER_DEFAULT(tlul_pkg_TL_A_USER_DEFAULT),
		.PutFullData(3'h0),
		.Get(3'h4)
	) reg_to_tlul_i2c_i(
		.tl_o(i2c_tl_h2d),
		.tl_i(i2c_tl_d2h),
		.reg_req_i(peripheral_slv_req[140+:70]),
		.reg_rsp_o(peripheral_slv_rsp[68+:34])
	);
	// Trace: design.sv:105524:3
	// removed localparam type spi_device_pkg_passthrough_req_t
	localparam [13:0] spi_device_pkg_PASSTHROUGH_REQ_DEFAULT = 14'h0200;
	spi_host_CA356 spi2_host(
		.clk_i(clk_cg),
		.rst_ni(rst_ni),
		.reg_req_i(peripheral_slv_req[280+:70]),
		.reg_rsp_o(peripheral_slv_rsp[136+:34]),
		.alert_rx_i(),
		.alert_tx_o(),
		.passthrough_i(spi_device_pkg_PASSTHROUGH_REQ_DEFAULT),
		.passthrough_o(),
		.cio_sck_o(spi2_sck_o),
		.cio_sck_en_o(spi2_sck_en_o),
		.cio_csb_o(spi2_csb_o),
		.cio_csb_en_o(spi2_csb_en_o),
		.cio_sd_o(spi2_sd_o),
		.cio_sd_en_o(spi2_sd_en_o),
		.cio_sd_i(spi2_sd_i),
		.rx_valid_o(),
		.tx_ready_o(),
		.intr_error_o(),
		.intr_spi_event_o(spi2_intr_event)
	);
	// Trace: design.sv:105550:3
	i2c i2c_i(
		.clk_i(clk_cg),
		.rst_ni(rst_ni),
		.tl_i(i2c_tl_h2d),
		.tl_o(i2c_tl_d2h),
		.cio_scl_i(cio_scl_i),
		.cio_scl_o(cio_scl_o),
		.cio_scl_en_o(cio_scl_en_o),
		.cio_sda_i(cio_sda_i),
		.cio_sda_o(cio_sda_o),
		.cio_sda_en_o(cio_sda_en_o),
		.intr_fmt_watermark_o(i2c_intr_fmt_watermark),
		.intr_rx_watermark_o(i2c_intr_rx_watermark),
		.intr_fmt_overflow_o(i2c_intr_fmt_overflow),
		.intr_rx_overflow_o(i2c_intr_rx_overflow),
		.intr_nak_o(i2c_intr_nak),
		.intr_scl_interference_o(i2c_intr_scl_interference),
		.intr_sda_interference_o(i2c_intr_sda_interference),
		.intr_stretch_timeout_o(i2c_intr_stretch_timeout),
		.intr_sda_unstable_o(i2c_intr_sda_unstable),
		.intr_trans_complete_o(i2c_intr_trans_complete),
		.intr_tx_empty_o(i2c_intr_tx_empty),
		.intr_tx_nonempty_o(i2c_intr_tx_nonempty),
		.intr_tx_overflow_o(i2c_intr_tx_overflow),
		.intr_acq_overflow_o(i2c_intr_acq_overflow),
		.intr_ack_stop_o(i2c_intr_ack_stop),
		.intr_host_timeout_o(i2c_intr_host_timeout)
	);
	// Trace: design.sv:105579:3
	reg_to_tlul_223C2_EF763 #(
		.tl_a_user_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_a_user_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_d2h_t_tlul_pkg_D2HRspIntgWidth(tlul_pkg_D2HRspIntgWidth),
		.tl_d2h_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_d2h_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_d2h_t_top_pkg_TL_DIW(top_pkg_TL_DIW),
		.tl_d2h_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_d2h_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.tl_h2d_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_h2d_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_h2d_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_h2d_t_top_pkg_TL_AW(top_pkg_TL_AW),
		.tl_h2d_t_top_pkg_TL_DBW(top_pkg_TL_DBW),
		.tl_h2d_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_h2d_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.TL_A_USER_DEFAULT(tlul_pkg_TL_A_USER_DEFAULT),
		.PutFullData(3'h0),
		.Get(3'h4)
	) rv_timer_reg_to_tlul_i(
		.tl_o(rv_timer_tl_h2d),
		.tl_i(rv_timer_tl_d2h),
		.reg_req_i(peripheral_slv_req[210+:70]),
		.reg_rsp_o(peripheral_slv_rsp[102+:34])
	);
	// Trace: design.sv:105596:3
	rv_timer rv_timer_2_3_i(
		.clk_i(clk_cg),
		.rst_ni(rst_ni),
		.tl_i(rv_timer_tl_h2d),
		.tl_o(rv_timer_tl_d2h),
		.intr_timer_expired_0_0_o(rv_timer_2_intr_o),
		.intr_timer_expired_1_0_o(rv_timer_3_intr_o)
	);
endmodule
module ao_peripheral_subsystem (
	clk_i,
	rst_ni,
	slave_req_i,
	slave_resp_o,
	boot_select_i,
	execute_from_flash_i,
	exit_valid_o,
	exit_value_o,
	spimemio_req_i,
	spimemio_resp_o,
	spi_flash_sck_o,
	spi_flash_sck_en_o,
	spi_flash_csb_o,
	spi_flash_csb_en_o,
	spi_flash_sd_o,
	spi_flash_sd_en_o,
	spi_flash_sd_i,
	spi_sck_o,
	spi_sck_en_o,
	spi_csb_o,
	spi_csb_en_o,
	spi_sd_o,
	spi_sd_en_o,
	spi_sd_i,
	spi_intr_event_o,
	spi_flash_intr_event_o,
	intr_i,
	intr_vector_ext_i,
	core_sleep_i,
	cpu_subsystem_powergate_switch_o,
	cpu_subsystem_powergate_switch_ack_i,
	cpu_subsystem_powergate_iso_o,
	cpu_subsystem_rst_no,
	peripheral_subsystem_powergate_switch_o,
	peripheral_subsystem_powergate_switch_ack_i,
	peripheral_subsystem_powergate_iso_o,
	peripheral_subsystem_rst_no,
	memory_subsystem_banks_powergate_switch_o,
	memory_subsystem_banks_powergate_switch_ack_i,
	memory_subsystem_banks_powergate_iso_o,
	memory_subsystem_banks_set_retentive_o,
	external_subsystem_powergate_switch_o,
	external_subsystem_powergate_switch_ack_i,
	external_subsystem_powergate_iso_o,
	external_subsystem_rst_no,
	external_ram_banks_set_retentive_o,
	peripheral_subsystem_clkgate_en_o,
	memory_subsystem_clkgate_en_o,
	rv_timer_0_intr_o,
	rv_timer_1_intr_o,
	dma_master0_ch0_req_o,
	dma_master0_ch0_resp_i,
	dma_master1_ch0_req_o,
	dma_master1_ch0_resp_i,
	dma_intr_o,
	pad_req_o,
	pad_resp_i,
	fast_intr_i,
	fast_intr_o,
	cio_gpio_i,
	cio_gpio_o,
	cio_gpio_en_o,
	intr_gpio_o,
	uart_rx_i,
	uart_tx_o,
	uart_intr_tx_watermark_o,
	uart_intr_rx_watermark_o,
	uart_intr_tx_empty_o,
	uart_intr_rx_overflow_o,
	uart_intr_rx_frame_err_o,
	uart_intr_rx_break_err_o,
	uart_intr_rx_timeout_o,
	uart_intr_rx_parity_err_o,
	ext_peripheral_slave_req_o,
	ext_peripheral_slave_resp_i
);
	// removed import obi_pkg::*;
	// removed import reg_pkg::*;
	// Trace: design.sv:105614:5
	input wire clk_i;
	// Trace: design.sv:105615:5
	input wire rst_ni;
	// Trace: design.sv:105617:5
	// removed localparam type obi_pkg_obi_req_t
	input wire [69:0] slave_req_i;
	// Trace: design.sv:105618:5
	// removed localparam type obi_pkg_obi_resp_t
	output wire [33:0] slave_resp_o;
	// Trace: design.sv:105621:5
	input wire boot_select_i;
	// Trace: design.sv:105622:5
	input wire execute_from_flash_i;
	// Trace: design.sv:105623:5
	output wire exit_valid_o;
	// Trace: design.sv:105624:5
	output wire [31:0] exit_value_o;
	// Trace: design.sv:105627:5
	input wire [69:0] spimemio_req_i;
	// Trace: design.sv:105628:5
	output wire [33:0] spimemio_resp_o;
	// Trace: design.sv:105631:5
	output wire spi_flash_sck_o;
	// Trace: design.sv:105632:5
	output wire spi_flash_sck_en_o;
	// Trace: design.sv:105633:5
	localparam signed [31:0] spi_host_reg_pkg_NumCS = 2;
	output wire [1:0] spi_flash_csb_o;
	// Trace: design.sv:105634:5
	output wire [1:0] spi_flash_csb_en_o;
	// Trace: design.sv:105635:5
	output wire [3:0] spi_flash_sd_o;
	// Trace: design.sv:105636:5
	output wire [3:0] spi_flash_sd_en_o;
	// Trace: design.sv:105637:5
	input wire [3:0] spi_flash_sd_i;
	// Trace: design.sv:105640:5
	output wire spi_sck_o;
	// Trace: design.sv:105641:5
	output wire spi_sck_en_o;
	// Trace: design.sv:105642:5
	output wire [1:0] spi_csb_o;
	// Trace: design.sv:105643:5
	output wire [1:0] spi_csb_en_o;
	// Trace: design.sv:105644:5
	output wire [3:0] spi_sd_o;
	// Trace: design.sv:105645:5
	output wire [3:0] spi_sd_en_o;
	// Trace: design.sv:105646:5
	input wire [3:0] spi_sd_i;
	// Trace: design.sv:105647:5
	output wire spi_intr_event_o;
	// Trace: design.sv:105648:5
	output wire spi_flash_intr_event_o;
	// Trace: design.sv:105651:5
	input wire [31:0] intr_i;
	// Trace: design.sv:105652:5
	localparam core_v_mini_mcu_pkg_PLIC_NINT = 64;
	localparam core_v_mini_mcu_pkg_PLIC_USED_NINT = 50;
	localparam core_v_mini_mcu_pkg_NEXT_INT = 14;
	input wire [13:0] intr_vector_ext_i;
	// Trace: design.sv:105653:5
	input wire core_sleep_i;
	// Trace: design.sv:105654:5
	output wire cpu_subsystem_powergate_switch_o;
	// Trace: design.sv:105655:5
	input wire cpu_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:105656:5
	output wire cpu_subsystem_powergate_iso_o;
	// Trace: design.sv:105657:5
	output wire cpu_subsystem_rst_no;
	// Trace: design.sv:105658:5
	output wire peripheral_subsystem_powergate_switch_o;
	// Trace: design.sv:105659:5
	input wire peripheral_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:105660:5
	output wire peripheral_subsystem_powergate_iso_o;
	// Trace: design.sv:105661:5
	output wire peripheral_subsystem_rst_no;
	// Trace: design.sv:105662:5
	localparam [31:0] core_v_mini_mcu_pkg_NUM_BANKS = 2;
	output wire [1:0] memory_subsystem_banks_powergate_switch_o;
	// Trace: design.sv:105663:5
	input wire [1:0] memory_subsystem_banks_powergate_switch_ack_i;
	// Trace: design.sv:105664:5
	output wire [1:0] memory_subsystem_banks_powergate_iso_o;
	// Trace: design.sv:105665:5
	output wire [1:0] memory_subsystem_banks_set_retentive_o;
	// Trace: design.sv:105666:5
	localparam [31:0] core_v_mini_mcu_pkg_EXTERNAL_DOMAINS = 0;
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_switch_o;
	// Trace: design.sv:105667:5
	input wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_switch_ack_i;
	// Trace: design.sv:105668:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_powergate_iso_o;
	// Trace: design.sv:105669:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_subsystem_rst_no;
	// Trace: design.sv:105670:5
	output wire [core_v_mini_mcu_pkg_EXTERNAL_DOMAINS - 1:0] external_ram_banks_set_retentive_o;
	// Trace: design.sv:105673:5
	output wire peripheral_subsystem_clkgate_en_o;
	// Trace: design.sv:105674:5
	output wire [1:0] memory_subsystem_clkgate_en_o;
	// Trace: design.sv:105677:5
	output wire rv_timer_0_intr_o;
	// Trace: design.sv:105678:5
	output wire rv_timer_1_intr_o;
	// Trace: design.sv:105681:5
	output wire [69:0] dma_master0_ch0_req_o;
	// Trace: design.sv:105682:5
	input wire [33:0] dma_master0_ch0_resp_i;
	// Trace: design.sv:105683:5
	output wire [69:0] dma_master1_ch0_req_o;
	// Trace: design.sv:105684:5
	input wire [33:0] dma_master1_ch0_resp_i;
	// Trace: design.sv:105685:5
	output wire dma_intr_o;
	// Trace: design.sv:105688:5
	// removed localparam type reg_pkg_reg_req_t
	output wire [69:0] pad_req_o;
	// Trace: design.sv:105689:5
	// removed localparam type reg_pkg_reg_rsp_t
	input wire [33:0] pad_resp_i;
	// Trace: design.sv:105692:5
	input wire [14:0] fast_intr_i;
	// Trace: design.sv:105693:5
	output wire [14:0] fast_intr_o;
	// Trace: design.sv:105696:5
	input wire [7:0] cio_gpio_i;
	// Trace: design.sv:105697:5
	output wire [7:0] cio_gpio_o;
	// Trace: design.sv:105698:5
	output wire [7:0] cio_gpio_en_o;
	// Trace: design.sv:105699:5
	output wire [7:0] intr_gpio_o;
	// Trace: design.sv:105702:5
	input wire uart_rx_i;
	// Trace: design.sv:105703:5
	output wire uart_tx_o;
	// Trace: design.sv:105704:5
	output wire uart_intr_tx_watermark_o;
	// Trace: design.sv:105705:5
	output wire uart_intr_rx_watermark_o;
	// Trace: design.sv:105706:5
	output wire uart_intr_tx_empty_o;
	// Trace: design.sv:105707:5
	output wire uart_intr_rx_overflow_o;
	// Trace: design.sv:105708:5
	output wire uart_intr_rx_frame_err_o;
	// Trace: design.sv:105709:5
	output wire uart_intr_rx_break_err_o;
	// Trace: design.sv:105710:5
	output wire uart_intr_rx_timeout_o;
	// Trace: design.sv:105711:5
	output wire uart_intr_rx_parity_err_o;
	// Trace: design.sv:105714:5
	output wire [69:0] ext_peripheral_slave_req_o;
	// Trace: design.sv:105715:5
	input wire [33:0] ext_peripheral_slave_resp_i;
	// Trace: design.sv:105718:3
	// removed import core_v_mini_mcu_pkg::*;
	// Trace: design.sv:105719:3
	// removed import tlul_pkg::*;
	// Trace: design.sv:105720:3
	// removed import rv_plic_reg_pkg::*;
	// Trace: design.sv:105722:3
	wire [69:0] peripheral_req;
	// Trace: design.sv:105723:3
	wire [33:0] peripheral_rsp;
	// Trace: design.sv:105725:3
	localparam core_v_mini_mcu_pkg_AO_PERIPHERALS = 13;
	wire [909:0] ao_peripheral_slv_req;
	// Trace: design.sv:105726:3
	wire [441:0] ao_peripheral_slv_rsp;
	// Trace: design.sv:105728:3
	// removed localparam type tlul_pkg_tl_a_op_e
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_type_e
	// removed localparam type tlul_pkg_tl_a_user_t
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	// removed localparam type tlul_pkg_tl_h2d_t
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] rv_timer_tl_h2d;
	// Trace: design.sv:105729:3
	// removed localparam type tlul_pkg_tl_d_op_e
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	// removed localparam type tlul_pkg_tl_d_user_t
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	// removed localparam type tlul_pkg_tl_d2h_t
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] rv_timer_tl_d2h;
	// Trace: design.sv:105731:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 21:0] uart_tl_h2d;
	// Trace: design.sv:105732:3
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] uart_tl_d2h;
	// Trace: design.sv:105734:3
	localparam [31:0] core_v_mini_mcu_pkg_AO_PERIPHERALS_PORT_SEL_WIDTH = 4;
	wire [3:0] peripheral_select;
	// Trace: design.sv:105736:3
	wire use_spimemio;
	// Trace: design.sv:105738:3
	wire spi_rx_valid;
	// Trace: design.sv:105739:3
	wire spi_tx_ready;
	// Trace: design.sv:105740:3
	wire spi_flash_rx_valid;
	// Trace: design.sv:105741:3
	wire spi_flash_tx_ready;
	// Trace: design.sv:105743:3
	wire [23:0] intr_gpio_unused;
	// Trace: design.sv:105744:3
	wire [23:0] cio_gpio_unused;
	// Trace: design.sv:105745:3
	wire [23:0] cio_gpio_en_unused;
	// Trace: design.sv:105747:3
	localparam [31:0] core_v_mini_mcu_pkg_EXT_PERIPHERAL_IDX = 32'd9;
	assign ext_peripheral_slave_req_o = ao_peripheral_slv_req[630+:70];
	// Trace: design.sv:105748:3
	assign ao_peripheral_slv_rsp[306+:34] = ext_peripheral_slave_resp_i;
	// Trace: design.sv:105750:3
	localparam [31:0] sv2v_uu_periph_to_reg_i_IW = 1;
	// removed localparam type sv2v_uu_periph_to_reg_i_id_i
	localparam [0:0] sv2v_uu_periph_to_reg_i_ext_id_i_0 = 1'sb0;
	periph_to_reg_35129 #(.IW(1)) periph_to_reg_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.req_i(slave_req_i[69]),
		.add_i(slave_req_i[63-:32]),
		.wen_i(~slave_req_i[68]),
		.wdata_i(slave_req_i[31-:32]),
		.be_i(slave_req_i[67-:4]),
		.id_i(sv2v_uu_periph_to_reg_i_ext_id_i_0),
		.gnt_o(slave_resp_o[33]),
		.r_rdata_o(slave_resp_o[31-:32]),
		.r_opc_o(),
		.r_id_o(),
		.r_valid_o(slave_resp_o[32]),
		.reg_req_o(peripheral_req),
		.reg_rsp_i(peripheral_rsp)
	);
	// Trace: design.sv:105772:3
	// removed localparam type addr_map_rule_pkg_addr_map_rule_t
	localparam [31:0] core_v_mini_mcu_pkg_BOOTROM_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS = 32'h20000000;
	localparam [31:0] core_v_mini_mcu_pkg_BOOTROM_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_BOOTROM_END_ADDRESS = core_v_mini_mcu_pkg_BOOTROM_START_ADDRESS + core_v_mini_mcu_pkg_BOOTROM_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_BOOTROM_IDX = 32'd1;
	localparam [31:0] core_v_mini_mcu_pkg_DMA_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_DMA_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00060000;
	localparam [31:0] core_v_mini_mcu_pkg_DMA_END_ADDRESS = core_v_mini_mcu_pkg_DMA_START_ADDRESS + core_v_mini_mcu_pkg_DMA_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_DMA_IDX = 32'd7;
	localparam [31:0] core_v_mini_mcu_pkg_EXT_PERIPHERAL_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_EXT_PERIPHERAL_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00080000;
	localparam [31:0] core_v_mini_mcu_pkg_EXT_PERIPHERAL_END_ADDRESS = core_v_mini_mcu_pkg_EXT_PERIPHERAL_START_ADDRESS + core_v_mini_mcu_pkg_EXT_PERIPHERAL_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_FAST_INTR_CTRL_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_FAST_INTR_CTRL_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00070000;
	localparam [31:0] core_v_mini_mcu_pkg_FAST_INTR_CTRL_END_ADDRESS = core_v_mini_mcu_pkg_FAST_INTR_CTRL_START_ADDRESS + core_v_mini_mcu_pkg_FAST_INTR_CTRL_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_FAST_INTR_CTRL_IDX = 32'd8;
	localparam [31:0] core_v_mini_mcu_pkg_GPIO_AO_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_GPIO_AO_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h000a0000;
	localparam [31:0] core_v_mini_mcu_pkg_GPIO_AO_END_ADDRESS = core_v_mini_mcu_pkg_GPIO_AO_START_ADDRESS + core_v_mini_mcu_pkg_GPIO_AO_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_GPIO_AO_IDX = 32'd11;
	localparam [31:0] core_v_mini_mcu_pkg_PAD_CONTROL_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_PAD_CONTROL_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00090000;
	localparam [31:0] core_v_mini_mcu_pkg_PAD_CONTROL_END_ADDRESS = core_v_mini_mcu_pkg_PAD_CONTROL_START_ADDRESS + core_v_mini_mcu_pkg_PAD_CONTROL_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_PAD_CONTROL_IDX = 32'd10;
	localparam [31:0] core_v_mini_mcu_pkg_POWER_MANAGER_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_POWER_MANAGER_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00040000;
	localparam [31:0] core_v_mini_mcu_pkg_POWER_MANAGER_END_ADDRESS = core_v_mini_mcu_pkg_POWER_MANAGER_START_ADDRESS + core_v_mini_mcu_pkg_POWER_MANAGER_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_POWER_MANAGER_IDX = 32'd5;
	localparam [31:0] core_v_mini_mcu_pkg_RV_TIMER_AO_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_RV_TIMER_AO_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00050000;
	localparam [31:0] core_v_mini_mcu_pkg_RV_TIMER_AO_END_ADDRESS = core_v_mini_mcu_pkg_RV_TIMER_AO_START_ADDRESS + core_v_mini_mcu_pkg_RV_TIMER_AO_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_RV_TIMER_AO_IDX = 32'd6;
	localparam [31:0] core_v_mini_mcu_pkg_SOC_CTRL_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_SOC_CTRL_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00000000;
	localparam [31:0] core_v_mini_mcu_pkg_SOC_CTRL_END_ADDRESS = core_v_mini_mcu_pkg_SOC_CTRL_START_ADDRESS + core_v_mini_mcu_pkg_SOC_CTRL_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_SOC_CTRL_IDX = 32'd0;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_FLASH_SIZE = 32'h00008000;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_FLASH_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00020000;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_FLASH_END_ADDRESS = core_v_mini_mcu_pkg_SPI_FLASH_START_ADDRESS + core_v_mini_mcu_pkg_SPI_FLASH_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_FLASH_IDX = 32'd2;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_HOST_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_HOST_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00030000;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_HOST_END_ADDRESS = core_v_mini_mcu_pkg_SPI_HOST_START_ADDRESS + core_v_mini_mcu_pkg_SPI_HOST_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_HOST_IDX = 32'd4;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_MEMIO_SIZE = 32'h00008000;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_MEMIO_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h00028000;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_MEMIO_END_ADDRESS = core_v_mini_mcu_pkg_SPI_MEMIO_START_ADDRESS + core_v_mini_mcu_pkg_SPI_MEMIO_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_SPI_MEMIO_IDX = 32'd3;
	localparam [31:0] core_v_mini_mcu_pkg_UART_SIZE = 32'h00010000;
	localparam [31:0] core_v_mini_mcu_pkg_UART_START_ADDRESS = core_v_mini_mcu_pkg_AO_PERIPHERAL_START_ADDRESS + 32'h000b0000;
	localparam [31:0] core_v_mini_mcu_pkg_UART_END_ADDRESS = core_v_mini_mcu_pkg_UART_START_ADDRESS + core_v_mini_mcu_pkg_UART_SIZE;
	localparam [31:0] core_v_mini_mcu_pkg_UART_IDX = 32'd12;
	localparam [1247:0] core_v_mini_mcu_pkg_AO_PERIPHERALS_ADDR_RULES = {core_v_mini_mcu_pkg_SOC_CTRL_IDX, core_v_mini_mcu_pkg_SOC_CTRL_START_ADDRESS, core_v_mini_mcu_pkg_SOC_CTRL_END_ADDRESS, core_v_mini_mcu_pkg_BOOTROM_IDX, core_v_mini_mcu_pkg_BOOTROM_START_ADDRESS, core_v_mini_mcu_pkg_BOOTROM_END_ADDRESS, core_v_mini_mcu_pkg_SPI_FLASH_IDX, core_v_mini_mcu_pkg_SPI_FLASH_START_ADDRESS, core_v_mini_mcu_pkg_SPI_FLASH_END_ADDRESS, core_v_mini_mcu_pkg_SPI_MEMIO_IDX, core_v_mini_mcu_pkg_SPI_MEMIO_START_ADDRESS, core_v_mini_mcu_pkg_SPI_MEMIO_END_ADDRESS, core_v_mini_mcu_pkg_SPI_HOST_IDX, core_v_mini_mcu_pkg_SPI_HOST_START_ADDRESS, core_v_mini_mcu_pkg_SPI_HOST_END_ADDRESS, core_v_mini_mcu_pkg_POWER_MANAGER_IDX, core_v_mini_mcu_pkg_POWER_MANAGER_START_ADDRESS, core_v_mini_mcu_pkg_POWER_MANAGER_END_ADDRESS, core_v_mini_mcu_pkg_RV_TIMER_AO_IDX, core_v_mini_mcu_pkg_RV_TIMER_AO_START_ADDRESS, core_v_mini_mcu_pkg_RV_TIMER_AO_END_ADDRESS, core_v_mini_mcu_pkg_DMA_IDX, core_v_mini_mcu_pkg_DMA_START_ADDRESS, core_v_mini_mcu_pkg_DMA_END_ADDRESS, core_v_mini_mcu_pkg_FAST_INTR_CTRL_IDX, core_v_mini_mcu_pkg_FAST_INTR_CTRL_START_ADDRESS, core_v_mini_mcu_pkg_FAST_INTR_CTRL_END_ADDRESS, core_v_mini_mcu_pkg_EXT_PERIPHERAL_IDX, core_v_mini_mcu_pkg_EXT_PERIPHERAL_START_ADDRESS, core_v_mini_mcu_pkg_EXT_PERIPHERAL_END_ADDRESS, core_v_mini_mcu_pkg_PAD_CONTROL_IDX, core_v_mini_mcu_pkg_PAD_CONTROL_START_ADDRESS, core_v_mini_mcu_pkg_PAD_CONTROL_END_ADDRESS, core_v_mini_mcu_pkg_GPIO_AO_IDX, core_v_mini_mcu_pkg_GPIO_AO_START_ADDRESS, core_v_mini_mcu_pkg_GPIO_AO_END_ADDRESS, core_v_mini_mcu_pkg_UART_IDX, core_v_mini_mcu_pkg_UART_START_ADDRESS, core_v_mini_mcu_pkg_UART_END_ADDRESS};
	localparam [31:0] sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_NoIndices = core_v_mini_mcu_pkg_AO_PERIPHERALS;
	function automatic [31:0] sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_cf_math_pkg_idx_width;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: ../src/pulp-platform.org__common_cells_1.28.0/src/cf_math_pkg.sv:58:9
		sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	localparam [31:0] sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_IdxWidth = sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_cf_math_pkg_idx_width(sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_NoIndices);
	// removed localparam type sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_idx_t
	// removed localparam type sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_default_idx_i
	localparam [sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_IdxWidth - 1:0] sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_ext_default_idx_i_0 = 1'sb0;
	addr_decode_6EF7A #(
		.NoIndices(core_v_mini_mcu_pkg_AO_PERIPHERALS),
		.NoRules(core_v_mini_mcu_pkg_AO_PERIPHERALS)
	) i_addr_decode_soc_regbus_periph_xbar(
		.addr_i(peripheral_req[63-:32]),
		.addr_map_i(core_v_mini_mcu_pkg_AO_PERIPHERALS_ADDR_RULES),
		.idx_o(peripheral_select),
		.dec_valid_o(),
		.dec_error_o(),
		.en_default_idx_i(1'b0),
		.default_idx_i(sv2v_uu_i_addr_decode_soc_regbus_periph_xbar_ext_default_idx_i_0)
	);
	// Trace: design.sv:105787:3
	reg_demux_64ED6 #(.NoPorts(core_v_mini_mcu_pkg_AO_PERIPHERALS)) reg_demux_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.in_select_i(peripheral_select),
		.in_req_i(peripheral_req),
		.in_rsp_o(peripheral_rsp),
		.out_req_o(ao_peripheral_slv_req),
		.out_rsp_i(ao_peripheral_slv_rsp)
	);
	// Trace: design.sv:105801:3
	soc_ctrl_E136A soc_ctrl_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(ao_peripheral_slv_req[0+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[0+:34]),
		.boot_select_i(boot_select_i),
		.execute_from_flash_i(execute_from_flash_i),
		.use_spimemio_o(use_spimemio),
		.exit_valid_o(exit_valid_o),
		.exit_value_o(exit_value_o)
	);
	// Trace: design.sv:105816:3
	boot_rom boot_rom_i(
		.reg_req_i(ao_peripheral_slv_req[70+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[34+:34])
	);
	// Trace: design.sv:105821:3
	spi_subsystem spi_subsystem_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.use_spimemio_i(use_spimemio),
		.spimemio_req_i(spimemio_req_i),
		.spimemio_resp_o(spimemio_resp_o),
		.yo_reg_req_i(ao_peripheral_slv_req[210+:70]),
		.yo_reg_rsp_o(ao_peripheral_slv_rsp[102+:34]),
		.ot_reg_req_i(ao_peripheral_slv_req[140+:70]),
		.ot_reg_rsp_o(ao_peripheral_slv_rsp[68+:34]),
		.spi_flash_sck_o(spi_flash_sck_o),
		.spi_flash_sck_en_o(spi_flash_sck_en_o),
		.spi_flash_csb_o(spi_flash_csb_o),
		.spi_flash_csb_en_o(spi_flash_csb_en_o),
		.spi_flash_sd_o(spi_flash_sd_o),
		.spi_flash_sd_en_o(spi_flash_sd_en_o),
		.spi_flash_sd_i(spi_flash_sd_i),
		.spi_flash_intr_error_o(),
		.spi_flash_intr_event_o(spi_flash_intr_event_o),
		.spi_flash_rx_valid_o(spi_flash_rx_valid),
		.spi_flash_tx_ready_o(spi_flash_tx_ready)
	);
	// Trace: design.sv:105844:3
	// removed localparam type spi_device_pkg_passthrough_req_t
	localparam [13:0] spi_device_pkg_PASSTHROUGH_REQ_DEFAULT = 14'h0200;
	spi_host_CA356 spi_host_dma_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(ao_peripheral_slv_req[280+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[136+:34]),
		.alert_rx_i(),
		.alert_tx_o(),
		.passthrough_i(spi_device_pkg_PASSTHROUGH_REQ_DEFAULT),
		.passthrough_o(),
		.cio_sck_o(spi_sck_o),
		.cio_sck_en_o(spi_sck_en_o),
		.cio_csb_o(spi_csb_o),
		.cio_csb_en_o(spi_csb_en_o),
		.cio_sd_o(spi_sd_o),
		.cio_sd_en_o(spi_sd_en_o),
		.cio_sd_i(spi_sd_i),
		.rx_valid_o(spi_rx_valid),
		.tx_ready_o(spi_tx_ready),
		.intr_error_o(),
		.intr_spi_event_o(spi_intr_event_o)
	);
	// Trace: design.sv:105869:3
	power_manager_2EE6F power_manager_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(ao_peripheral_slv_req[350+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[170+:34]),
		.intr_i(intr_i),
		.ext_irq_i(intr_vector_ext_i),
		.core_sleep_i(core_sleep_i),
		.cpu_subsystem_powergate_switch_o(cpu_subsystem_powergate_switch_o),
		.cpu_subsystem_powergate_switch_ack_i(cpu_subsystem_powergate_switch_ack_i),
		.cpu_subsystem_powergate_iso_o(cpu_subsystem_powergate_iso_o),
		.cpu_subsystem_rst_no(cpu_subsystem_rst_no),
		.peripheral_subsystem_powergate_switch_o(peripheral_subsystem_powergate_switch_o),
		.peripheral_subsystem_powergate_switch_ack_i(peripheral_subsystem_powergate_switch_ack_i),
		.peripheral_subsystem_powergate_iso_o(peripheral_subsystem_powergate_iso_o),
		.peripheral_subsystem_rst_no(peripheral_subsystem_rst_no),
		.memory_subsystem_banks_powergate_switch_o(memory_subsystem_banks_powergate_switch_o),
		.memory_subsystem_banks_powergate_switch_ack_i(memory_subsystem_banks_powergate_switch_ack_i),
		.memory_subsystem_banks_powergate_iso_o(memory_subsystem_banks_powergate_iso_o),
		.memory_subsystem_banks_set_retentive_o(memory_subsystem_banks_set_retentive_o),
		.external_subsystem_powergate_switch_o(external_subsystem_powergate_switch_o),
		.external_subsystem_powergate_switch_ack_i(external_subsystem_powergate_switch_ack_i),
		.external_subsystem_powergate_iso_o(external_subsystem_powergate_iso_o),
		.external_subsystem_rst_no(external_subsystem_rst_no),
		.external_ram_banks_set_retentive_o(external_ram_banks_set_retentive_o),
		.peripheral_subsystem_clkgate_en_o(peripheral_subsystem_clkgate_en_o),
		.memory_subsystem_clkgate_en_o(memory_subsystem_clkgate_en_o)
	);
	// Trace: design.sv:105901:3
	function automatic [6:0] sv2v_cast_65793;
		input reg [6:0] inp;
		sv2v_cast_65793 = inp;
	endfunction
	function automatic [6:0] sv2v_cast_F1979;
		input reg [6:0] inp;
		sv2v_cast_F1979 = inp;
	endfunction
	localparam [20:0] tlul_pkg_TL_A_USER_DEFAULT = {7'b0000010, sv2v_cast_65793(1'sb0), sv2v_cast_F1979(1'sb0)};
	reg_to_tlul_223C2_EF763 #(
		.tl_a_user_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_a_user_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_d2h_t_tlul_pkg_D2HRspIntgWidth(tlul_pkg_D2HRspIntgWidth),
		.tl_d2h_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_d2h_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_d2h_t_top_pkg_TL_DIW(top_pkg_TL_DIW),
		.tl_d2h_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_d2h_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.tl_h2d_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_h2d_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_h2d_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_h2d_t_top_pkg_TL_AW(top_pkg_TL_AW),
		.tl_h2d_t_top_pkg_TL_DBW(top_pkg_TL_DBW),
		.tl_h2d_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_h2d_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.TL_A_USER_DEFAULT(tlul_pkg_TL_A_USER_DEFAULT),
		.PutFullData(3'h0),
		.Get(3'h4)
	) rv_timer_reg_to_tlul_i(
		.tl_o(rv_timer_tl_h2d),
		.tl_i(rv_timer_tl_d2h),
		.reg_req_i(ao_peripheral_slv_req[420+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[204+:34])
	);
	// Trace: design.sv:105918:3
	rv_timer rv_timer_0_1_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(rv_timer_tl_h2d),
		.tl_o(rv_timer_tl_d2h),
		.intr_timer_expired_0_0_o(rv_timer_0_intr_o),
		.intr_timer_expired_1_0_o(rv_timer_1_intr_o)
	);
	// Trace: design.sv:105927:3
	dma_689DF dma_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(ao_peripheral_slv_req[490+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[238+:34]),
		.dma_master0_ch0_req_o(dma_master0_ch0_req_o),
		.dma_master0_ch0_resp_i(dma_master0_ch0_resp_i),
		.dma_master1_ch0_req_o(dma_master1_ch0_req_o),
		.dma_master1_ch0_resp_i(dma_master1_ch0_resp_i),
		.spi_rx_valid_i(spi_rx_valid),
		.spi_tx_ready_i(spi_tx_ready),
		.spi_flash_rx_valid_i(spi_flash_rx_valid),
		.spi_flash_tx_ready_i(spi_flash_tx_ready),
		.dma_intr_o(dma_intr_o)
	);
	// Trace: design.sv:105948:3
	assign pad_req_o = ao_peripheral_slv_req[700+:70];
	// Trace: design.sv:105949:3
	assign ao_peripheral_slv_rsp[340+:34] = pad_resp_i;
	// Trace: design.sv:105951:3
	fast_intr_ctrl_65415 fast_intr_ctrl_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(ao_peripheral_slv_req[560+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[272+:34]),
		.fast_intr_i(fast_intr_i),
		.fast_intr_o(fast_intr_o)
	);
	// Trace: design.sv:105963:3
	gpio_B7E66 gpio_ao_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.reg_req_i(ao_peripheral_slv_req[770+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[374+:34]),
		.gpio_in({24'b000000000000000000000000, cio_gpio_i}),
		.gpio_out({cio_gpio_unused, cio_gpio_o}),
		.gpio_tx_en_o({cio_gpio_en_unused, cio_gpio_en_o}),
		.gpio_in_sync_o(),
		.pin_level_interrupts_o({intr_gpio_unused, intr_gpio_o}),
		.global_interrupt_o()
	);
	// Trace: design.sv:105979:3
	reg_to_tlul_223C2_EF763 #(
		.tl_a_user_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_a_user_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_d2h_t_tlul_pkg_D2HRspIntgWidth(tlul_pkg_D2HRspIntgWidth),
		.tl_d2h_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_d2h_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_d2h_t_top_pkg_TL_DIW(top_pkg_TL_DIW),
		.tl_d2h_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_d2h_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.tl_h2d_t_tlul_pkg_DataIntgWidth(tlul_pkg_DataIntgWidth),
		.tl_h2d_t_tlul_pkg_H2DCmdIntgWidth(tlul_pkg_H2DCmdIntgWidth),
		.tl_h2d_t_top_pkg_TL_AIW(top_pkg_TL_AIW),
		.tl_h2d_t_top_pkg_TL_AW(top_pkg_TL_AW),
		.tl_h2d_t_top_pkg_TL_DBW(top_pkg_TL_DBW),
		.tl_h2d_t_top_pkg_TL_DW(top_pkg_TL_DW),
		.tl_h2d_t_top_pkg_TL_SZW(top_pkg_TL_SZW),
		.TL_A_USER_DEFAULT(tlul_pkg_TL_A_USER_DEFAULT),
		.PutFullData(3'h0),
		.Get(3'h4)
	) reg_to_tlul_uart_i(
		.tl_o(uart_tl_h2d),
		.tl_i(uart_tl_d2h),
		.reg_req_i(ao_peripheral_slv_req[840+:70]),
		.reg_rsp_o(ao_peripheral_slv_rsp[408+:34])
	);
	// Trace: design.sv:105996:3
	uart uart_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(uart_tl_h2d),
		.tl_o(uart_tl_d2h),
		.cio_rx_i(uart_rx_i),
		.cio_tx_o(uart_tx_o),
		.cio_tx_en_o(),
		.intr_tx_watermark_o(uart_intr_tx_watermark_o),
		.intr_rx_watermark_o(uart_intr_rx_watermark_o),
		.intr_tx_empty_o(uart_intr_tx_empty_o),
		.intr_rx_overflow_o(uart_intr_rx_overflow_o),
		.intr_rx_frame_err_o(uart_intr_rx_frame_err_o),
		.intr_rx_break_err_o(uart_intr_rx_break_err_o),
		.intr_rx_timeout_o(uart_intr_rx_timeout_o),
		.intr_rx_parity_err_o(uart_intr_rx_parity_err_o)
	);
endmodule
module sram_wrapper (
	clk_i,
	rst_ni,
	req_i,
	we_i,
	addr_i,
	wdata_i,
	be_i,
	set_retentive_i,
	rdata_o
);
	reg _sv2v_0;
	// Trace: design.sv:106021:15
	parameter [31:0] NumWords = 32'd1024;
	// Trace: design.sv:106022:15
	parameter [31:0] DataWidth = 32'd32;
	// Trace: design.sv:106024:15
	parameter [31:0] AddrWidth = (NumWords > 32'd1 ? $clog2(NumWords) : 32'd1);
	// Trace: design.sv:106026:5
	input wire clk_i;
	// Trace: design.sv:106027:5
	input wire rst_ni;
	// Trace: design.sv:106029:5
	input wire req_i;
	// Trace: design.sv:106030:5
	input wire we_i;
	// Trace: design.sv:106031:5
	input wire [AddrWidth - 1:0] addr_i;
	// Trace: design.sv:106032:5
	input wire [31:0] wdata_i;
	// Trace: design.sv:106033:5
	input wire [3:0] be_i;
	// Trace: design.sv:106034:5
	input wire set_retentive_i;
	// Trace: design.sv:106036:5
	output wire [31:0] rdata_o;
	// Trace: design.sv:106039:3
	wire [7:0] unused;
	// Trace: design.sv:106040:3
	reg [7:0] cs;
	// Trace: design.sv:106042:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:106044:5
		cs = 1'sb0;
		// Trace: design.sv:106045:5
		cs[addr_i[AddrWidth - 1:AddrWidth - 3]] = 1'b1;
	end
	// Trace: design.sv:106048:3
	sky130_sram_4kbyte_1rw_32x1024_8 cut0_i(
		.clk0(clk_i),
		.csb0(~cs[0]),
		.web0(~we_i),
		.wmask0(be_i),
		.addr0($unsigned(addr_i[AddrWidth - 4:0])),
		.din0({1'b0, wdata_i}),
		.dout0({unused[0], rdata_o})
	);
	// Trace: design.sv:106067:3
	sky130_sram_4kbyte_1rw_32x1024_8 cut1_i(
		.clk0(clk_i),
		.csb0(~cs[1]),
		.web0(~we_i),
		.wmask0(be_i),
		.addr0($unsigned(addr_i[AddrWidth - 4:0])),
		.din0({1'b0, wdata_i}),
		.dout0({unused[1], rdata_o})
	);
	// Trace: design.sv:106086:3
	sky130_sram_4kbyte_1rw_32x1024_8 cut2_i(
		.clk0(clk_i),
		.csb0(~cs[2]),
		.web0(~we_i),
		.wmask0(be_i),
		.addr0($unsigned(addr_i[AddrWidth - 4:0])),
		.din0({1'b0, wdata_i}),
		.dout0({unused[2], rdata_o})
	);
	// Trace: design.sv:106106:3
	sky130_sram_4kbyte_1rw_32x1024_8 cut3_i(
		.clk0(clk_i),
		.csb0(~cs[3]),
		.web0(~we_i),
		.wmask0(be_i),
		.addr0($unsigned(addr_i[AddrWidth - 4:0])),
		.din0({1'b0, wdata_i}),
		.dout0({unused[3], rdata_o})
	);
	// Trace: design.sv:106125:3
	sky130_sram_4kbyte_1rw_32x1024_8 cut4_i(
		.clk0(clk_i),
		.csb0(~cs[4]),
		.web0(~we_i),
		.wmask0(be_i),
		.addr0($unsigned(addr_i[AddrWidth - 4:0])),
		.din0({1'b0, wdata_i}),
		.dout0({unused[4], rdata_o})
	);
	// Trace: design.sv:106144:3
	sky130_sram_4kbyte_1rw_32x1024_8 cut5_i(
		.clk0(clk_i),
		.csb0(~cs[5]),
		.web0(~we_i),
		.wmask0(be_i),
		.addr0($unsigned(addr_i[AddrWidth - 4:0])),
		.din0({1'b0, wdata_i}),
		.dout0({unused[5], rdata_o})
	);
	// Trace: design.sv:106163:3
	sky130_sram_4kbyte_1rw_32x1024_8 cut6_i(
		.clk0(clk_i),
		.csb0(~cs[6]),
		.web0(~we_i),
		.wmask0(be_i),
		.addr0($unsigned(addr_i[AddrWidth - 4:0])),
		.din0({1'b0, wdata_i}),
		.dout0({unused[6], rdata_o})
	);
	// Trace: design.sv:106182:3
	sky130_sram_4kbyte_1rw_32x1024_8 cut7_i(
		.clk0(clk_i),
		.csb0(~cs[7]),
		.web0(~we_i),
		.wmask0(be_i),
		.addr0($unsigned(addr_i[AddrWidth - 4:0])),
		.din0({1'b0, wdata_i}),
		.dout0({unused[7], rdata_o})
	);
	initial _sv2v_0 = 0;
endmodule
module cve2_clock_gate (
	clk_i,
	en_i,
	scan_cg_en_i,
	clk_o
);
	reg _sv2v_0;
	// Trace: design.sv:106216:5
	input wire clk_i;
	// Trace: design.sv:106217:5
	input wire en_i;
	// Trace: design.sv:106218:5
	input wire scan_cg_en_i;
	// Trace: design.sv:106219:5
	output wire clk_o;
	// Trace: design.sv:106222:3
	reg clk_en;
	// Trace: design.sv:106224:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:106225:5
		if (clk_i == 1'b0)
			// Trace: design.sv:106225:24
			clk_en <= en_i | scan_cg_en_i;
	end
	// Trace: design.sv:106228:3
	assign clk_o = clk_i & clk_en;
	initial _sv2v_0 = 0;
endmodule
module cv32e40p_clock_gate (
	clk_i,
	en_i,
	scan_cg_en_i,
	clk_o
);
	reg _sv2v_0;
	// Trace: design.sv:106246:5
	input wire clk_i;
	// Trace: design.sv:106247:5
	input wire en_i;
	// Trace: design.sv:106248:5
	input wire scan_cg_en_i;
	// Trace: design.sv:106249:5
	output wire clk_o;
	// Trace: design.sv:106252:3
	reg clk_en;
	// Trace: design.sv:106254:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:106255:5
		if (clk_i == 1'b0)
			// Trace: design.sv:106255:24
			clk_en <= en_i | scan_cg_en_i;
	end
	// Trace: design.sv:106258:3
	assign clk_o = clk_i & clk_en;
	initial _sv2v_0 = 0;
endmodule
module pulp_clock_and2 (
	clk0_i,
	clk1_i,
	clk_o
);
	// Trace: design.sv:106272:3
	input wire clk0_i;
	// Trace: design.sv:106273:3
	input wire clk1_i;
	// Trace: design.sv:106274:3
	output wire clk_o;
	// Trace: design.sv:106277:3
	tc_clk_and2 i_tc_clk_and2(
		.clk0_i(clk0_i),
		.clk1_i(clk1_i),
		.clk_o(clk_o)
	);
endmodule
module pulp_clock_buffer (
	clk_i,
	clk_o
);
	// Trace: design.sv:106286:3
	input wire clk_i;
	// Trace: design.sv:106287:3
	output wire clk_o;
	// Trace: design.sv:106290:3
	tc_clk_buffer i_tc_clk_buffer(
		.clk_i(clk_i),
		.clk_o(clk_o)
	);
endmodule
module pulp_clock_gating (
	clk_i,
	en_i,
	test_en_i,
	clk_o
);
	// Trace: design.sv:106299:4
	input wire clk_i;
	// Trace: design.sv:106300:4
	input wire en_i;
	// Trace: design.sv:106301:4
	input wire test_en_i;
	// Trace: design.sv:106302:4
	output wire clk_o;
	// Trace: design.sv:106305:3
	tc_clk_gating i_tc_clk_gating(
		.clk_i(clk_i),
		.en_i(en_i),
		.test_en_i(test_en_i),
		.clk_o(clk_o)
	);
endmodule
module pulp_clock_inverter (
	clk_i,
	clk_o
);
	// Trace: design.sv:106315:3
	input wire clk_i;
	// Trace: design.sv:106316:3
	output wire clk_o;
	// Trace: design.sv:106319:3
	tc_clk_inverter i_tc_clk_inverter(
		.clk_i(clk_i),
		.clk_o(clk_o)
	);
endmodule
module pulp_clock_mux2 (
	clk0_i,
	clk1_i,
	clk_sel_i,
	clk_o
);
	// Trace: design.sv:106327:3
	input wire clk0_i;
	// Trace: design.sv:106328:3
	input wire clk1_i;
	// Trace: design.sv:106329:3
	input wire clk_sel_i;
	// Trace: design.sv:106330:3
	output wire clk_o;
	// Trace: design.sv:106333:3
	tc_clk_mux2 i_tc_clk_mux2(
		.clk0_i(clk0_i),
		.clk1_i(clk1_i),
		.clk_sel_i(clk_sel_i),
		.clk_o(clk_o)
	);
endmodule
module pulp_clock_xor2 (
	clk0_i,
	clk1_i,
	clk_o
);
	// Trace: design.sv:106343:3
	input wire clk0_i;
	// Trace: design.sv:106344:3
	input wire clk1_i;
	// Trace: design.sv:106345:3
	output wire clk_o;
	// Trace: design.sv:106348:3
	tc_clk_xor2 i_tc_clk_xor2(
		.clk0_i(clk0_i),
		.clk1_i(clk1_i),
		.clk_o(clk_o)
	);
endmodule
module cluster_clock_and2 (
	clk0_i,
	clk1_i,
	clk_o
);
	// Trace: design.sv:106379:3
	input wire clk0_i;
	// Trace: design.sv:106380:3
	input wire clk1_i;
	// Trace: design.sv:106381:3
	output wire clk_o;
	// Trace: design.sv:106384:3
	tc_clk_and2 i_tc_clk_and2(
		.clk0_i(clk0_i),
		.clk1_i(clk1_i),
		.clk_o(clk_o)
	);
endmodule
module cluster_clock_buffer (
	clk_i,
	clk_o
);
	// Trace: design.sv:106393:3
	input wire clk_i;
	// Trace: design.sv:106394:3
	output wire clk_o;
	// Trace: design.sv:106397:3
	tc_clk_buffer i_tc_clk_buffer(
		.clk_i(clk_i),
		.clk_o(clk_o)
	);
endmodule
module cluster_clock_gating (
	clk_i,
	en_i,
	test_en_i,
	clk_o
);
	// Trace: design.sv:106406:4
	input wire clk_i;
	// Trace: design.sv:106407:4
	input wire en_i;
	// Trace: design.sv:106408:4
	input wire test_en_i;
	// Trace: design.sv:106409:4
	output wire clk_o;
	// Trace: design.sv:106412:3
	tc_clk_gating i_tc_clk_gating(
		.clk_i(clk_i),
		.en_i(en_i),
		.test_en_i(test_en_i),
		.clk_o(clk_o)
	);
endmodule
module cluster_clock_inverter (
	clk_i,
	clk_o
);
	// Trace: design.sv:106422:3
	input wire clk_i;
	// Trace: design.sv:106423:3
	output wire clk_o;
	// Trace: design.sv:106426:3
	tc_clk_inverter i_tc_clk_inverter(
		.clk_i(clk_i),
		.clk_o(clk_o)
	);
endmodule
module cluster_clock_mux2 (
	clk0_i,
	clk1_i,
	clk_sel_i,
	clk_o
);
	// Trace: design.sv:106434:3
	input wire clk0_i;
	// Trace: design.sv:106435:3
	input wire clk1_i;
	// Trace: design.sv:106436:3
	input wire clk_sel_i;
	// Trace: design.sv:106437:3
	output wire clk_o;
	// Trace: design.sv:106440:3
	tc_clk_mux2 i_tc_clk_mux2(
		.clk0_i(clk0_i),
		.clk1_i(clk1_i),
		.clk_sel_i(clk_sel_i),
		.clk_o(clk_o)
	);
endmodule
module cluster_clock_xor2 (
	clk0_i,
	clk1_i,
	clk_o
);
	// Trace: design.sv:106450:3
	input wire clk0_i;
	// Trace: design.sv:106451:3
	input wire clk1_i;
	// Trace: design.sv:106452:3
	output wire clk_o;
	// Trace: design.sv:106455:3
	tc_clk_xor2 i_tc_clk_xor2(
		.clk0_i(clk0_i),
		.clk1_i(clk1_i),
		.clk_o(clk_o)
	);
endmodule
module tc_clk_and2 (
	clk0_i,
	clk1_i,
	clk_o
);
	// Trace: design.sv:106473:3
	input wire clk0_i;
	// Trace: design.sv:106474:3
	input wire clk1_i;
	// Trace: design.sv:106475:3
	output wire clk_o;
	// Trace: design.sv:106478:3
	assign clk_o = clk0_i & clk1_i;
endmodule
module tc_clk_buffer (
	clk_i,
	clk_o
);
	// Trace: design.sv:106483:3
	input wire clk_i;
	// Trace: design.sv:106484:3
	output wire clk_o;
	// Trace: design.sv:106487:3
	assign clk_o = clk_i;
endmodule
module tc_clk_gating (
	clk_i,
	en_i,
	test_en_i,
	clk_o
);
	reg _sv2v_0;
	// Trace: design.sv:106498:13
	parameter [0:0] IS_FUNCTIONAL = 1'b1;
	// Trace: design.sv:106500:4
	input wire clk_i;
	// Trace: design.sv:106501:4
	input wire en_i;
	// Trace: design.sv:106502:4
	input wire test_en_i;
	// Trace: design.sv:106503:4
	output wire clk_o;
	// Trace: design.sv:106506:3
	reg clk_en;
	// Trace: design.sv:106508:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: design.sv:106509:5
		if (clk_i == 1'b0)
			// Trace: design.sv:106509:24
			clk_en <= en_i | test_en_i;
	end
	// Trace: design.sv:106512:3
	assign clk_o = clk_i & clk_en;
	initial _sv2v_0 = 0;
endmodule
module tc_clk_inverter (
	clk_i,
	clk_o
);
	// Trace: design.sv:106517:3
	input wire clk_i;
	// Trace: design.sv:106518:3
	output wire clk_o;
	// Trace: design.sv:106521:3
	assign clk_o = ~clk_i;
endmodule
module tc_clk_mux2 (
	clk0_i,
	clk1_i,
	clk_sel_i,
	clk_o
);
	// Trace: design.sv:106526:3
	input wire clk0_i;
	// Trace: design.sv:106527:3
	input wire clk1_i;
	// Trace: design.sv:106528:3
	input wire clk_sel_i;
	// Trace: design.sv:106529:3
	output wire clk_o;
	// Trace: design.sv:106532:3
	assign clk_o = (clk_sel_i ? clk1_i : clk0_i);
endmodule
module tc_clk_xor2 (
	clk0_i,
	clk1_i,
	clk_o
);
	// Trace: design.sv:106537:3
	input wire clk0_i;
	// Trace: design.sv:106538:3
	input wire clk1_i;
	// Trace: design.sv:106539:3
	output wire clk_o;
	// Trace: design.sv:106542:3
	assign clk_o = clk0_i ^ clk1_i;
endmodule
module spimemio (
	clk,
	resetn,
	start_spi_i,
	valid,
	ready,
	addr,
	rdata,
	flash_csb,
	flash_clk,
	flash_io0_oe,
	flash_io1_oe,
	flash_io2_oe,
	flash_io3_oe,
	flash_io0_do,
	flash_io1_do,
	flash_io2_do,
	flash_io3_do,
	flash_io0_di,
	flash_io1_di,
	flash_io2_di,
	flash_io3_di,
	cfgreg_we,
	cfgreg_di,
	cfgreg_do
);
	// Trace: design.sv:106584:2
	input clk;
	input resetn;
	// Trace: design.sv:106585:2
	input start_spi_i;
	// Trace: design.sv:106586:2
	input valid;
	// Trace: design.sv:106587:2
	output wire ready;
	// Trace: design.sv:106588:2
	input [23:0] addr;
	// Trace: design.sv:106589:2
	output reg [31:0] rdata;
	// Trace: design.sv:106591:2
	output wire flash_csb;
	// Trace: design.sv:106592:2
	output wire flash_clk;
	// Trace: design.sv:106594:2
	output wire flash_io0_oe;
	// Trace: design.sv:106595:2
	output wire flash_io1_oe;
	// Trace: design.sv:106596:2
	output wire flash_io2_oe;
	// Trace: design.sv:106597:2
	output wire flash_io3_oe;
	// Trace: design.sv:106599:2
	output wire flash_io0_do;
	// Trace: design.sv:106600:2
	output wire flash_io1_do;
	// Trace: design.sv:106601:2
	output wire flash_io2_do;
	// Trace: design.sv:106602:2
	output wire flash_io3_do;
	// Trace: design.sv:106604:2
	input flash_io0_di;
	// Trace: design.sv:106605:2
	input flash_io1_di;
	// Trace: design.sv:106606:2
	input flash_io2_di;
	// Trace: design.sv:106607:2
	input flash_io3_di;
	// Trace: design.sv:106609:2
	input [3:0] cfgreg_we;
	// Trace: design.sv:106610:2
	input [31:0] cfgreg_di;
	// Trace: design.sv:106611:2
	output wire [31:0] cfgreg_do;
	// Trace: design.sv:106613:2
	reg xfer_resetn;
	// Trace: design.sv:106614:2
	reg din_valid;
	// Trace: design.sv:106615:2
	wire din_ready;
	// Trace: design.sv:106616:2
	reg [7:0] din_data;
	// Trace: design.sv:106617:2
	reg [3:0] din_tag;
	// Trace: design.sv:106618:2
	reg din_cont;
	// Trace: design.sv:106619:2
	reg din_qspi;
	// Trace: design.sv:106620:2
	reg din_ddr;
	// Trace: design.sv:106621:2
	reg din_rd;
	// Trace: design.sv:106623:2
	wire dout_valid;
	// Trace: design.sv:106624:2
	wire [7:0] dout_data;
	// Trace: design.sv:106625:2
	wire [3:0] dout_tag;
	// Trace: design.sv:106627:2
	reg [23:0] buffer;
	// Trace: design.sv:106629:2
	reg [23:0] rd_addr;
	// Trace: design.sv:106630:2
	reg rd_valid;
	// Trace: design.sv:106631:2
	reg rd_wait;
	// Trace: design.sv:106632:2
	reg rd_inc;
	// Trace: design.sv:106634:2
	assign ready = (valid && (addr == rd_addr)) && rd_valid;
	// Trace: design.sv:106635:2
	wire jump = ((valid && !ready) && (addr != (rd_addr + 4))) && rd_valid;
	// Trace: design.sv:106637:2
	reg softreset;
	// Trace: design.sv:106639:2
	reg config_en;
	// Trace: design.sv:106640:2
	reg config_ddr;
	// Trace: design.sv:106641:2
	reg config_qspi;
	// Trace: design.sv:106642:2
	reg config_cont;
	// Trace: design.sv:106643:2
	reg [3:0] config_dummy;
	// Trace: design.sv:106644:2
	reg [3:0] config_oe;
	// Trace: design.sv:106645:2
	reg config_csb;
	// Trace: design.sv:106646:2
	reg config_clk;
	// Trace: design.sv:106647:2
	reg [3:0] config_do;
	// Trace: design.sv:106649:2
	assign cfgreg_do[31] = config_en;
	// Trace: design.sv:106650:2
	assign cfgreg_do[30:23] = 0;
	// Trace: design.sv:106651:2
	assign cfgreg_do[22] = config_ddr;
	// Trace: design.sv:106652:2
	assign cfgreg_do[21] = config_qspi;
	// Trace: design.sv:106653:2
	assign cfgreg_do[20] = config_cont;
	// Trace: design.sv:106654:2
	assign cfgreg_do[19:16] = config_dummy;
	// Trace: design.sv:106655:2
	assign cfgreg_do[15:12] = 0;
	// Trace: design.sv:106656:2
	assign cfgreg_do[11:8] = {flash_io3_oe, flash_io2_oe, flash_io1_oe, flash_io0_oe};
	// Trace: design.sv:106657:2
	assign cfgreg_do[7:6] = 0;
	// Trace: design.sv:106658:2
	assign cfgreg_do[5] = flash_csb;
	// Trace: design.sv:106659:2
	assign cfgreg_do[4] = flash_clk;
	// Trace: design.sv:106660:2
	assign cfgreg_do[3:0] = {flash_io3_di, flash_io2_di, flash_io1_di, flash_io0_di};
	// Trace: design.sv:106662:2
	always @(posedge clk or negedge resetn)
		// Trace: design.sv:106663:3
		if (!resetn) begin
			// Trace: design.sv:106664:4
			softreset <= 1;
			// Trace: design.sv:106665:4
			config_en <= 1;
			// Trace: design.sv:106666:4
			config_csb <= 0;
			// Trace: design.sv:106667:4
			config_clk <= 0;
			// Trace: design.sv:106668:4
			config_oe <= 0;
			// Trace: design.sv:106669:4
			config_do <= 0;
			// Trace: design.sv:106670:4
			config_ddr <= 0;
			// Trace: design.sv:106671:4
			config_qspi <= 0;
			// Trace: design.sv:106672:4
			config_cont <= 0;
			// Trace: design.sv:106673:4
			config_dummy <= 8;
		end
		else begin
			// Trace: design.sv:106675:4
			softreset <= !config_en || cfgreg_we;
			// Trace: design.sv:106676:4
			if (cfgreg_we[0]) begin
				// Trace: design.sv:106677:5
				config_csb <= cfgreg_di[5];
				// Trace: design.sv:106678:5
				config_clk <= cfgreg_di[4];
				// Trace: design.sv:106679:5
				config_do <= cfgreg_di[3:0];
			end
			if (cfgreg_we[1])
				// Trace: design.sv:106682:5
				config_oe <= cfgreg_di[11:8];
			if (cfgreg_we[2]) begin
				// Trace: design.sv:106685:5
				config_ddr <= cfgreg_di[22];
				// Trace: design.sv:106686:5
				config_qspi <= cfgreg_di[21];
				// Trace: design.sv:106687:5
				config_cont <= cfgreg_di[20];
				// Trace: design.sv:106688:5
				config_dummy <= cfgreg_di[19:16];
			end
			if (cfgreg_we[3])
				// Trace: design.sv:106691:5
				config_en <= cfgreg_di[31];
		end
	// Trace: design.sv:106696:2
	wire xfer_csb;
	// Trace: design.sv:106697:2
	wire xfer_clk;
	// Trace: design.sv:106699:2
	wire xfer_io0_oe;
	// Trace: design.sv:106700:2
	wire xfer_io1_oe;
	// Trace: design.sv:106701:2
	wire xfer_io2_oe;
	// Trace: design.sv:106702:2
	wire xfer_io3_oe;
	// Trace: design.sv:106704:2
	wire xfer_io0_do;
	// Trace: design.sv:106705:2
	wire xfer_io1_do;
	// Trace: design.sv:106706:2
	wire xfer_io2_do;
	// Trace: design.sv:106707:2
	wire xfer_io3_do;
	// Trace: design.sv:106709:2
	reg xfer_io0_90;
	// Trace: design.sv:106710:2
	reg xfer_io1_90;
	// Trace: design.sv:106711:2
	reg xfer_io2_90;
	// Trace: design.sv:106712:2
	reg xfer_io3_90;
	// Trace: design.sv:106714:2
	always @(negedge clk) begin
		// Trace: design.sv:106715:3
		xfer_io0_90 <= xfer_io0_do;
		// Trace: design.sv:106716:3
		xfer_io1_90 <= xfer_io1_do;
		// Trace: design.sv:106717:3
		xfer_io2_90 <= xfer_io2_do;
		// Trace: design.sv:106718:3
		xfer_io3_90 <= xfer_io3_do;
	end
	// Trace: design.sv:106721:2
	assign flash_csb = (config_en ? xfer_csb : config_csb);
	// Trace: design.sv:106722:2
	assign flash_clk = (config_en ? xfer_clk : config_clk);
	// Trace: design.sv:106724:2
	assign flash_io0_oe = (config_en ? xfer_io0_oe : config_oe[0]);
	// Trace: design.sv:106725:2
	assign flash_io1_oe = (config_en ? xfer_io1_oe : config_oe[1]);
	// Trace: design.sv:106726:2
	assign flash_io2_oe = (config_en ? xfer_io2_oe : config_oe[2]);
	// Trace: design.sv:106727:2
	assign flash_io3_oe = (config_en ? xfer_io3_oe : config_oe[3]);
	// Trace: design.sv:106729:2
	assign flash_io0_do = (config_en ? (config_ddr ? xfer_io0_90 : xfer_io0_do) : config_do[0]);
	// Trace: design.sv:106730:2
	assign flash_io1_do = (config_en ? (config_ddr ? xfer_io1_90 : xfer_io1_do) : config_do[1]);
	// Trace: design.sv:106731:2
	assign flash_io2_do = (config_en ? (config_ddr ? xfer_io2_90 : xfer_io2_do) : config_do[2]);
	// Trace: design.sv:106732:2
	assign flash_io3_do = (config_en ? (config_ddr ? xfer_io3_90 : xfer_io3_do) : config_do[3]);
	// Trace: design.sv:106734:2
	wire xfer_dspi = din_ddr && !din_qspi;
	// Trace: design.sv:106735:2
	wire xfer_ddr = din_ddr && din_qspi;
	// Trace: design.sv:106737:2
	spimemio_xfer xfer(
		.clk(clk),
		.resetn(xfer_resetn),
		.din_valid(din_valid),
		.din_ready(din_ready),
		.din_data(din_data),
		.din_tag(din_tag),
		.din_cont(din_cont),
		.din_dspi(xfer_dspi),
		.din_qspi(din_qspi),
		.din_ddr(xfer_ddr),
		.din_rd(din_rd),
		.dout_valid(dout_valid),
		.dout_data(dout_data),
		.dout_tag(dout_tag),
		.flash_csb(xfer_csb),
		.flash_clk(xfer_clk),
		.flash_io0_oe(xfer_io0_oe),
		.flash_io1_oe(xfer_io1_oe),
		.flash_io2_oe(xfer_io2_oe),
		.flash_io3_oe(xfer_io3_oe),
		.flash_io0_do(xfer_io0_do),
		.flash_io1_do(xfer_io1_do),
		.flash_io2_do(xfer_io2_do),
		.flash_io3_do(xfer_io3_do),
		.flash_io0_di(flash_io0_di),
		.flash_io1_di(flash_io1_di),
		.flash_io2_di(flash_io2_di),
		.flash_io3_di(flash_io3_di)
	);
	// Trace: design.sv:106768:2
	reg [3:0] state;
	// Trace: design.sv:106770:2
	always @(posedge clk or negedge resetn)
		// Trace: design.sv:106771:3
		if (!resetn) begin
			// Trace: design.sv:106772:4
			xfer_resetn <= 1;
			// Trace: design.sv:106773:4
			din_valid <= 0;
			// Trace: design.sv:106774:4
			state <= 0;
			// Trace: design.sv:106775:4
			xfer_resetn <= 0;
			// Trace: design.sv:106776:4
			rd_valid <= 0;
			// Trace: design.sv:106777:4
			din_tag <= 0;
			// Trace: design.sv:106778:4
			din_cont <= 0;
			// Trace: design.sv:106779:4
			din_qspi <= 0;
			// Trace: design.sv:106780:4
			din_ddr <= 0;
			// Trace: design.sv:106781:4
			din_rd <= 0;
		end
		else
			// Trace: design.sv:106784:4
			if (softreset) begin
				// Trace: design.sv:106785:5
				xfer_resetn <= 1;
				// Trace: design.sv:106786:5
				din_valid <= 0;
				// Trace: design.sv:106787:5
				state <= 0;
				// Trace: design.sv:106788:5
				xfer_resetn <= 0;
				// Trace: design.sv:106789:5
				rd_valid <= 0;
				// Trace: design.sv:106790:5
				din_tag <= 0;
				// Trace: design.sv:106791:5
				din_cont <= 0;
				// Trace: design.sv:106792:5
				din_qspi <= 0;
				// Trace: design.sv:106793:5
				din_ddr <= 0;
				// Trace: design.sv:106794:5
				din_rd <= 0;
			end
			else begin
				// Trace: design.sv:106796:5
				xfer_resetn <= 1;
				// Trace: design.sv:106797:5
				din_valid <= 0;
				// Trace: design.sv:106798:5
				if (dout_valid && (dout_tag == 1))
					// Trace: design.sv:106798:38
					buffer[7:0] <= dout_data;
				if (dout_valid && (dout_tag == 2))
					// Trace: design.sv:106799:38
					buffer[15:8] <= dout_data;
				if (dout_valid && (dout_tag == 3))
					// Trace: design.sv:106800:38
					buffer[23:16] <= dout_data;
				if (dout_valid && (dout_tag == 4)) begin
					// Trace: design.sv:106802:6
					rdata <= {dout_data, buffer};
					// Trace: design.sv:106803:6
					rd_addr <= (rd_inc ? rd_addr + 4 : addr);
					// Trace: design.sv:106804:6
					rd_valid <= 1;
					// Trace: design.sv:106805:6
					rd_wait <= rd_inc;
					// Trace: design.sv:106806:6
					rd_inc <= 1;
				end
				if (valid)
					// Trace: design.sv:106810:6
					rd_wait <= 0;
				case (state)
					0: begin
						// Trace: design.sv:106814:7
						din_valid <= start_spi_i;
						// Trace: design.sv:106815:7
						din_data <= 8'hff;
						// Trace: design.sv:106816:7
						din_tag <= 0;
						// Trace: design.sv:106817:7
						if (din_ready) begin
							// Trace: design.sv:106818:8
							din_valid <= 0;
							// Trace: design.sv:106819:8
							state <= 1;
						end
					end
					1:
						// Trace: design.sv:106823:7
						if (dout_valid) begin
							// Trace: design.sv:106824:8
							xfer_resetn <= 0;
							// Trace: design.sv:106825:8
							state <= 2;
						end
					2: begin
						// Trace: design.sv:106829:7
						din_valid <= 1;
						// Trace: design.sv:106830:7
						din_data <= 8'hab;
						// Trace: design.sv:106831:7
						din_tag <= 0;
						// Trace: design.sv:106832:7
						if (din_ready) begin
							// Trace: design.sv:106833:8
							din_valid <= 0;
							// Trace: design.sv:106834:8
							state <= 3;
						end
					end
					3:
						// Trace: design.sv:106838:7
						if (dout_valid) begin
							// Trace: design.sv:106839:8
							xfer_resetn <= 0;
							// Trace: design.sv:106840:8
							state <= 4;
						end
					4: begin
						// Trace: design.sv:106844:7
						rd_inc <= 0;
						// Trace: design.sv:106845:7
						din_valid <= 1;
						// Trace: design.sv:106846:7
						din_tag <= 0;
						// Trace: design.sv:106847:7
						case ({config_ddr, config_qspi})
							2'b11:
								// Trace: design.sv:106848:15
								din_data <= 8'hed;
							2'b01:
								// Trace: design.sv:106849:15
								din_data <= 8'heb;
							2'b10:
								// Trace: design.sv:106850:15
								din_data <= 8'hbb;
							2'b00:
								// Trace: design.sv:106851:15
								din_data <= 8'h03;
						endcase
						if (din_ready) begin
							// Trace: design.sv:106854:8
							din_valid <= 0;
							// Trace: design.sv:106855:8
							state <= 5;
						end
					end
					5:
						// Trace: design.sv:106859:7
						if (valid && !ready) begin
							// Trace: design.sv:106860:8
							din_valid <= 1;
							// Trace: design.sv:106861:8
							din_tag <= 0;
							// Trace: design.sv:106862:8
							din_data <= addr[23:16];
							// Trace: design.sv:106863:8
							din_qspi <= config_qspi;
							// Trace: design.sv:106864:8
							din_ddr <= config_ddr;
							// Trace: design.sv:106865:8
							if (din_ready) begin
								// Trace: design.sv:106866:9
								din_valid <= 0;
								// Trace: design.sv:106867:9
								state <= 6;
							end
						end
					6: begin
						// Trace: design.sv:106872:7
						din_valid <= 1;
						// Trace: design.sv:106873:7
						din_tag <= 0;
						// Trace: design.sv:106874:7
						din_data <= addr[15:8];
						// Trace: design.sv:106875:7
						if (din_ready) begin
							// Trace: design.sv:106876:8
							din_valid <= 0;
							// Trace: design.sv:106877:8
							state <= 7;
						end
					end
					7: begin
						// Trace: design.sv:106881:7
						din_valid <= 1;
						// Trace: design.sv:106882:7
						din_tag <= 0;
						// Trace: design.sv:106883:7
						din_data <= addr[7:0];
						// Trace: design.sv:106884:7
						if (din_ready) begin
							// Trace: design.sv:106885:8
							din_valid <= 0;
							// Trace: design.sv:106886:8
							din_data <= 0;
							// Trace: design.sv:106887:8
							state <= (config_qspi || config_ddr ? 8 : 9);
						end
					end
					8: begin
						// Trace: design.sv:106891:7
						din_valid <= 1;
						// Trace: design.sv:106892:7
						din_tag <= 0;
						// Trace: design.sv:106893:7
						din_data <= (config_cont ? 8'ha5 : 8'hff);
						// Trace: design.sv:106894:7
						if (din_ready) begin
							// Trace: design.sv:106895:8
							din_rd <= 1;
							// Trace: design.sv:106896:8
							din_data <= config_dummy;
							// Trace: design.sv:106897:8
							din_valid <= 0;
							// Trace: design.sv:106898:8
							state <= 9;
						end
					end
					9: begin
						// Trace: design.sv:106902:7
						din_valid <= 1;
						// Trace: design.sv:106903:7
						din_tag <= 1;
						// Trace: design.sv:106904:7
						if (din_ready) begin
							// Trace: design.sv:106905:8
							din_valid <= 0;
							// Trace: design.sv:106906:8
							state <= 10;
						end
					end
					10: begin
						// Trace: design.sv:106910:7
						din_valid <= 1;
						// Trace: design.sv:106911:7
						din_data <= 8'h00;
						// Trace: design.sv:106912:7
						din_tag <= 2;
						// Trace: design.sv:106913:7
						if (din_ready) begin
							// Trace: design.sv:106914:8
							din_valid <= 0;
							// Trace: design.sv:106915:8
							state <= 11;
						end
					end
					11: begin
						// Trace: design.sv:106919:7
						din_valid <= 1;
						// Trace: design.sv:106920:7
						din_tag <= 3;
						// Trace: design.sv:106921:7
						if (din_ready) begin
							// Trace: design.sv:106922:8
							din_valid <= 0;
							// Trace: design.sv:106923:8
							state <= 12;
						end
					end
					12:
						// Trace: design.sv:106927:7
						if (!rd_wait || valid) begin
							// Trace: design.sv:106928:8
							din_valid <= 1;
							// Trace: design.sv:106929:8
							din_tag <= 4;
							// Trace: design.sv:106930:8
							if (din_ready) begin
								// Trace: design.sv:106931:9
								din_valid <= 0;
								// Trace: design.sv:106932:9
								state <= 9;
							end
						end
				endcase
				if (jump) begin
					// Trace: design.sv:106939:6
					rd_inc <= 0;
					// Trace: design.sv:106940:6
					rd_valid <= 0;
					// Trace: design.sv:106941:6
					xfer_resetn <= 0;
					// Trace: design.sv:106942:6
					if (config_cont)
						// Trace: design.sv:106943:7
						state <= 5;
					else begin
						// Trace: design.sv:106945:7
						state <= 4;
						// Trace: design.sv:106946:7
						din_qspi <= 0;
						// Trace: design.sv:106947:7
						din_ddr <= 0;
					end
					// Trace: design.sv:106949:6
					din_rd <= 0;
				end
			end
endmodule
module spimemio_xfer (
	clk,
	resetn,
	din_valid,
	din_ready,
	din_data,
	din_tag,
	din_cont,
	din_dspi,
	din_qspi,
	din_ddr,
	din_rd,
	dout_valid,
	dout_data,
	dout_tag,
	flash_csb,
	flash_clk,
	flash_io0_oe,
	flash_io1_oe,
	flash_io2_oe,
	flash_io3_oe,
	flash_io0_do,
	flash_io1_do,
	flash_io2_do,
	flash_io3_do,
	flash_io0_di,
	flash_io1_di,
	flash_io2_di,
	flash_io3_di
);
	// Trace: design.sv:106957:2
	input clk;
	input resetn;
	// Trace: design.sv:106959:2
	input din_valid;
	// Trace: design.sv:106960:2
	output wire din_ready;
	// Trace: design.sv:106961:2
	input [7:0] din_data;
	// Trace: design.sv:106962:2
	input [3:0] din_tag;
	// Trace: design.sv:106963:2
	input din_cont;
	// Trace: design.sv:106964:2
	input din_dspi;
	// Trace: design.sv:106965:2
	input din_qspi;
	// Trace: design.sv:106966:2
	input din_ddr;
	// Trace: design.sv:106967:2
	input din_rd;
	// Trace: design.sv:106969:2
	output wire dout_valid;
	// Trace: design.sv:106970:2
	output wire [7:0] dout_data;
	// Trace: design.sv:106971:2
	output wire [3:0] dout_tag;
	// Trace: design.sv:106973:2
	output reg flash_csb;
	// Trace: design.sv:106974:2
	output reg flash_clk;
	// Trace: design.sv:106976:2
	output reg flash_io0_oe;
	// Trace: design.sv:106977:2
	output reg flash_io1_oe;
	// Trace: design.sv:106978:2
	output reg flash_io2_oe;
	// Trace: design.sv:106979:2
	output reg flash_io3_oe;
	// Trace: design.sv:106981:2
	output reg flash_io0_do;
	// Trace: design.sv:106982:2
	output reg flash_io1_do;
	// Trace: design.sv:106983:2
	output reg flash_io2_do;
	// Trace: design.sv:106984:2
	output reg flash_io3_do;
	// Trace: design.sv:106986:2
	input flash_io0_di;
	// Trace: design.sv:106987:2
	input flash_io1_di;
	// Trace: design.sv:106988:2
	input flash_io2_di;
	// Trace: design.sv:106989:2
	input flash_io3_di;
	// Trace: design.sv:106991:2
	reg [7:0] obuffer;
	// Trace: design.sv:106992:2
	reg [7:0] ibuffer;
	// Trace: design.sv:106994:2
	reg [3:0] count;
	// Trace: design.sv:106995:2
	reg [3:0] dummy_count;
	// Trace: design.sv:106997:2
	reg xfer_cont;
	// Trace: design.sv:106998:2
	reg xfer_dspi;
	// Trace: design.sv:106999:2
	reg xfer_qspi;
	// Trace: design.sv:107000:2
	reg xfer_ddr;
	// Trace: design.sv:107001:2
	reg xfer_ddr_q;
	// Trace: design.sv:107002:2
	reg xfer_rd;
	// Trace: design.sv:107003:2
	reg [3:0] xfer_tag;
	// Trace: design.sv:107004:2
	reg [3:0] xfer_tag_q;
	// Trace: design.sv:107006:2
	reg [7:0] next_obuffer;
	// Trace: design.sv:107007:2
	reg [7:0] next_ibuffer;
	// Trace: design.sv:107008:2
	reg [3:0] next_count;
	// Trace: design.sv:107010:2
	reg fetch;
	// Trace: design.sv:107011:2
	reg next_fetch;
	// Trace: design.sv:107012:2
	reg last_fetch;
	// Trace: design.sv:107014:2
	always @(posedge clk) begin
		// Trace: design.sv:107015:3
		xfer_ddr_q <= xfer_ddr;
		// Trace: design.sv:107016:3
		xfer_tag_q <= xfer_tag;
	end
	// Trace: design.sv:107019:2
	assign din_ready = (din_valid && resetn) && next_fetch;
	// Trace: design.sv:107021:2
	assign dout_valid = (xfer_ddr_q ? fetch && !last_fetch : next_fetch && !fetch) && resetn;
	// Trace: design.sv:107022:2
	assign dout_data = ibuffer;
	// Trace: design.sv:107023:2
	assign dout_tag = xfer_tag_q;
	// Trace: design.sv:107025:2
	always @(*) begin
		// Trace: design.sv:107026:3
		flash_io0_oe = 0;
		// Trace: design.sv:107027:3
		flash_io1_oe = 0;
		// Trace: design.sv:107028:3
		flash_io2_oe = 0;
		// Trace: design.sv:107029:3
		flash_io3_oe = 0;
		// Trace: design.sv:107031:3
		flash_io0_do = 0;
		// Trace: design.sv:107032:3
		flash_io1_do = 0;
		// Trace: design.sv:107033:3
		flash_io2_do = 0;
		// Trace: design.sv:107034:3
		flash_io3_do = 0;
		// Trace: design.sv:107036:3
		next_obuffer = obuffer;
		// Trace: design.sv:107037:3
		next_ibuffer = ibuffer;
		// Trace: design.sv:107038:3
		next_count = count;
		// Trace: design.sv:107039:3
		next_fetch = 0;
		// Trace: design.sv:107041:3
		if (dummy_count == 0)
			// Trace: design.sv:107042:4
			casez ({xfer_ddr, xfer_qspi, xfer_dspi})
				3'b000: begin
					// Trace: design.sv:107044:6
					flash_io0_oe = 1;
					// Trace: design.sv:107045:6
					flash_io0_do = obuffer[7];
					// Trace: design.sv:107047:6
					if (flash_clk) begin
						// Trace: design.sv:107048:7
						next_obuffer = {obuffer[6:0], 1'b0};
						// Trace: design.sv:107049:7
						next_count = count - |count;
					end
					else
						// Trace: design.sv:107051:7
						next_ibuffer = {ibuffer[6:0], flash_io1_di};
					// Trace: design.sv:107054:6
					next_fetch = next_count == 0;
				end
				3'b01z: begin
					// Trace: design.sv:107057:6
					flash_io0_oe = !xfer_rd;
					// Trace: design.sv:107058:6
					flash_io1_oe = !xfer_rd;
					// Trace: design.sv:107059:6
					flash_io2_oe = !xfer_rd;
					// Trace: design.sv:107060:6
					flash_io3_oe = !xfer_rd;
					// Trace: design.sv:107062:6
					flash_io0_do = obuffer[4];
					// Trace: design.sv:107063:6
					flash_io1_do = obuffer[5];
					// Trace: design.sv:107064:6
					flash_io2_do = obuffer[6];
					// Trace: design.sv:107065:6
					flash_io3_do = obuffer[7];
					// Trace: design.sv:107067:6
					if (flash_clk) begin
						// Trace: design.sv:107068:7
						next_obuffer = {obuffer[3:0], 4'b0000};
						// Trace: design.sv:107069:7
						next_count = count - {|count, 2'b00};
					end
					else
						// Trace: design.sv:107071:7
						next_ibuffer = {ibuffer[3:0], flash_io3_di, flash_io2_di, flash_io1_di, flash_io0_di};
					// Trace: design.sv:107074:6
					next_fetch = next_count == 0;
				end
				3'b11z: begin
					// Trace: design.sv:107077:6
					flash_io0_oe = !xfer_rd;
					// Trace: design.sv:107078:6
					flash_io1_oe = !xfer_rd;
					// Trace: design.sv:107079:6
					flash_io2_oe = !xfer_rd;
					// Trace: design.sv:107080:6
					flash_io3_oe = !xfer_rd;
					// Trace: design.sv:107082:6
					flash_io0_do = obuffer[4];
					// Trace: design.sv:107083:6
					flash_io1_do = obuffer[5];
					// Trace: design.sv:107084:6
					flash_io2_do = obuffer[6];
					// Trace: design.sv:107085:6
					flash_io3_do = obuffer[7];
					// Trace: design.sv:107087:6
					next_obuffer = {obuffer[3:0], 4'b0000};
					// Trace: design.sv:107088:6
					next_ibuffer = {ibuffer[3:0], flash_io3_di, flash_io2_di, flash_io1_di, flash_io0_di};
					// Trace: design.sv:107089:6
					next_count = count - {|count, 2'b00};
					// Trace: design.sv:107091:6
					next_fetch = next_count == 0;
				end
				3'bzz1: begin
					// Trace: design.sv:107094:6
					flash_io0_oe = !xfer_rd;
					// Trace: design.sv:107095:6
					flash_io1_oe = !xfer_rd;
					// Trace: design.sv:107097:6
					flash_io0_do = obuffer[6];
					// Trace: design.sv:107098:6
					flash_io1_do = obuffer[7];
					// Trace: design.sv:107100:6
					if (flash_clk) begin
						// Trace: design.sv:107101:7
						next_obuffer = {obuffer[5:0], 2'b00};
						// Trace: design.sv:107102:7
						next_count = count - {|count, 1'b0};
					end
					else
						// Trace: design.sv:107104:7
						next_ibuffer = {ibuffer[5:0], flash_io1_di, flash_io0_di};
					// Trace: design.sv:107107:6
					next_fetch = next_count == 0;
				end
			endcase
	end
	// Trace: design.sv:107113:2
	always @(posedge clk or negedge resetn)
		// Trace: design.sv:107114:3
		if (!resetn) begin
			// Trace: design.sv:107115:4
			fetch <= 1;
			// Trace: design.sv:107116:4
			last_fetch <= 1;
			// Trace: design.sv:107117:4
			flash_csb <= 1;
			// Trace: design.sv:107118:4
			flash_clk <= 0;
			// Trace: design.sv:107119:4
			count <= 0;
			// Trace: design.sv:107120:4
			dummy_count <= 0;
			// Trace: design.sv:107121:4
			xfer_tag <= 0;
			// Trace: design.sv:107122:4
			xfer_cont <= 0;
			// Trace: design.sv:107123:4
			xfer_dspi <= 0;
			// Trace: design.sv:107124:4
			xfer_qspi <= 0;
			// Trace: design.sv:107125:4
			xfer_ddr <= 0;
			// Trace: design.sv:107126:4
			xfer_rd <= 0;
		end
		else begin
			// Trace: design.sv:107128:4
			fetch <= next_fetch;
			// Trace: design.sv:107129:4
			last_fetch <= (xfer_ddr ? fetch : 1);
			// Trace: design.sv:107130:4
			if (dummy_count) begin
				// Trace: design.sv:107131:5
				flash_clk <= !flash_clk && !flash_csb;
				// Trace: design.sv:107132:5
				dummy_count <= dummy_count - flash_clk;
			end
			else if (count) begin
				// Trace: design.sv:107135:5
				flash_clk <= !flash_clk && !flash_csb;
				// Trace: design.sv:107136:5
				obuffer <= next_obuffer;
				// Trace: design.sv:107137:5
				ibuffer <= next_ibuffer;
				// Trace: design.sv:107138:5
				count <= next_count;
			end
			if (din_valid && din_ready) begin
				// Trace: design.sv:107141:5
				flash_csb <= 0;
				// Trace: design.sv:107142:5
				flash_clk <= 0;
				// Trace: design.sv:107144:5
				count <= 8;
				// Trace: design.sv:107145:5
				dummy_count <= (din_rd ? din_data : 0);
				// Trace: design.sv:107146:5
				obuffer <= din_data;
				// Trace: design.sv:107148:5
				xfer_tag <= din_tag;
				// Trace: design.sv:107149:5
				xfer_cont <= din_cont;
				// Trace: design.sv:107150:5
				xfer_dspi <= din_dspi;
				// Trace: design.sv:107151:5
				xfer_qspi <= din_qspi;
				// Trace: design.sv:107152:5
				xfer_ddr <= din_ddr;
				// Trace: design.sv:107153:5
				xfer_rd <= din_rd;
			end
		end
endmodule
